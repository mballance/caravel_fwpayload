VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1496.910 84.900 1497.230 84.960 ;
        RECT 1555.790 84.900 1556.110 84.960 ;
        RECT 1496.910 84.760 1556.110 84.900 ;
        RECT 1496.910 84.700 1497.230 84.760 ;
        RECT 1555.790 84.700 1556.110 84.760 ;
        RECT 2089.390 83.880 2089.710 83.940 ;
        RECT 2090.770 83.880 2091.090 83.940 ;
        RECT 2089.390 83.740 2091.090 83.880 ;
        RECT 2089.390 83.680 2089.710 83.740 ;
        RECT 2090.770 83.680 2091.090 83.740 ;
        RECT 2185.990 83.880 2186.310 83.940 ;
        RECT 2187.370 83.880 2187.690 83.940 ;
        RECT 2185.990 83.740 2187.690 83.880 ;
        RECT 2185.990 83.680 2186.310 83.740 ;
        RECT 2187.370 83.680 2187.690 83.740 ;
        RECT 2318.930 83.540 2319.250 83.600 ;
        RECT 2332.730 83.540 2333.050 83.600 ;
        RECT 2318.930 83.400 2333.050 83.540 ;
        RECT 2318.930 83.340 2319.250 83.400 ;
        RECT 2332.730 83.340 2333.050 83.400 ;
      LAYER via ;
        RECT 1496.940 84.700 1497.200 84.960 ;
        RECT 1555.820 84.700 1556.080 84.960 ;
        RECT 2089.420 83.680 2089.680 83.940 ;
        RECT 2090.800 83.680 2091.060 83.940 ;
        RECT 2186.020 83.680 2186.280 83.940 ;
        RECT 2187.400 83.680 2187.660 83.940 ;
        RECT 2318.960 83.340 2319.220 83.600 ;
        RECT 2332.760 83.340 2333.020 83.600 ;
      LAYER met2 ;
        RECT 1154.165 2896.530 1154.445 2900.000 ;
        RECT 1155.610 2896.530 1155.890 2896.645 ;
        RECT 1154.165 2896.390 1155.890 2896.530 ;
        RECT 1154.165 2896.000 1154.445 2896.390 ;
        RECT 1155.610 2896.275 1155.890 2896.390 ;
        RECT 2414.630 85.835 2414.910 86.205 ;
        RECT 1555.810 85.155 1556.090 85.525 ;
        RECT 1586.630 85.155 1586.910 85.525 ;
        RECT 1683.230 85.155 1683.510 85.525 ;
        RECT 1555.880 84.990 1556.020 85.155 ;
        RECT 1328.110 84.475 1328.390 84.845 ;
        RECT 1441.730 84.475 1442.010 84.845 ;
        RECT 1496.940 84.670 1497.200 84.990 ;
        RECT 1555.820 84.670 1556.080 84.990 ;
        RECT 1328.180 82.125 1328.320 84.475 ;
        RECT 1441.800 84.165 1441.940 84.475 ;
        RECT 1497.000 84.165 1497.140 84.670 ;
        RECT 1441.730 83.795 1442.010 84.165 ;
        RECT 1496.930 83.795 1497.210 84.165 ;
        RECT 1586.700 83.485 1586.840 85.155 ;
        RECT 1611.010 83.795 1611.290 84.165 ;
        RECT 1586.630 83.115 1586.910 83.485 ;
        RECT 1611.080 82.125 1611.220 83.795 ;
        RECT 1683.300 83.485 1683.440 85.155 ;
        RECT 2332.750 84.475 2333.030 84.845 ;
        RECT 2089.410 83.795 2089.690 84.165 ;
        RECT 2090.790 83.795 2091.070 84.165 ;
        RECT 2186.010 83.795 2186.290 84.165 ;
        RECT 2187.390 83.795 2187.670 84.165 ;
        RECT 2089.420 83.650 2089.680 83.795 ;
        RECT 2090.800 83.650 2091.060 83.795 ;
        RECT 2186.020 83.650 2186.280 83.795 ;
        RECT 2187.400 83.650 2187.660 83.795 ;
        RECT 2332.820 83.630 2332.960 84.475 ;
        RECT 2414.700 84.165 2414.840 85.835 ;
        RECT 2439.010 85.155 2439.290 85.525 ;
        RECT 2414.630 83.795 2414.910 84.165 ;
        RECT 2318.960 83.485 2319.220 83.630 ;
        RECT 1683.230 83.115 1683.510 83.485 ;
        RECT 2318.950 83.115 2319.230 83.485 ;
        RECT 2332.760 83.310 2333.020 83.630 ;
        RECT 2439.080 83.485 2439.220 85.155 ;
        RECT 2439.010 83.115 2439.290 83.485 ;
        RECT 1328.110 81.755 1328.390 82.125 ;
        RECT 1611.010 81.755 1611.290 82.125 ;
      LAYER via2 ;
        RECT 1155.610 2896.320 1155.890 2896.600 ;
        RECT 2414.630 85.880 2414.910 86.160 ;
        RECT 1555.810 85.200 1556.090 85.480 ;
        RECT 1586.630 85.200 1586.910 85.480 ;
        RECT 1683.230 85.200 1683.510 85.480 ;
        RECT 1328.110 84.520 1328.390 84.800 ;
        RECT 1441.730 84.520 1442.010 84.800 ;
        RECT 1441.730 83.840 1442.010 84.120 ;
        RECT 1496.930 83.840 1497.210 84.120 ;
        RECT 1611.010 83.840 1611.290 84.120 ;
        RECT 1586.630 83.160 1586.910 83.440 ;
        RECT 2332.750 84.520 2333.030 84.800 ;
        RECT 2089.410 83.840 2089.690 84.120 ;
        RECT 2090.790 83.840 2091.070 84.120 ;
        RECT 2186.010 83.840 2186.290 84.120 ;
        RECT 2187.390 83.840 2187.670 84.120 ;
        RECT 2439.010 85.200 2439.290 85.480 ;
        RECT 2414.630 83.840 2414.910 84.120 ;
        RECT 1683.230 83.160 1683.510 83.440 ;
        RECT 2318.950 83.160 2319.230 83.440 ;
        RECT 2439.010 83.160 2439.290 83.440 ;
        RECT 1328.110 81.800 1328.390 82.080 ;
        RECT 1611.010 81.800 1611.290 82.080 ;
      LAYER met3 ;
        RECT 1155.585 2896.610 1155.915 2896.625 ;
        RECT 1158.550 2896.610 1158.930 2896.620 ;
        RECT 1155.585 2896.310 1158.930 2896.610 ;
        RECT 1155.585 2896.295 1155.915 2896.310 ;
        RECT 1158.550 2896.300 1158.930 2896.310 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2916.710 87.910 2924.800 88.210 ;
        RECT 2366.510 86.170 2366.890 86.180 ;
        RECT 2414.605 86.170 2414.935 86.185 ;
        RECT 2366.510 85.870 2414.935 86.170 ;
        RECT 2366.510 85.860 2366.890 85.870 ;
        RECT 2414.605 85.855 2414.935 85.870 ;
        RECT 1555.785 85.490 1556.115 85.505 ;
        RECT 1586.605 85.490 1586.935 85.505 ;
        RECT 1683.205 85.490 1683.535 85.505 ;
        RECT 2027.030 85.490 2027.410 85.500 ;
        RECT 2316.830 85.490 2317.210 85.500 ;
        RECT 2438.985 85.490 2439.315 85.505 ;
        RECT 1555.785 85.190 1586.935 85.490 ;
        RECT 1555.785 85.175 1556.115 85.190 ;
        RECT 1586.605 85.175 1586.935 85.190 ;
        RECT 1635.150 85.190 1683.535 85.490 ;
        RECT 1328.085 84.810 1328.415 84.825 ;
        RECT 1441.705 84.810 1442.035 84.825 ;
        RECT 1328.085 84.510 1352.090 84.810 ;
        RECT 1328.085 84.495 1328.415 84.510 ;
        RECT 1158.550 84.130 1158.930 84.140 ;
        RECT 1158.550 83.830 1225.130 84.130 ;
        RECT 1158.550 83.820 1158.930 83.830 ;
        RECT 1224.830 83.450 1225.130 83.830 ;
        RECT 1224.830 83.150 1249.970 83.450 ;
        RECT 1249.670 82.090 1249.970 83.150 ;
        RECT 1351.790 82.770 1352.090 84.510 ;
        RECT 1441.705 84.510 1448.690 84.810 ;
        RECT 1441.705 84.495 1442.035 84.510 ;
        RECT 1441.705 84.130 1442.035 84.145 ;
        RECT 1394.110 83.830 1442.035 84.130 ;
        RECT 1448.390 84.130 1448.690 84.510 ;
        RECT 1496.905 84.130 1497.235 84.145 ;
        RECT 1448.390 83.830 1497.235 84.130 ;
        RECT 1394.110 83.450 1394.410 83.830 ;
        RECT 1441.705 83.815 1442.035 83.830 ;
        RECT 1496.905 83.815 1497.235 83.830 ;
        RECT 1610.985 84.130 1611.315 84.145 ;
        RECT 1635.150 84.130 1635.450 85.190 ;
        RECT 1683.205 85.175 1683.535 85.190 ;
        RECT 1993.030 85.190 2027.410 85.490 ;
        RECT 1610.985 83.830 1635.450 84.130 ;
        RECT 1704.150 84.510 1801.050 84.810 ;
        RECT 1610.985 83.815 1611.315 83.830 ;
        RECT 1366.510 83.150 1394.410 83.450 ;
        RECT 1586.605 83.450 1586.935 83.465 ;
        RECT 1683.205 83.450 1683.535 83.465 ;
        RECT 1704.150 83.450 1704.450 84.510 ;
        RECT 1800.750 84.130 1801.050 84.510 ;
        RECT 1993.030 84.130 1993.330 85.190 ;
        RECT 2027.030 85.180 2027.410 85.190 ;
        RECT 2282.830 85.190 2317.210 85.490 ;
        RECT 2089.385 84.130 2089.715 84.145 ;
        RECT 1800.750 83.830 1848.890 84.130 ;
        RECT 1586.605 83.150 1587.610 83.450 ;
        RECT 1366.510 82.770 1366.810 83.150 ;
        RECT 1586.605 83.135 1586.935 83.150 ;
        RECT 1351.790 82.470 1366.810 82.770 ;
        RECT 1328.085 82.090 1328.415 82.105 ;
        RECT 1249.670 81.790 1328.415 82.090 ;
        RECT 1587.310 82.090 1587.610 83.150 ;
        RECT 1683.205 83.150 1704.450 83.450 ;
        RECT 1848.590 83.450 1848.890 83.830 ;
        RECT 1942.430 83.830 1993.330 84.130 ;
        RECT 2042.710 83.830 2089.715 84.130 ;
        RECT 1942.430 83.450 1942.730 83.830 ;
        RECT 1848.590 83.150 1942.730 83.450 ;
        RECT 2027.950 83.450 2028.330 83.460 ;
        RECT 2042.710 83.450 2043.010 83.830 ;
        RECT 2089.385 83.815 2089.715 83.830 ;
        RECT 2090.765 84.130 2091.095 84.145 ;
        RECT 2185.985 84.130 2186.315 84.145 ;
        RECT 2090.765 83.830 2124.890 84.130 ;
        RECT 2090.765 83.815 2091.095 83.830 ;
        RECT 2027.950 83.150 2043.010 83.450 ;
        RECT 2124.590 83.450 2124.890 83.830 ;
        RECT 2139.310 83.830 2186.315 84.130 ;
        RECT 2139.310 83.450 2139.610 83.830 ;
        RECT 2185.985 83.815 2186.315 83.830 ;
        RECT 2187.365 84.130 2187.695 84.145 ;
        RECT 2282.830 84.130 2283.130 85.190 ;
        RECT 2316.830 85.180 2317.210 85.190 ;
        RECT 2415.310 85.190 2439.315 85.490 ;
        RECT 2332.725 84.810 2333.055 84.825 ;
        RECT 2366.510 84.810 2366.890 84.820 ;
        RECT 2332.725 84.510 2366.890 84.810 ;
        RECT 2332.725 84.495 2333.055 84.510 ;
        RECT 2366.510 84.500 2366.890 84.510 ;
        RECT 2187.365 83.830 2221.490 84.130 ;
        RECT 2187.365 83.815 2187.695 83.830 ;
        RECT 2124.590 83.150 2139.610 83.450 ;
        RECT 2221.190 83.450 2221.490 83.830 ;
        RECT 2235.910 83.830 2283.130 84.130 ;
        RECT 2414.605 84.130 2414.935 84.145 ;
        RECT 2415.310 84.130 2415.610 85.190 ;
        RECT 2438.985 85.175 2439.315 85.190 ;
        RECT 2463.110 84.810 2463.490 84.820 ;
        RECT 2463.110 84.510 2546.250 84.810 ;
        RECT 2463.110 84.500 2463.490 84.510 ;
        RECT 2414.605 83.830 2415.610 84.130 ;
        RECT 2545.950 84.130 2546.250 84.510 ;
        RECT 2594.710 84.510 2642.850 84.810 ;
        RECT 2545.950 83.830 2594.090 84.130 ;
        RECT 2235.910 83.450 2236.210 83.830 ;
        RECT 2414.605 83.815 2414.935 83.830 ;
        RECT 2221.190 83.150 2236.210 83.450 ;
        RECT 2317.750 83.450 2318.130 83.460 ;
        RECT 2318.925 83.450 2319.255 83.465 ;
        RECT 2317.750 83.150 2319.255 83.450 ;
        RECT 1683.205 83.135 1683.535 83.150 ;
        RECT 2027.950 83.140 2028.330 83.150 ;
        RECT 2317.750 83.140 2318.130 83.150 ;
        RECT 2318.925 83.135 2319.255 83.150 ;
        RECT 2438.985 83.450 2439.315 83.465 ;
        RECT 2463.110 83.450 2463.490 83.460 ;
        RECT 2438.985 83.150 2463.490 83.450 ;
        RECT 2593.790 83.450 2594.090 83.830 ;
        RECT 2594.710 83.450 2595.010 84.510 ;
        RECT 2642.550 84.130 2642.850 84.510 ;
        RECT 2691.310 84.510 2739.450 84.810 ;
        RECT 2642.550 83.830 2690.690 84.130 ;
        RECT 2593.790 83.150 2595.010 83.450 ;
        RECT 2690.390 83.450 2690.690 83.830 ;
        RECT 2691.310 83.450 2691.610 84.510 ;
        RECT 2739.150 84.130 2739.450 84.510 ;
        RECT 2787.910 84.510 2836.050 84.810 ;
        RECT 2739.150 83.830 2787.290 84.130 ;
        RECT 2690.390 83.150 2691.610 83.450 ;
        RECT 2786.990 83.450 2787.290 83.830 ;
        RECT 2787.910 83.450 2788.210 84.510 ;
        RECT 2835.750 84.130 2836.050 84.510 ;
        RECT 2916.710 84.130 2917.010 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
        RECT 2835.750 83.830 2883.890 84.130 ;
        RECT 2786.990 83.150 2788.210 83.450 ;
        RECT 2883.590 83.450 2883.890 83.830 ;
        RECT 2884.510 83.830 2917.010 84.130 ;
        RECT 2884.510 83.450 2884.810 83.830 ;
        RECT 2883.590 83.150 2884.810 83.450 ;
        RECT 2438.985 83.135 2439.315 83.150 ;
        RECT 2463.110 83.140 2463.490 83.150 ;
        RECT 1610.985 82.090 1611.315 82.105 ;
        RECT 1587.310 81.790 1611.315 82.090 ;
        RECT 1328.085 81.775 1328.415 81.790 ;
        RECT 1610.985 81.775 1611.315 81.790 ;
      LAYER via3 ;
        RECT 1158.580 2896.300 1158.900 2896.620 ;
        RECT 2366.540 85.860 2366.860 86.180 ;
        RECT 1158.580 83.820 1158.900 84.140 ;
        RECT 2027.060 85.180 2027.380 85.500 ;
        RECT 2027.980 83.140 2028.300 83.460 ;
        RECT 2316.860 85.180 2317.180 85.500 ;
        RECT 2366.540 84.500 2366.860 84.820 ;
        RECT 2463.140 84.500 2463.460 84.820 ;
        RECT 2317.780 83.140 2318.100 83.460 ;
        RECT 2463.140 83.140 2463.460 83.460 ;
      LAYER met4 ;
        RECT 1158.575 2896.295 1158.905 2896.625 ;
        RECT 1158.590 84.145 1158.890 2896.295 ;
        RECT 2366.535 85.855 2366.865 86.185 ;
        RECT 2027.055 85.175 2027.385 85.505 ;
        RECT 2316.855 85.175 2317.185 85.505 ;
        RECT 1158.575 83.815 1158.905 84.145 ;
        RECT 2027.070 83.450 2027.370 85.175 ;
        RECT 2027.975 83.450 2028.305 83.465 ;
        RECT 2027.070 83.150 2028.305 83.450 ;
        RECT 2316.870 83.450 2317.170 85.175 ;
        RECT 2366.550 84.825 2366.850 85.855 ;
        RECT 2366.535 84.495 2366.865 84.825 ;
        RECT 2463.135 84.495 2463.465 84.825 ;
        RECT 2463.150 83.465 2463.450 84.495 ;
        RECT 2317.775 83.450 2318.105 83.465 ;
        RECT 2316.870 83.150 2318.105 83.450 ;
        RECT 2027.975 83.135 2028.305 83.150 ;
        RECT 2317.775 83.135 2318.105 83.150 ;
        RECT 2463.135 83.135 2463.465 83.465 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1469.790 2915.315 1470.070 2915.685 ;
        RECT 1469.860 2900.000 1470.000 2915.315 ;
        RECT 1469.725 2896.000 1470.005 2900.000 ;
      LAYER via2 ;
        RECT 1469.790 2915.360 1470.070 2915.640 ;
      LAYER met3 ;
        RECT 1469.765 2915.650 1470.095 2915.665 ;
        RECT 2327.870 2915.650 2328.250 2915.660 ;
        RECT 1469.765 2915.350 2328.250 2915.650 ;
        RECT 1469.765 2915.335 1470.095 2915.350 ;
        RECT 2327.870 2915.340 2328.250 2915.350 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2916.710 2433.910 2924.800 2434.210 ;
        RECT 2329.710 2430.810 2330.090 2430.820 ;
        RECT 2329.710 2430.510 2353.050 2430.810 ;
        RECT 2329.710 2430.500 2330.090 2430.510 ;
        RECT 2352.750 2430.130 2353.050 2430.510 ;
        RECT 2401.510 2430.510 2449.650 2430.810 ;
        RECT 2352.750 2429.830 2400.890 2430.130 ;
        RECT 2400.590 2429.450 2400.890 2429.830 ;
        RECT 2401.510 2429.450 2401.810 2430.510 ;
        RECT 2449.350 2430.130 2449.650 2430.510 ;
        RECT 2498.110 2430.510 2546.250 2430.810 ;
        RECT 2449.350 2429.830 2497.490 2430.130 ;
        RECT 2400.590 2429.150 2401.810 2429.450 ;
        RECT 2497.190 2429.450 2497.490 2429.830 ;
        RECT 2498.110 2429.450 2498.410 2430.510 ;
        RECT 2545.950 2430.130 2546.250 2430.510 ;
        RECT 2594.710 2430.510 2642.850 2430.810 ;
        RECT 2545.950 2429.830 2594.090 2430.130 ;
        RECT 2497.190 2429.150 2498.410 2429.450 ;
        RECT 2593.790 2429.450 2594.090 2429.830 ;
        RECT 2594.710 2429.450 2595.010 2430.510 ;
        RECT 2642.550 2430.130 2642.850 2430.510 ;
        RECT 2691.310 2430.510 2739.450 2430.810 ;
        RECT 2642.550 2429.830 2690.690 2430.130 ;
        RECT 2593.790 2429.150 2595.010 2429.450 ;
        RECT 2690.390 2429.450 2690.690 2429.830 ;
        RECT 2691.310 2429.450 2691.610 2430.510 ;
        RECT 2739.150 2430.130 2739.450 2430.510 ;
        RECT 2787.910 2430.510 2836.050 2430.810 ;
        RECT 2739.150 2429.830 2787.290 2430.130 ;
        RECT 2690.390 2429.150 2691.610 2429.450 ;
        RECT 2786.990 2429.450 2787.290 2429.830 ;
        RECT 2787.910 2429.450 2788.210 2430.510 ;
        RECT 2835.750 2430.130 2836.050 2430.510 ;
        RECT 2916.710 2430.130 2917.010 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
        RECT 2835.750 2429.830 2883.890 2430.130 ;
        RECT 2786.990 2429.150 2788.210 2429.450 ;
        RECT 2883.590 2429.450 2883.890 2429.830 ;
        RECT 2884.510 2429.830 2917.010 2430.130 ;
        RECT 2884.510 2429.450 2884.810 2429.830 ;
        RECT 2883.590 2429.150 2884.810 2429.450 ;
      LAYER via3 ;
        RECT 2327.900 2915.340 2328.220 2915.660 ;
        RECT 2329.740 2430.500 2330.060 2430.820 ;
      LAYER met4 ;
        RECT 2327.895 2915.335 2328.225 2915.665 ;
        RECT 2327.910 2439.650 2328.210 2915.335 ;
        RECT 2327.910 2439.350 2330.050 2439.650 ;
        RECT 2329.750 2430.825 2330.050 2439.350 ;
        RECT 2329.735 2430.495 2330.065 2430.825 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1501.530 2915.995 1501.810 2916.365 ;
        RECT 1501.600 2900.000 1501.740 2915.995 ;
        RECT 1501.465 2896.000 1501.745 2900.000 ;
      LAYER via2 ;
        RECT 1501.530 2916.040 1501.810 2916.320 ;
      LAYER met3 ;
        RECT 1501.505 2916.330 1501.835 2916.345 ;
        RECT 2328.790 2916.330 2329.170 2916.340 ;
        RECT 1501.505 2916.030 2329.170 2916.330 ;
        RECT 1501.505 2916.015 1501.835 2916.030 ;
        RECT 2328.790 2916.020 2329.170 2916.030 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2916.710 2669.190 2924.800 2669.490 ;
        RECT 2328.790 2665.410 2329.170 2665.420 ;
        RECT 2328.790 2665.110 2353.050 2665.410 ;
        RECT 2328.790 2665.100 2329.170 2665.110 ;
        RECT 2352.750 2664.730 2353.050 2665.110 ;
        RECT 2401.510 2665.110 2449.650 2665.410 ;
        RECT 2352.750 2664.430 2400.890 2664.730 ;
        RECT 2400.590 2664.050 2400.890 2664.430 ;
        RECT 2401.510 2664.050 2401.810 2665.110 ;
        RECT 2449.350 2664.730 2449.650 2665.110 ;
        RECT 2498.110 2665.110 2546.250 2665.410 ;
        RECT 2449.350 2664.430 2497.490 2664.730 ;
        RECT 2400.590 2663.750 2401.810 2664.050 ;
        RECT 2497.190 2664.050 2497.490 2664.430 ;
        RECT 2498.110 2664.050 2498.410 2665.110 ;
        RECT 2545.950 2664.730 2546.250 2665.110 ;
        RECT 2594.710 2665.110 2642.850 2665.410 ;
        RECT 2545.950 2664.430 2594.090 2664.730 ;
        RECT 2497.190 2663.750 2498.410 2664.050 ;
        RECT 2593.790 2664.050 2594.090 2664.430 ;
        RECT 2594.710 2664.050 2595.010 2665.110 ;
        RECT 2642.550 2664.730 2642.850 2665.110 ;
        RECT 2691.310 2665.110 2739.450 2665.410 ;
        RECT 2642.550 2664.430 2690.690 2664.730 ;
        RECT 2593.790 2663.750 2595.010 2664.050 ;
        RECT 2690.390 2664.050 2690.690 2664.430 ;
        RECT 2691.310 2664.050 2691.610 2665.110 ;
        RECT 2739.150 2664.730 2739.450 2665.110 ;
        RECT 2787.910 2665.110 2836.050 2665.410 ;
        RECT 2739.150 2664.430 2787.290 2664.730 ;
        RECT 2690.390 2663.750 2691.610 2664.050 ;
        RECT 2786.990 2664.050 2787.290 2664.430 ;
        RECT 2787.910 2664.050 2788.210 2665.110 ;
        RECT 2835.750 2664.730 2836.050 2665.110 ;
        RECT 2916.710 2664.730 2917.010 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
        RECT 2835.750 2664.430 2883.890 2664.730 ;
        RECT 2786.990 2663.750 2788.210 2664.050 ;
        RECT 2883.590 2664.050 2883.890 2664.430 ;
        RECT 2884.510 2664.430 2917.010 2664.730 ;
        RECT 2884.510 2664.050 2884.810 2664.430 ;
        RECT 2883.590 2663.750 2884.810 2664.050 ;
      LAYER via3 ;
        RECT 2328.820 2916.020 2329.140 2916.340 ;
        RECT 2328.820 2665.100 2329.140 2665.420 ;
      LAYER met4 ;
        RECT 2328.815 2916.015 2329.145 2916.345 ;
        RECT 2328.830 2665.425 2329.130 2916.015 ;
        RECT 2328.815 2665.095 2329.145 2665.425 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1532.790 2901.120 1533.110 2901.180 ;
        RECT 2900.830 2901.120 2901.150 2901.180 ;
        RECT 1532.790 2900.980 2901.150 2901.120 ;
        RECT 1532.790 2900.920 1533.110 2900.980 ;
        RECT 2900.830 2900.920 2901.150 2900.980 ;
      LAYER via ;
        RECT 1532.820 2900.920 1533.080 2901.180 ;
        RECT 2900.860 2900.920 2901.120 2901.180 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2901.210 2901.060 2903.755 ;
        RECT 1532.820 2900.890 1533.080 2901.210 ;
        RECT 2900.860 2900.890 2901.120 2901.210 ;
        RECT 1532.880 2900.000 1533.020 2900.890 ;
        RECT 1532.745 2896.000 1533.025 2900.000 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1565.910 3133.000 1566.230 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 1565.910 3132.860 2901.150 3133.000 ;
        RECT 1565.910 3132.800 1566.230 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
      LAYER via ;
        RECT 1565.940 3132.800 1566.200 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 1565.940 3132.770 1566.200 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 1564.485 2899.930 1564.765 2900.000 ;
        RECT 1566.000 2899.930 1566.140 3132.770 ;
        RECT 1564.485 2899.790 1566.140 2899.930 ;
        RECT 1564.485 2896.000 1564.765 2899.790 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1600.410 3367.600 1600.730 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 1600.410 3367.460 2901.150 3367.600 ;
        RECT 1600.410 3367.400 1600.730 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
      LAYER via ;
        RECT 1600.440 3367.400 1600.700 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 1600.440 3367.370 1600.700 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 1600.500 2900.610 1600.640 3367.370 ;
        RECT 1598.660 2900.470 1600.640 2900.610 ;
        RECT 1596.225 2899.250 1596.505 2900.000 ;
        RECT 1598.660 2899.250 1598.800 2900.470 ;
        RECT 1596.225 2899.110 1598.800 2899.250 ;
        RECT 1596.225 2896.000 1596.505 2899.110 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2796.485 3332.765 2796.655 3422.355 ;
        RECT 2795.565 3008.405 2795.735 3042.915 ;
        RECT 2796.485 2946.525 2796.655 2994.635 ;
      LAYER mcon ;
        RECT 2796.485 3422.185 2796.655 3422.355 ;
        RECT 2795.565 3042.745 2795.735 3042.915 ;
        RECT 2796.485 2994.465 2796.655 2994.635 ;
      LAYER met1 ;
        RECT 2795.490 3443.080 2795.810 3443.140 ;
        RECT 2798.250 3443.080 2798.570 3443.140 ;
        RECT 2795.490 3442.940 2798.570 3443.080 ;
        RECT 2795.490 3442.880 2795.810 3442.940 ;
        RECT 2798.250 3442.880 2798.570 3442.940 ;
        RECT 2795.030 3422.340 2795.350 3422.400 ;
        RECT 2796.425 3422.340 2796.715 3422.385 ;
        RECT 2795.030 3422.200 2796.715 3422.340 ;
        RECT 2795.030 3422.140 2795.350 3422.200 ;
        RECT 2796.425 3422.155 2796.715 3422.200 ;
        RECT 2796.425 3332.920 2796.715 3332.965 ;
        RECT 2796.870 3332.920 2797.190 3332.980 ;
        RECT 2796.425 3332.780 2797.190 3332.920 ;
        RECT 2796.425 3332.735 2796.715 3332.780 ;
        RECT 2796.870 3332.720 2797.190 3332.780 ;
        RECT 2795.490 3236.360 2795.810 3236.420 ;
        RECT 2795.950 3236.360 2796.270 3236.420 ;
        RECT 2795.490 3236.220 2796.270 3236.360 ;
        RECT 2795.490 3236.160 2795.810 3236.220 ;
        RECT 2795.950 3236.160 2796.270 3236.220 ;
        RECT 2795.490 3202.020 2795.810 3202.080 ;
        RECT 2795.950 3202.020 2796.270 3202.080 ;
        RECT 2795.490 3201.880 2796.270 3202.020 ;
        RECT 2795.490 3201.820 2795.810 3201.880 ;
        RECT 2795.950 3201.820 2796.270 3201.880 ;
        RECT 2795.030 3153.400 2795.350 3153.460 ;
        RECT 2795.950 3153.400 2796.270 3153.460 ;
        RECT 2795.030 3153.260 2796.270 3153.400 ;
        RECT 2795.030 3153.200 2795.350 3153.260 ;
        RECT 2795.950 3153.200 2796.270 3153.260 ;
        RECT 2795.030 3056.840 2795.350 3056.900 ;
        RECT 2795.950 3056.840 2796.270 3056.900 ;
        RECT 2795.030 3056.700 2796.270 3056.840 ;
        RECT 2795.030 3056.640 2795.350 3056.700 ;
        RECT 2795.950 3056.640 2796.270 3056.700 ;
        RECT 2795.490 3042.900 2795.810 3042.960 ;
        RECT 2795.295 3042.760 2795.810 3042.900 ;
        RECT 2795.490 3042.700 2795.810 3042.760 ;
        RECT 2795.505 3008.560 2795.795 3008.605 ;
        RECT 2796.410 3008.560 2796.730 3008.620 ;
        RECT 2795.505 3008.420 2796.730 3008.560 ;
        RECT 2795.505 3008.375 2795.795 3008.420 ;
        RECT 2796.410 3008.360 2796.730 3008.420 ;
        RECT 2796.410 2994.620 2796.730 2994.680 ;
        RECT 2796.215 2994.480 2796.730 2994.620 ;
        RECT 2796.410 2994.420 2796.730 2994.480 ;
        RECT 2796.425 2946.680 2796.715 2946.725 ;
        RECT 2796.870 2946.680 2797.190 2946.740 ;
        RECT 2796.425 2946.540 2797.190 2946.680 ;
        RECT 2796.425 2946.495 2796.715 2946.540 ;
        RECT 2796.870 2946.480 2797.190 2946.540 ;
        RECT 1627.550 2922.200 1627.870 2922.260 ;
        RECT 2796.870 2922.200 2797.190 2922.260 ;
        RECT 1627.550 2922.060 2797.190 2922.200 ;
        RECT 1627.550 2922.000 1627.870 2922.060 ;
        RECT 2796.870 2922.000 2797.190 2922.060 ;
      LAYER via ;
        RECT 2795.520 3442.880 2795.780 3443.140 ;
        RECT 2798.280 3442.880 2798.540 3443.140 ;
        RECT 2795.060 3422.140 2795.320 3422.400 ;
        RECT 2796.900 3332.720 2797.160 3332.980 ;
        RECT 2795.520 3236.160 2795.780 3236.420 ;
        RECT 2795.980 3236.160 2796.240 3236.420 ;
        RECT 2795.520 3201.820 2795.780 3202.080 ;
        RECT 2795.980 3201.820 2796.240 3202.080 ;
        RECT 2795.060 3153.200 2795.320 3153.460 ;
        RECT 2795.980 3153.200 2796.240 3153.460 ;
        RECT 2795.060 3056.640 2795.320 3056.900 ;
        RECT 2795.980 3056.640 2796.240 3056.900 ;
        RECT 2795.520 3042.700 2795.780 3042.960 ;
        RECT 2796.440 3008.360 2796.700 3008.620 ;
        RECT 2796.440 2994.420 2796.700 2994.680 ;
        RECT 2796.900 2946.480 2797.160 2946.740 ;
        RECT 1627.580 2922.000 1627.840 2922.260 ;
        RECT 2796.900 2922.000 2797.160 2922.260 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3443.170 2798.480 3517.600 ;
        RECT 2795.520 3442.850 2795.780 3443.170 ;
        RECT 2798.280 3442.850 2798.540 3443.170 ;
        RECT 2795.580 3429.650 2795.720 3442.850 ;
        RECT 2795.120 3429.510 2795.720 3429.650 ;
        RECT 2795.120 3422.430 2795.260 3429.510 ;
        RECT 2795.060 3422.110 2795.320 3422.430 ;
        RECT 2796.900 3332.690 2797.160 3333.010 ;
        RECT 2796.960 3298.410 2797.100 3332.690 ;
        RECT 2796.040 3298.270 2797.100 3298.410 ;
        RECT 2796.040 3236.450 2796.180 3298.270 ;
        RECT 2795.520 3236.130 2795.780 3236.450 ;
        RECT 2795.980 3236.130 2796.240 3236.450 ;
        RECT 2795.580 3202.110 2795.720 3236.130 ;
        RECT 2795.520 3201.790 2795.780 3202.110 ;
        RECT 2795.980 3201.790 2796.240 3202.110 ;
        RECT 2796.040 3153.490 2796.180 3201.790 ;
        RECT 2795.060 3153.170 2795.320 3153.490 ;
        RECT 2795.980 3153.170 2796.240 3153.490 ;
        RECT 2795.120 3152.890 2795.260 3153.170 ;
        RECT 2795.120 3152.750 2795.720 3152.890 ;
        RECT 2795.580 3105.290 2795.720 3152.750 ;
        RECT 2795.580 3105.150 2796.180 3105.290 ;
        RECT 2796.040 3056.930 2796.180 3105.150 ;
        RECT 2795.060 3056.610 2795.320 3056.930 ;
        RECT 2795.980 3056.610 2796.240 3056.930 ;
        RECT 2795.120 3056.330 2795.260 3056.610 ;
        RECT 2795.120 3056.190 2795.720 3056.330 ;
        RECT 2795.580 3042.990 2795.720 3056.190 ;
        RECT 2795.520 3042.670 2795.780 3042.990 ;
        RECT 2796.440 3008.330 2796.700 3008.650 ;
        RECT 2796.500 2994.710 2796.640 3008.330 ;
        RECT 2796.440 2994.390 2796.700 2994.710 ;
        RECT 2796.900 2946.450 2797.160 2946.770 ;
        RECT 2796.960 2922.290 2797.100 2946.450 ;
        RECT 1627.580 2921.970 1627.840 2922.290 ;
        RECT 2796.900 2921.970 2797.160 2922.290 ;
        RECT 1627.640 2900.000 1627.780 2921.970 ;
        RECT 1627.505 2896.000 1627.785 2900.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2470.345 3332.765 2470.515 3380.875 ;
      LAYER mcon ;
        RECT 2470.345 3380.705 2470.515 3380.875 ;
      LAYER met1 ;
        RECT 2470.270 3380.860 2470.590 3380.920 ;
        RECT 2470.075 3380.720 2470.590 3380.860 ;
        RECT 2470.270 3380.660 2470.590 3380.720 ;
        RECT 2470.285 3332.920 2470.575 3332.965 ;
        RECT 2470.730 3332.920 2471.050 3332.980 ;
        RECT 2470.285 3332.780 2471.050 3332.920 ;
        RECT 2470.285 3332.735 2470.575 3332.780 ;
        RECT 2470.730 3332.720 2471.050 3332.780 ;
        RECT 2470.270 3270.700 2470.590 3270.760 ;
        RECT 2471.190 3270.700 2471.510 3270.760 ;
        RECT 2470.270 3270.560 2471.510 3270.700 ;
        RECT 2470.270 3270.500 2470.590 3270.560 ;
        RECT 2471.190 3270.500 2471.510 3270.560 ;
        RECT 2470.270 3174.140 2470.590 3174.200 ;
        RECT 2471.190 3174.140 2471.510 3174.200 ;
        RECT 2470.270 3174.000 2471.510 3174.140 ;
        RECT 2470.270 3173.940 2470.590 3174.000 ;
        RECT 2471.190 3173.940 2471.510 3174.000 ;
        RECT 2470.270 3077.580 2470.590 3077.640 ;
        RECT 2471.190 3077.580 2471.510 3077.640 ;
        RECT 2470.270 3077.440 2471.510 3077.580 ;
        RECT 2470.270 3077.380 2470.590 3077.440 ;
        RECT 2471.190 3077.380 2471.510 3077.440 ;
        RECT 2470.270 2981.020 2470.590 2981.080 ;
        RECT 2471.190 2981.020 2471.510 2981.080 ;
        RECT 2470.270 2980.880 2471.510 2981.020 ;
        RECT 2470.270 2980.820 2470.590 2980.880 ;
        RECT 2471.190 2980.820 2471.510 2980.880 ;
        RECT 1659.290 2922.540 1659.610 2922.600 ;
        RECT 2471.190 2922.540 2471.510 2922.600 ;
        RECT 1659.290 2922.400 2471.510 2922.540 ;
        RECT 1659.290 2922.340 1659.610 2922.400 ;
        RECT 2471.190 2922.340 2471.510 2922.400 ;
      LAYER via ;
        RECT 2470.300 3380.660 2470.560 3380.920 ;
        RECT 2470.760 3332.720 2471.020 3332.980 ;
        RECT 2470.300 3270.500 2470.560 3270.760 ;
        RECT 2471.220 3270.500 2471.480 3270.760 ;
        RECT 2470.300 3173.940 2470.560 3174.200 ;
        RECT 2471.220 3173.940 2471.480 3174.200 ;
        RECT 2470.300 3077.380 2470.560 3077.640 ;
        RECT 2471.220 3077.380 2471.480 3077.640 ;
        RECT 2470.300 2980.820 2470.560 2981.080 ;
        RECT 2471.220 2980.820 2471.480 2981.080 ;
        RECT 1659.320 2922.340 1659.580 2922.600 ;
        RECT 2471.220 2922.340 2471.480 2922.600 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3517.370 2474.180 3517.600 ;
        RECT 2474.040 3517.230 2474.640 3517.370 ;
        RECT 2474.500 3430.445 2474.640 3517.230 ;
        RECT 2474.430 3430.075 2474.710 3430.445 ;
        RECT 2471.210 3429.395 2471.490 3429.765 ;
        RECT 2471.280 3394.970 2471.420 3429.395 ;
        RECT 2470.360 3394.830 2471.420 3394.970 ;
        RECT 2470.360 3380.950 2470.500 3394.830 ;
        RECT 2470.300 3380.630 2470.560 3380.950 ;
        RECT 2470.760 3332.690 2471.020 3333.010 ;
        RECT 2470.820 3298.410 2470.960 3332.690 ;
        RECT 2470.820 3298.270 2471.420 3298.410 ;
        RECT 2471.280 3270.790 2471.420 3298.270 ;
        RECT 2470.300 3270.470 2470.560 3270.790 ;
        RECT 2471.220 3270.470 2471.480 3270.790 ;
        RECT 2470.360 3222.250 2470.500 3270.470 ;
        RECT 2470.360 3222.110 2471.420 3222.250 ;
        RECT 2471.280 3174.230 2471.420 3222.110 ;
        RECT 2470.300 3173.910 2470.560 3174.230 ;
        RECT 2471.220 3173.910 2471.480 3174.230 ;
        RECT 2470.360 3125.690 2470.500 3173.910 ;
        RECT 2470.360 3125.550 2471.420 3125.690 ;
        RECT 2471.280 3077.670 2471.420 3125.550 ;
        RECT 2470.300 3077.350 2470.560 3077.670 ;
        RECT 2471.220 3077.350 2471.480 3077.670 ;
        RECT 2470.360 3029.130 2470.500 3077.350 ;
        RECT 2470.360 3028.990 2471.420 3029.130 ;
        RECT 2471.280 2981.110 2471.420 3028.990 ;
        RECT 2470.300 2980.850 2470.560 2981.110 ;
        RECT 2470.300 2980.790 2470.960 2980.850 ;
        RECT 2471.220 2980.790 2471.480 2981.110 ;
        RECT 2470.360 2980.710 2470.960 2980.790 ;
        RECT 2470.820 2980.170 2470.960 2980.710 ;
        RECT 2470.820 2980.030 2471.420 2980.170 ;
        RECT 2471.280 2922.630 2471.420 2980.030 ;
        RECT 1659.320 2922.310 1659.580 2922.630 ;
        RECT 2471.220 2922.310 2471.480 2922.630 ;
        RECT 1659.380 2900.000 1659.520 2922.310 ;
        RECT 1659.245 2896.000 1659.525 2900.000 ;
      LAYER via2 ;
        RECT 2474.430 3430.120 2474.710 3430.400 ;
        RECT 2471.210 3429.440 2471.490 3429.720 ;
      LAYER met3 ;
        RECT 2474.405 3430.410 2474.735 3430.425 ;
        RECT 2470.510 3430.110 2474.735 3430.410 ;
        RECT 2470.510 3429.730 2470.810 3430.110 ;
        RECT 2474.405 3430.095 2474.735 3430.110 ;
        RECT 2471.185 3429.730 2471.515 3429.745 ;
        RECT 2470.510 3429.430 2471.515 3429.730 ;
        RECT 2471.185 3429.415 2471.515 3429.430 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2147.885 3332.765 2148.055 3422.355 ;
        RECT 2146.965 3008.405 2147.135 3042.915 ;
        RECT 2147.885 2946.525 2148.055 2994.635 ;
      LAYER mcon ;
        RECT 2147.885 3422.185 2148.055 3422.355 ;
        RECT 2146.965 3042.745 2147.135 3042.915 ;
        RECT 2147.885 2994.465 2148.055 2994.635 ;
      LAYER met1 ;
        RECT 2146.890 3443.080 2147.210 3443.140 ;
        RECT 2149.190 3443.080 2149.510 3443.140 ;
        RECT 2146.890 3442.940 2149.510 3443.080 ;
        RECT 2146.890 3442.880 2147.210 3442.940 ;
        RECT 2149.190 3442.880 2149.510 3442.940 ;
        RECT 2146.430 3422.340 2146.750 3422.400 ;
        RECT 2147.825 3422.340 2148.115 3422.385 ;
        RECT 2146.430 3422.200 2148.115 3422.340 ;
        RECT 2146.430 3422.140 2146.750 3422.200 ;
        RECT 2147.825 3422.155 2148.115 3422.200 ;
        RECT 2147.825 3332.920 2148.115 3332.965 ;
        RECT 2148.270 3332.920 2148.590 3332.980 ;
        RECT 2147.825 3332.780 2148.590 3332.920 ;
        RECT 2147.825 3332.735 2148.115 3332.780 ;
        RECT 2148.270 3332.720 2148.590 3332.780 ;
        RECT 2146.890 3236.360 2147.210 3236.420 ;
        RECT 2147.350 3236.360 2147.670 3236.420 ;
        RECT 2146.890 3236.220 2147.670 3236.360 ;
        RECT 2146.890 3236.160 2147.210 3236.220 ;
        RECT 2147.350 3236.160 2147.670 3236.220 ;
        RECT 2146.890 3202.020 2147.210 3202.080 ;
        RECT 2147.350 3202.020 2147.670 3202.080 ;
        RECT 2146.890 3201.880 2147.670 3202.020 ;
        RECT 2146.890 3201.820 2147.210 3201.880 ;
        RECT 2147.350 3201.820 2147.670 3201.880 ;
        RECT 2146.430 3153.400 2146.750 3153.460 ;
        RECT 2147.350 3153.400 2147.670 3153.460 ;
        RECT 2146.430 3153.260 2147.670 3153.400 ;
        RECT 2146.430 3153.200 2146.750 3153.260 ;
        RECT 2147.350 3153.200 2147.670 3153.260 ;
        RECT 2146.430 3056.840 2146.750 3056.900 ;
        RECT 2147.350 3056.840 2147.670 3056.900 ;
        RECT 2146.430 3056.700 2147.670 3056.840 ;
        RECT 2146.430 3056.640 2146.750 3056.700 ;
        RECT 2147.350 3056.640 2147.670 3056.700 ;
        RECT 2146.890 3042.900 2147.210 3042.960 ;
        RECT 2146.695 3042.760 2147.210 3042.900 ;
        RECT 2146.890 3042.700 2147.210 3042.760 ;
        RECT 2146.905 3008.560 2147.195 3008.605 ;
        RECT 2147.810 3008.560 2148.130 3008.620 ;
        RECT 2146.905 3008.420 2148.130 3008.560 ;
        RECT 2146.905 3008.375 2147.195 3008.420 ;
        RECT 2147.810 3008.360 2148.130 3008.420 ;
        RECT 2147.810 2994.620 2148.130 2994.680 ;
        RECT 2147.615 2994.480 2148.130 2994.620 ;
        RECT 2147.810 2994.420 2148.130 2994.480 ;
        RECT 2147.825 2946.680 2148.115 2946.725 ;
        RECT 2148.270 2946.680 2148.590 2946.740 ;
        RECT 2147.825 2946.540 2148.590 2946.680 ;
        RECT 2147.825 2946.495 2148.115 2946.540 ;
        RECT 2148.270 2946.480 2148.590 2946.540 ;
        RECT 1691.030 2922.880 1691.350 2922.940 ;
        RECT 2148.270 2922.880 2148.590 2922.940 ;
        RECT 1691.030 2922.740 2148.590 2922.880 ;
        RECT 1691.030 2922.680 1691.350 2922.740 ;
        RECT 2148.270 2922.680 2148.590 2922.740 ;
      LAYER via ;
        RECT 2146.920 3442.880 2147.180 3443.140 ;
        RECT 2149.220 3442.880 2149.480 3443.140 ;
        RECT 2146.460 3422.140 2146.720 3422.400 ;
        RECT 2148.300 3332.720 2148.560 3332.980 ;
        RECT 2146.920 3236.160 2147.180 3236.420 ;
        RECT 2147.380 3236.160 2147.640 3236.420 ;
        RECT 2146.920 3201.820 2147.180 3202.080 ;
        RECT 2147.380 3201.820 2147.640 3202.080 ;
        RECT 2146.460 3153.200 2146.720 3153.460 ;
        RECT 2147.380 3153.200 2147.640 3153.460 ;
        RECT 2146.460 3056.640 2146.720 3056.900 ;
        RECT 2147.380 3056.640 2147.640 3056.900 ;
        RECT 2146.920 3042.700 2147.180 3042.960 ;
        RECT 2147.840 3008.360 2148.100 3008.620 ;
        RECT 2147.840 2994.420 2148.100 2994.680 ;
        RECT 2148.300 2946.480 2148.560 2946.740 ;
        RECT 1691.060 2922.680 1691.320 2922.940 ;
        RECT 2148.300 2922.680 2148.560 2922.940 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3443.170 2149.420 3517.600 ;
        RECT 2146.920 3442.850 2147.180 3443.170 ;
        RECT 2149.220 3442.850 2149.480 3443.170 ;
        RECT 2146.980 3429.650 2147.120 3442.850 ;
        RECT 2146.520 3429.510 2147.120 3429.650 ;
        RECT 2146.520 3422.430 2146.660 3429.510 ;
        RECT 2146.460 3422.110 2146.720 3422.430 ;
        RECT 2148.300 3332.690 2148.560 3333.010 ;
        RECT 2148.360 3298.410 2148.500 3332.690 ;
        RECT 2147.440 3298.270 2148.500 3298.410 ;
        RECT 2147.440 3236.450 2147.580 3298.270 ;
        RECT 2146.920 3236.130 2147.180 3236.450 ;
        RECT 2147.380 3236.130 2147.640 3236.450 ;
        RECT 2146.980 3202.110 2147.120 3236.130 ;
        RECT 2146.920 3201.790 2147.180 3202.110 ;
        RECT 2147.380 3201.790 2147.640 3202.110 ;
        RECT 2147.440 3153.490 2147.580 3201.790 ;
        RECT 2146.460 3153.170 2146.720 3153.490 ;
        RECT 2147.380 3153.170 2147.640 3153.490 ;
        RECT 2146.520 3152.890 2146.660 3153.170 ;
        RECT 2146.520 3152.750 2147.120 3152.890 ;
        RECT 2146.980 3105.290 2147.120 3152.750 ;
        RECT 2146.980 3105.150 2147.580 3105.290 ;
        RECT 2147.440 3056.930 2147.580 3105.150 ;
        RECT 2146.460 3056.610 2146.720 3056.930 ;
        RECT 2147.380 3056.610 2147.640 3056.930 ;
        RECT 2146.520 3056.330 2146.660 3056.610 ;
        RECT 2146.520 3056.190 2147.120 3056.330 ;
        RECT 2146.980 3042.990 2147.120 3056.190 ;
        RECT 2146.920 3042.670 2147.180 3042.990 ;
        RECT 2147.840 3008.330 2148.100 3008.650 ;
        RECT 2147.900 2994.710 2148.040 3008.330 ;
        RECT 2147.840 2994.390 2148.100 2994.710 ;
        RECT 2148.300 2946.450 2148.560 2946.770 ;
        RECT 2148.360 2922.970 2148.500 2946.450 ;
        RECT 1691.060 2922.650 1691.320 2922.970 ;
        RECT 2148.300 2922.650 2148.560 2922.970 ;
        RECT 1691.120 2900.000 1691.260 2922.650 ;
        RECT 1690.985 2896.000 1691.265 2900.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1822.665 3381.045 1822.835 3429.155 ;
        RECT 1822.665 3043.085 1822.835 3091.195 ;
        RECT 1823.125 2946.525 1823.295 2994.635 ;
      LAYER mcon ;
        RECT 1822.665 3428.985 1822.835 3429.155 ;
        RECT 1822.665 3091.025 1822.835 3091.195 ;
        RECT 1823.125 2994.465 1823.295 2994.635 ;
      LAYER met1 ;
        RECT 1823.050 3439.000 1823.370 3439.060 ;
        RECT 1825.810 3439.000 1826.130 3439.060 ;
        RECT 1823.050 3438.860 1826.130 3439.000 ;
        RECT 1823.050 3438.800 1823.370 3438.860 ;
        RECT 1825.810 3438.800 1826.130 3438.860 ;
        RECT 1822.605 3429.140 1822.895 3429.185 ;
        RECT 1823.050 3429.140 1823.370 3429.200 ;
        RECT 1822.605 3429.000 1823.370 3429.140 ;
        RECT 1822.605 3428.955 1822.895 3429.000 ;
        RECT 1823.050 3428.940 1823.370 3429.000 ;
        RECT 1822.590 3381.200 1822.910 3381.260 ;
        RECT 1822.395 3381.060 1822.910 3381.200 ;
        RECT 1822.590 3381.000 1822.910 3381.060 ;
        RECT 1822.605 3091.180 1822.895 3091.225 ;
        RECT 1823.050 3091.180 1823.370 3091.240 ;
        RECT 1822.605 3091.040 1823.370 3091.180 ;
        RECT 1822.605 3090.995 1822.895 3091.040 ;
        RECT 1823.050 3090.980 1823.370 3091.040 ;
        RECT 1822.590 3043.240 1822.910 3043.300 ;
        RECT 1822.395 3043.100 1822.910 3043.240 ;
        RECT 1822.590 3043.040 1822.910 3043.100 ;
        RECT 1823.050 2994.620 1823.370 2994.680 ;
        RECT 1822.855 2994.480 1823.370 2994.620 ;
        RECT 1823.050 2994.420 1823.370 2994.480 ;
        RECT 1823.065 2946.680 1823.355 2946.725 ;
        RECT 1823.510 2946.680 1823.830 2946.740 ;
        RECT 1823.065 2946.540 1823.830 2946.680 ;
        RECT 1823.065 2946.495 1823.355 2946.540 ;
        RECT 1823.510 2946.480 1823.830 2946.540 ;
        RECT 1722.310 2923.560 1722.630 2923.620 ;
        RECT 1823.510 2923.560 1823.830 2923.620 ;
        RECT 1722.310 2923.420 1823.830 2923.560 ;
        RECT 1722.310 2923.360 1722.630 2923.420 ;
        RECT 1823.510 2923.360 1823.830 2923.420 ;
      LAYER via ;
        RECT 1823.080 3438.800 1823.340 3439.060 ;
        RECT 1825.840 3438.800 1826.100 3439.060 ;
        RECT 1823.080 3428.940 1823.340 3429.200 ;
        RECT 1822.620 3381.000 1822.880 3381.260 ;
        RECT 1823.080 3090.980 1823.340 3091.240 ;
        RECT 1822.620 3043.040 1822.880 3043.300 ;
        RECT 1823.080 2994.420 1823.340 2994.680 ;
        RECT 1823.540 2946.480 1823.800 2946.740 ;
        RECT 1722.340 2923.360 1722.600 2923.620 ;
        RECT 1823.540 2923.360 1823.800 2923.620 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3517.370 1825.120 3517.600 ;
        RECT 1824.980 3517.230 1826.040 3517.370 ;
        RECT 1825.900 3439.090 1826.040 3517.230 ;
        RECT 1823.080 3438.770 1823.340 3439.090 ;
        RECT 1825.840 3438.770 1826.100 3439.090 ;
        RECT 1823.140 3429.230 1823.280 3438.770 ;
        RECT 1823.080 3428.910 1823.340 3429.230 ;
        RECT 1822.620 3380.970 1822.880 3381.290 ;
        RECT 1822.680 3346.690 1822.820 3380.970 ;
        RECT 1822.680 3346.550 1823.740 3346.690 ;
        RECT 1823.600 3250.130 1823.740 3346.550 ;
        RECT 1822.680 3249.990 1823.740 3250.130 ;
        RECT 1822.680 3153.570 1822.820 3249.990 ;
        RECT 1822.680 3153.430 1823.280 3153.570 ;
        RECT 1823.140 3091.270 1823.280 3153.430 ;
        RECT 1823.080 3090.950 1823.340 3091.270 ;
        RECT 1822.620 3043.010 1822.880 3043.330 ;
        RECT 1822.680 3008.730 1822.820 3043.010 ;
        RECT 1822.680 3008.590 1823.280 3008.730 ;
        RECT 1823.140 2994.710 1823.280 3008.590 ;
        RECT 1823.080 2994.390 1823.340 2994.710 ;
        RECT 1823.540 2946.450 1823.800 2946.770 ;
        RECT 1823.600 2923.650 1823.740 2946.450 ;
        RECT 1722.340 2923.330 1722.600 2923.650 ;
        RECT 1823.540 2923.330 1823.800 2923.650 ;
        RECT 1722.400 2900.000 1722.540 2923.330 ;
        RECT 1722.265 2896.000 1722.545 2900.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1500.590 3498.500 1500.910 3498.560 ;
        RECT 1503.810 3498.500 1504.130 3498.560 ;
        RECT 1500.590 3498.360 1504.130 3498.500 ;
        RECT 1500.590 3498.300 1500.910 3498.360 ;
        RECT 1503.810 3498.300 1504.130 3498.360 ;
        RECT 1503.810 2923.220 1504.130 2923.280 ;
        RECT 1754.050 2923.220 1754.370 2923.280 ;
        RECT 1503.810 2923.080 1754.370 2923.220 ;
        RECT 1503.810 2923.020 1504.130 2923.080 ;
        RECT 1754.050 2923.020 1754.370 2923.080 ;
      LAYER via ;
        RECT 1500.620 3498.300 1500.880 3498.560 ;
        RECT 1503.840 3498.300 1504.100 3498.560 ;
        RECT 1503.840 2923.020 1504.100 2923.280 ;
        RECT 1754.080 2923.020 1754.340 2923.280 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3498.590 1500.820 3517.600 ;
        RECT 1500.620 3498.270 1500.880 3498.590 ;
        RECT 1503.840 3498.270 1504.100 3498.590 ;
        RECT 1503.900 2923.310 1504.040 3498.270 ;
        RECT 1503.840 2922.990 1504.100 2923.310 ;
        RECT 1754.080 2922.990 1754.340 2923.310 ;
        RECT 1754.140 2900.000 1754.280 2922.990 ;
        RECT 1754.005 2896.000 1754.285 2900.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1891.130 319.500 1891.450 319.560 ;
        RECT 1931.610 319.500 1931.930 319.560 ;
        RECT 1891.130 319.360 1931.930 319.500 ;
        RECT 1891.130 319.300 1891.450 319.360 ;
        RECT 1931.610 319.300 1931.930 319.360 ;
        RECT 2089.390 318.480 2089.710 318.540 ;
        RECT 2090.770 318.480 2091.090 318.540 ;
        RECT 2089.390 318.340 2091.090 318.480 ;
        RECT 2089.390 318.280 2089.710 318.340 ;
        RECT 2090.770 318.280 2091.090 318.340 ;
        RECT 2185.990 318.480 2186.310 318.540 ;
        RECT 2187.370 318.480 2187.690 318.540 ;
        RECT 2185.990 318.340 2187.690 318.480 ;
        RECT 2185.990 318.280 2186.310 318.340 ;
        RECT 2187.370 318.280 2187.690 318.340 ;
        RECT 2282.590 318.480 2282.910 318.540 ;
        RECT 2284.430 318.480 2284.750 318.540 ;
        RECT 2282.590 318.340 2284.750 318.480 ;
        RECT 2282.590 318.280 2282.910 318.340 ;
        RECT 2284.430 318.280 2284.750 318.340 ;
      LAYER via ;
        RECT 1891.160 319.300 1891.420 319.560 ;
        RECT 1931.640 319.300 1931.900 319.560 ;
        RECT 2089.420 318.280 2089.680 318.540 ;
        RECT 2090.800 318.280 2091.060 318.540 ;
        RECT 2186.020 318.280 2186.280 318.540 ;
        RECT 2187.400 318.280 2187.660 318.540 ;
        RECT 2282.620 318.280 2282.880 318.540 ;
        RECT 2284.460 318.280 2284.720 318.540 ;
      LAYER met2 ;
        RECT 1185.445 2896.530 1185.725 2900.000 ;
        RECT 1185.970 2896.530 1186.250 2896.645 ;
        RECT 1185.445 2896.390 1186.250 2896.530 ;
        RECT 1185.445 2896.000 1185.725 2896.390 ;
        RECT 1185.970 2896.275 1186.250 2896.390 ;
        RECT 1891.160 319.445 1891.420 319.590 ;
        RECT 1931.640 319.445 1931.900 319.590 ;
        RECT 1891.150 319.075 1891.430 319.445 ;
        RECT 1931.630 319.075 1931.910 319.445 ;
        RECT 1800.530 318.650 1800.810 318.765 ;
        RECT 1801.450 318.650 1801.730 318.765 ;
        RECT 1800.530 318.510 1801.730 318.650 ;
        RECT 1800.530 318.395 1800.810 318.510 ;
        RECT 1801.450 318.395 1801.730 318.510 ;
        RECT 2089.410 318.395 2089.690 318.765 ;
        RECT 2090.790 318.395 2091.070 318.765 ;
        RECT 2186.010 318.395 2186.290 318.765 ;
        RECT 2187.390 318.395 2187.670 318.765 ;
        RECT 2282.610 318.395 2282.890 318.765 ;
        RECT 2284.450 318.395 2284.730 318.765 ;
        RECT 2089.420 318.250 2089.680 318.395 ;
        RECT 2090.800 318.250 2091.060 318.395 ;
        RECT 2186.020 318.250 2186.280 318.395 ;
        RECT 2187.400 318.250 2187.660 318.395 ;
        RECT 2282.620 318.250 2282.880 318.395 ;
        RECT 2284.460 318.250 2284.720 318.395 ;
      LAYER via2 ;
        RECT 1185.970 2896.320 1186.250 2896.600 ;
        RECT 1891.150 319.120 1891.430 319.400 ;
        RECT 1931.630 319.120 1931.910 319.400 ;
        RECT 1800.530 318.440 1800.810 318.720 ;
        RECT 1801.450 318.440 1801.730 318.720 ;
        RECT 2089.410 318.440 2089.690 318.720 ;
        RECT 2090.790 318.440 2091.070 318.720 ;
        RECT 2186.010 318.440 2186.290 318.720 ;
        RECT 2187.390 318.440 2187.670 318.720 ;
        RECT 2282.610 318.440 2282.890 318.720 ;
        RECT 2284.450 318.440 2284.730 318.720 ;
      LAYER met3 ;
        RECT 1185.945 2896.620 1186.275 2896.625 ;
        RECT 1185.945 2896.610 1186.530 2896.620 ;
        RECT 1185.945 2896.310 1186.730 2896.610 ;
        RECT 1185.945 2896.300 1186.530 2896.310 ;
        RECT 1185.945 2896.295 1186.275 2896.300 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2916.710 322.510 2924.800 322.810 ;
        RECT 1586.350 320.090 1586.730 320.100 ;
        RECT 2027.030 320.090 2027.410 320.100 ;
        RECT 1538.550 319.790 1586.730 320.090 ;
        RECT 1400.510 319.410 1400.890 319.420 ;
        RECT 1376.630 319.110 1400.890 319.410 ;
        RECT 1186.150 318.730 1186.530 318.740 ;
        RECT 1186.150 318.430 1280.330 318.730 ;
        RECT 1186.150 318.420 1186.530 318.430 ;
        RECT 1280.030 318.050 1280.330 318.430 ;
        RECT 1376.630 318.050 1376.930 319.110 ;
        RECT 1400.510 319.100 1400.890 319.110 ;
        RECT 1442.830 318.730 1443.210 318.740 ;
        RECT 1538.550 318.730 1538.850 319.790 ;
        RECT 1586.350 319.780 1586.730 319.790 ;
        RECT 1993.030 319.790 2027.410 320.090 ;
        RECT 1635.110 319.410 1635.490 319.420 ;
        RECT 1891.125 319.410 1891.455 319.425 ;
        RECT 1635.110 319.110 1704.450 319.410 ;
        RECT 1635.110 319.100 1635.490 319.110 ;
        RECT 1442.830 318.430 1538.850 318.730 ;
        RECT 1442.830 318.420 1443.210 318.430 ;
        RECT 1280.030 317.750 1376.930 318.050 ;
        RECT 1400.510 318.050 1400.890 318.060 ;
        RECT 1441.910 318.050 1442.290 318.060 ;
        RECT 1400.510 317.750 1442.290 318.050 ;
        RECT 1400.510 317.740 1400.890 317.750 ;
        RECT 1441.910 317.740 1442.290 317.750 ;
        RECT 1586.350 318.050 1586.730 318.060 ;
        RECT 1635.110 318.050 1635.490 318.060 ;
        RECT 1586.350 317.750 1635.490 318.050 ;
        RECT 1704.150 318.050 1704.450 319.110 ;
        RECT 1849.510 319.110 1891.455 319.410 ;
        RECT 1800.505 318.730 1800.835 318.745 ;
        RECT 1752.910 318.430 1800.835 318.730 ;
        RECT 1752.910 318.050 1753.210 318.430 ;
        RECT 1800.505 318.415 1800.835 318.430 ;
        RECT 1801.425 318.730 1801.755 318.745 ;
        RECT 1801.425 318.430 1848.890 318.730 ;
        RECT 1801.425 318.415 1801.755 318.430 ;
        RECT 1704.150 317.750 1753.210 318.050 ;
        RECT 1848.590 318.050 1848.890 318.430 ;
        RECT 1849.510 318.050 1849.810 319.110 ;
        RECT 1891.125 319.095 1891.455 319.110 ;
        RECT 1931.605 319.410 1931.935 319.425 ;
        RECT 1931.605 319.110 1945.490 319.410 ;
        RECT 1931.605 319.095 1931.935 319.110 ;
        RECT 1848.590 317.750 1849.810 318.050 ;
        RECT 1945.190 318.050 1945.490 319.110 ;
        RECT 1993.030 318.730 1993.330 319.790 ;
        RECT 2027.030 319.780 2027.410 319.790 ;
        RECT 2352.750 319.110 2400.890 319.410 ;
        RECT 2089.385 318.730 2089.715 318.745 ;
        RECT 1946.110 318.430 1993.330 318.730 ;
        RECT 2042.710 318.430 2089.715 318.730 ;
        RECT 1946.110 318.050 1946.410 318.430 ;
        RECT 1945.190 317.750 1946.410 318.050 ;
        RECT 2027.950 318.050 2028.330 318.060 ;
        RECT 2042.710 318.050 2043.010 318.430 ;
        RECT 2089.385 318.415 2089.715 318.430 ;
        RECT 2090.765 318.730 2091.095 318.745 ;
        RECT 2185.985 318.730 2186.315 318.745 ;
        RECT 2090.765 318.430 2124.890 318.730 ;
        RECT 2090.765 318.415 2091.095 318.430 ;
        RECT 2027.950 317.750 2043.010 318.050 ;
        RECT 2124.590 318.050 2124.890 318.430 ;
        RECT 2139.310 318.430 2186.315 318.730 ;
        RECT 2139.310 318.050 2139.610 318.430 ;
        RECT 2185.985 318.415 2186.315 318.430 ;
        RECT 2187.365 318.730 2187.695 318.745 ;
        RECT 2282.585 318.730 2282.915 318.745 ;
        RECT 2187.365 318.430 2221.490 318.730 ;
        RECT 2187.365 318.415 2187.695 318.430 ;
        RECT 2124.590 317.750 2139.610 318.050 ;
        RECT 2221.190 318.050 2221.490 318.430 ;
        RECT 2235.910 318.430 2282.915 318.730 ;
        RECT 2235.910 318.050 2236.210 318.430 ;
        RECT 2282.585 318.415 2282.915 318.430 ;
        RECT 2284.425 318.730 2284.755 318.745 ;
        RECT 2284.425 318.430 2331.890 318.730 ;
        RECT 2284.425 318.415 2284.755 318.430 ;
        RECT 2221.190 317.750 2236.210 318.050 ;
        RECT 2331.590 318.050 2331.890 318.430 ;
        RECT 2352.750 318.050 2353.050 319.110 ;
        RECT 2331.590 317.750 2353.050 318.050 ;
        RECT 2400.590 318.050 2400.890 319.110 ;
        RECT 2401.510 319.110 2449.650 319.410 ;
        RECT 2401.510 318.050 2401.810 319.110 ;
        RECT 2449.350 318.730 2449.650 319.110 ;
        RECT 2498.110 319.110 2546.250 319.410 ;
        RECT 2449.350 318.430 2497.490 318.730 ;
        RECT 2400.590 317.750 2401.810 318.050 ;
        RECT 2497.190 318.050 2497.490 318.430 ;
        RECT 2498.110 318.050 2498.410 319.110 ;
        RECT 2545.950 318.730 2546.250 319.110 ;
        RECT 2594.710 319.110 2642.850 319.410 ;
        RECT 2545.950 318.430 2594.090 318.730 ;
        RECT 2497.190 317.750 2498.410 318.050 ;
        RECT 2593.790 318.050 2594.090 318.430 ;
        RECT 2594.710 318.050 2595.010 319.110 ;
        RECT 2642.550 318.730 2642.850 319.110 ;
        RECT 2691.310 319.110 2739.450 319.410 ;
        RECT 2642.550 318.430 2690.690 318.730 ;
        RECT 2593.790 317.750 2595.010 318.050 ;
        RECT 2690.390 318.050 2690.690 318.430 ;
        RECT 2691.310 318.050 2691.610 319.110 ;
        RECT 2739.150 318.730 2739.450 319.110 ;
        RECT 2787.910 319.110 2836.050 319.410 ;
        RECT 2739.150 318.430 2787.290 318.730 ;
        RECT 2690.390 317.750 2691.610 318.050 ;
        RECT 2786.990 318.050 2787.290 318.430 ;
        RECT 2787.910 318.050 2788.210 319.110 ;
        RECT 2835.750 318.730 2836.050 319.110 ;
        RECT 2916.710 318.730 2917.010 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
        RECT 2835.750 318.430 2883.890 318.730 ;
        RECT 2786.990 317.750 2788.210 318.050 ;
        RECT 2883.590 318.050 2883.890 318.430 ;
        RECT 2884.510 318.430 2917.010 318.730 ;
        RECT 2884.510 318.050 2884.810 318.430 ;
        RECT 2883.590 317.750 2884.810 318.050 ;
        RECT 1586.350 317.740 1586.730 317.750 ;
        RECT 1635.110 317.740 1635.490 317.750 ;
        RECT 2027.950 317.740 2028.330 317.750 ;
      LAYER via3 ;
        RECT 1186.180 2896.300 1186.500 2896.620 ;
        RECT 1186.180 318.420 1186.500 318.740 ;
        RECT 1400.540 319.100 1400.860 319.420 ;
        RECT 1442.860 318.420 1443.180 318.740 ;
        RECT 1586.380 319.780 1586.700 320.100 ;
        RECT 1635.140 319.100 1635.460 319.420 ;
        RECT 1400.540 317.740 1400.860 318.060 ;
        RECT 1441.940 317.740 1442.260 318.060 ;
        RECT 1586.380 317.740 1586.700 318.060 ;
        RECT 1635.140 317.740 1635.460 318.060 ;
        RECT 2027.060 319.780 2027.380 320.100 ;
        RECT 2027.980 317.740 2028.300 318.060 ;
      LAYER met4 ;
        RECT 1186.175 2896.295 1186.505 2896.625 ;
        RECT 1186.190 318.745 1186.490 2896.295 ;
        RECT 1586.375 319.775 1586.705 320.105 ;
        RECT 2027.055 319.775 2027.385 320.105 ;
        RECT 1400.535 319.095 1400.865 319.425 ;
        RECT 1186.175 318.415 1186.505 318.745 ;
        RECT 1400.550 318.065 1400.850 319.095 ;
        RECT 1442.855 318.415 1443.185 318.745 ;
        RECT 1400.535 317.735 1400.865 318.065 ;
        RECT 1441.935 318.050 1442.265 318.065 ;
        RECT 1442.870 318.050 1443.170 318.415 ;
        RECT 1586.390 318.065 1586.690 319.775 ;
        RECT 1635.135 319.095 1635.465 319.425 ;
        RECT 1635.150 318.065 1635.450 319.095 ;
        RECT 1441.935 317.750 1443.170 318.050 ;
        RECT 1441.935 317.735 1442.265 317.750 ;
        RECT 1586.375 317.735 1586.705 318.065 ;
        RECT 1635.135 317.735 1635.465 318.065 ;
        RECT 2027.070 318.050 2027.370 319.775 ;
        RECT 2027.975 318.050 2028.305 318.065 ;
        RECT 2027.070 317.750 2028.305 318.050 ;
        RECT 2027.975 317.735 2028.305 317.750 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3500.200 1176.150 3500.260 ;
        RECT 1780.270 3500.200 1780.590 3500.260 ;
        RECT 1175.830 3500.060 1780.590 3500.200 ;
        RECT 1175.830 3500.000 1176.150 3500.060 ;
        RECT 1780.270 3500.000 1780.590 3500.060 ;
      LAYER via ;
        RECT 1175.860 3500.000 1176.120 3500.260 ;
        RECT 1780.300 3500.000 1780.560 3500.260 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3500.290 1176.060 3517.600 ;
        RECT 1175.860 3499.970 1176.120 3500.290 ;
        RECT 1780.300 3499.970 1780.560 3500.290 ;
        RECT 1780.360 2899.250 1780.500 3499.970 ;
        RECT 1785.745 2899.250 1786.025 2900.000 ;
        RECT 1780.360 2899.110 1786.025 2899.250 ;
        RECT 1785.745 2896.000 1786.025 2899.110 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 851.530 3504.620 851.850 3504.680 ;
        RECT 1814.770 3504.620 1815.090 3504.680 ;
        RECT 851.530 3504.480 1815.090 3504.620 ;
        RECT 851.530 3504.420 851.850 3504.480 ;
        RECT 1814.770 3504.420 1815.090 3504.480 ;
      LAYER via ;
        RECT 851.560 3504.420 851.820 3504.680 ;
        RECT 1814.800 3504.420 1815.060 3504.680 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3504.710 851.760 3517.600 ;
        RECT 851.560 3504.390 851.820 3504.710 ;
        RECT 1814.800 3504.390 1815.060 3504.710 ;
        RECT 1814.860 2899.930 1815.000 3504.390 ;
        RECT 1817.025 2899.930 1817.305 2900.000 ;
        RECT 1814.860 2899.790 1817.305 2899.930 ;
        RECT 1817.025 2896.000 1817.305 2899.790 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 527.230 3502.920 527.550 3502.980 ;
        RECT 1842.370 3502.920 1842.690 3502.980 ;
        RECT 527.230 3502.780 1842.690 3502.920 ;
        RECT 527.230 3502.720 527.550 3502.780 ;
        RECT 1842.370 3502.720 1842.690 3502.780 ;
      LAYER via ;
        RECT 527.260 3502.720 527.520 3502.980 ;
        RECT 1842.400 3502.720 1842.660 3502.980 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3503.010 527.460 3517.600 ;
        RECT 527.260 3502.690 527.520 3503.010 ;
        RECT 1842.400 3502.690 1842.660 3503.010 ;
        RECT 1842.460 2900.610 1842.600 3502.690 ;
        RECT 1842.460 2900.470 1846.740 2900.610 ;
        RECT 1846.600 2899.250 1846.740 2900.470 ;
        RECT 1848.765 2899.250 1849.045 2900.000 ;
        RECT 1846.600 2899.110 1849.045 2899.250 ;
        RECT 1848.765 2896.000 1849.045 2899.110 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 1876.870 3501.900 1877.190 3501.960 ;
        RECT 202.470 3501.760 1877.190 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 1876.870 3501.700 1877.190 3501.760 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 1876.900 3501.700 1877.160 3501.960 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 1876.900 3501.670 1877.160 3501.990 ;
        RECT 1876.960 2899.250 1877.100 3501.670 ;
        RECT 1880.505 2899.250 1880.785 2900.000 ;
        RECT 1876.960 2899.110 1880.785 2899.250 ;
        RECT 1880.505 2896.000 1880.785 2899.110 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.550 3408.740 17.870 3408.800 ;
        RECT 1911.370 3408.740 1911.690 3408.800 ;
        RECT 17.550 3408.600 1911.690 3408.740 ;
        RECT 17.550 3408.540 17.870 3408.600 ;
        RECT 1911.370 3408.540 1911.690 3408.600 ;
      LAYER via ;
        RECT 17.580 3408.540 17.840 3408.800 ;
        RECT 1911.400 3408.540 1911.660 3408.800 ;
      LAYER met2 ;
        RECT 17.570 3411.035 17.850 3411.405 ;
        RECT 17.640 3408.830 17.780 3411.035 ;
        RECT 17.580 3408.510 17.840 3408.830 ;
        RECT 1911.400 3408.510 1911.660 3408.830 ;
        RECT 1911.460 2899.930 1911.600 3408.510 ;
        RECT 1911.785 2899.930 1912.065 2900.000 ;
        RECT 1911.460 2899.790 1912.065 2899.930 ;
        RECT 1911.785 2896.000 1912.065 2899.790 ;
      LAYER via2 ;
        RECT 17.570 3411.080 17.850 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.545 3411.370 17.875 3411.385 ;
        RECT -4.800 3411.070 17.875 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.545 3411.055 17.875 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 17.090 3119.060 17.410 3119.120 ;
        RECT 1938.970 3119.060 1939.290 3119.120 ;
        RECT 17.090 3118.920 1939.290 3119.060 ;
        RECT 17.090 3118.860 17.410 3118.920 ;
        RECT 1938.970 3118.860 1939.290 3118.920 ;
      LAYER via ;
        RECT 17.120 3118.860 17.380 3119.120 ;
        RECT 1939.000 3118.860 1939.260 3119.120 ;
      LAYER met2 ;
        RECT 17.110 3124.075 17.390 3124.445 ;
        RECT 17.180 3119.150 17.320 3124.075 ;
        RECT 17.120 3118.830 17.380 3119.150 ;
        RECT 1939.000 3118.830 1939.260 3119.150 ;
        RECT 1939.060 2899.250 1939.200 3118.830 ;
        RECT 1943.525 2899.250 1943.805 2900.000 ;
        RECT 1939.060 2899.110 1943.805 2899.250 ;
        RECT 1943.525 2896.000 1943.805 2899.110 ;
      LAYER via2 ;
        RECT 17.110 3124.120 17.390 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 17.085 3124.410 17.415 3124.425 ;
        RECT -4.800 3124.110 17.415 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 17.085 3124.095 17.415 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 33.650 2900.780 33.970 2900.840 ;
        RECT 1975.310 2900.780 1975.630 2900.840 ;
        RECT 33.650 2900.640 1975.630 2900.780 ;
        RECT 33.650 2900.580 33.970 2900.640 ;
        RECT 1975.310 2900.580 1975.630 2900.640 ;
        RECT 15.710 2841.620 16.030 2841.680 ;
        RECT 33.650 2841.620 33.970 2841.680 ;
        RECT 15.710 2841.480 33.970 2841.620 ;
        RECT 15.710 2841.420 16.030 2841.480 ;
        RECT 33.650 2841.420 33.970 2841.480 ;
      LAYER via ;
        RECT 33.680 2900.580 33.940 2900.840 ;
        RECT 1975.340 2900.580 1975.600 2900.840 ;
        RECT 15.740 2841.420 16.000 2841.680 ;
        RECT 33.680 2841.420 33.940 2841.680 ;
      LAYER met2 ;
        RECT 33.680 2900.550 33.940 2900.870 ;
        RECT 1975.340 2900.550 1975.600 2900.870 ;
        RECT 33.740 2841.710 33.880 2900.550 ;
        RECT 1975.400 2900.000 1975.540 2900.550 ;
        RECT 1975.265 2896.000 1975.545 2900.000 ;
        RECT 15.740 2841.390 16.000 2841.710 ;
        RECT 33.680 2841.390 33.940 2841.710 ;
        RECT 15.800 2836.805 15.940 2841.390 ;
        RECT 15.730 2836.435 16.010 2836.805 ;
      LAYER via2 ;
        RECT 15.730 2836.480 16.010 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 15.705 2836.770 16.035 2836.785 ;
        RECT -4.800 2836.470 16.035 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 15.705 2836.455 16.035 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 32.270 2900.440 32.590 2900.500 ;
        RECT 2006.590 2900.440 2006.910 2900.500 ;
        RECT 32.270 2900.300 2006.910 2900.440 ;
        RECT 32.270 2900.240 32.590 2900.300 ;
        RECT 2006.590 2900.240 2006.910 2900.300 ;
        RECT 15.710 2551.260 16.030 2551.320 ;
        RECT 32.270 2551.260 32.590 2551.320 ;
        RECT 15.710 2551.120 32.590 2551.260 ;
        RECT 15.710 2551.060 16.030 2551.120 ;
        RECT 32.270 2551.060 32.590 2551.120 ;
      LAYER via ;
        RECT 32.300 2900.240 32.560 2900.500 ;
        RECT 2006.620 2900.240 2006.880 2900.500 ;
        RECT 15.740 2551.060 16.000 2551.320 ;
        RECT 32.300 2551.060 32.560 2551.320 ;
      LAYER met2 ;
        RECT 32.300 2900.210 32.560 2900.530 ;
        RECT 2006.620 2900.210 2006.880 2900.530 ;
        RECT 32.360 2551.350 32.500 2900.210 ;
        RECT 2006.680 2900.000 2006.820 2900.210 ;
        RECT 2006.545 2896.000 2006.825 2900.000 ;
        RECT 15.740 2551.030 16.000 2551.350 ;
        RECT 32.300 2551.030 32.560 2551.350 ;
        RECT 15.800 2549.845 15.940 2551.030 ;
        RECT 15.730 2549.475 16.010 2549.845 ;
      LAYER via2 ;
        RECT 15.730 2549.520 16.010 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 15.705 2549.810 16.035 2549.825 ;
        RECT -4.800 2549.510 16.035 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 15.705 2549.495 16.035 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 2915.400 16.490 2915.460 ;
        RECT 2038.330 2915.400 2038.650 2915.460 ;
        RECT 16.170 2915.260 2038.650 2915.400 ;
        RECT 16.170 2915.200 16.490 2915.260 ;
        RECT 2038.330 2915.200 2038.650 2915.260 ;
      LAYER via ;
        RECT 16.200 2915.200 16.460 2915.460 ;
        RECT 2038.360 2915.200 2038.620 2915.460 ;
      LAYER met2 ;
        RECT 16.200 2915.170 16.460 2915.490 ;
        RECT 2038.360 2915.170 2038.620 2915.490 ;
        RECT 16.260 2262.205 16.400 2915.170 ;
        RECT 2038.420 2900.000 2038.560 2915.170 ;
        RECT 2038.285 2896.000 2038.565 2900.000 ;
        RECT 16.190 2261.835 16.470 2262.205 ;
      LAYER via2 ;
        RECT 16.190 2261.880 16.470 2262.160 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 16.165 2262.170 16.495 2262.185 ;
        RECT -4.800 2261.870 16.495 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 16.165 2261.855 16.495 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 31.350 2900.100 31.670 2900.160 ;
        RECT 2070.530 2900.100 2070.850 2900.160 ;
        RECT 31.350 2899.960 2070.850 2900.100 ;
        RECT 31.350 2899.900 31.670 2899.960 ;
        RECT 2070.530 2899.900 2070.850 2899.960 ;
        RECT 16.170 1979.380 16.490 1979.440 ;
        RECT 31.350 1979.380 31.670 1979.440 ;
        RECT 16.170 1979.240 31.670 1979.380 ;
        RECT 16.170 1979.180 16.490 1979.240 ;
        RECT 31.350 1979.180 31.670 1979.240 ;
      LAYER via ;
        RECT 31.380 2899.900 31.640 2900.160 ;
        RECT 2070.560 2899.900 2070.820 2900.160 ;
        RECT 16.200 1979.180 16.460 1979.440 ;
        RECT 31.380 1979.180 31.640 1979.440 ;
      LAYER met2 ;
        RECT 31.380 2899.870 31.640 2900.190 ;
        RECT 2070.025 2899.930 2070.305 2900.000 ;
        RECT 2070.560 2899.930 2070.820 2900.190 ;
        RECT 2070.025 2899.870 2070.820 2899.930 ;
        RECT 31.440 1979.470 31.580 2899.870 ;
        RECT 2070.025 2899.790 2070.760 2899.870 ;
        RECT 2070.025 2896.000 2070.305 2899.790 ;
        RECT 16.200 1979.150 16.460 1979.470 ;
        RECT 31.380 1979.150 31.640 1979.470 ;
        RECT 16.260 1975.245 16.400 1979.150 ;
        RECT 16.190 1974.875 16.470 1975.245 ;
      LAYER via2 ;
        RECT 16.190 1974.920 16.470 1975.200 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 16.165 1975.210 16.495 1975.225 ;
        RECT -4.800 1974.910 16.495 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 16.165 1974.895 16.495 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1531.410 554.100 1531.730 554.160 ;
        RECT 1579.710 554.100 1580.030 554.160 ;
        RECT 1531.410 553.960 1580.030 554.100 ;
        RECT 1531.410 553.900 1531.730 553.960 ;
        RECT 1579.710 553.900 1580.030 553.960 ;
        RECT 1242.070 553.760 1242.390 553.820 ;
        RECT 1270.590 553.760 1270.910 553.820 ;
        RECT 1242.070 553.620 1270.910 553.760 ;
        RECT 1242.070 553.560 1242.390 553.620 ;
        RECT 1270.590 553.560 1270.910 553.620 ;
        RECT 2282.590 553.760 2282.910 553.820 ;
        RECT 2287.190 553.760 2287.510 553.820 ;
        RECT 2282.590 553.620 2287.510 553.760 ;
        RECT 2282.590 553.560 2282.910 553.620 ;
        RECT 2287.190 553.560 2287.510 553.620 ;
        RECT 1296.810 553.080 1297.130 553.140 ;
        RECT 1338.210 553.080 1338.530 553.140 ;
        RECT 1296.810 552.940 1338.530 553.080 ;
        RECT 1296.810 552.880 1297.130 552.940 ;
        RECT 1338.210 552.880 1338.530 552.940 ;
        RECT 2089.390 553.080 2089.710 553.140 ;
        RECT 2090.770 553.080 2091.090 553.140 ;
        RECT 2089.390 552.940 2091.090 553.080 ;
        RECT 2089.390 552.880 2089.710 552.940 ;
        RECT 2090.770 552.880 2091.090 552.940 ;
        RECT 2185.990 553.080 2186.310 553.140 ;
        RECT 2187.370 553.080 2187.690 553.140 ;
        RECT 2185.990 552.940 2187.690 553.080 ;
        RECT 2185.990 552.880 2186.310 552.940 ;
        RECT 2187.370 552.880 2187.690 552.940 ;
      LAYER via ;
        RECT 1531.440 553.900 1531.700 554.160 ;
        RECT 1579.740 553.900 1580.000 554.160 ;
        RECT 1242.100 553.560 1242.360 553.820 ;
        RECT 1270.620 553.560 1270.880 553.820 ;
        RECT 2282.620 553.560 2282.880 553.820 ;
        RECT 2287.220 553.560 2287.480 553.820 ;
        RECT 1296.840 552.880 1297.100 553.140 ;
        RECT 1338.240 552.880 1338.500 553.140 ;
        RECT 2089.420 552.880 2089.680 553.140 ;
        RECT 2090.800 552.880 2091.060 553.140 ;
        RECT 2186.020 552.880 2186.280 553.140 ;
        RECT 2187.400 552.880 2187.660 553.140 ;
      LAYER met2 ;
        RECT 1217.185 2896.530 1217.465 2900.000 ;
        RECT 1218.170 2896.530 1218.450 2896.645 ;
        RECT 1217.185 2896.390 1218.450 2896.530 ;
        RECT 1217.185 2896.000 1217.465 2896.390 ;
        RECT 1218.170 2896.275 1218.450 2896.390 ;
        RECT 1628.030 555.035 1628.310 555.405 ;
        RECT 1531.440 554.045 1531.700 554.190 ;
        RECT 1579.740 554.045 1580.000 554.190 ;
        RECT 1628.100 554.045 1628.240 555.035 ;
        RECT 2439.010 554.355 2439.290 554.725 ;
        RECT 1242.090 553.675 1242.370 554.045 ;
        RECT 1242.100 553.530 1242.360 553.675 ;
        RECT 1270.620 553.530 1270.880 553.850 ;
        RECT 1531.430 553.675 1531.710 554.045 ;
        RECT 1579.730 553.675 1580.010 554.045 ;
        RECT 1628.030 553.675 1628.310 554.045 ;
        RECT 1675.870 553.675 1676.150 554.045 ;
        RECT 2282.610 553.675 2282.890 554.045 ;
        RECT 1270.680 553.365 1270.820 553.530 ;
        RECT 1675.940 553.365 1676.080 553.675 ;
        RECT 2282.620 553.530 2282.880 553.675 ;
        RECT 2287.220 553.530 2287.480 553.850 ;
        RECT 2359.430 553.675 2359.710 554.045 ;
        RECT 2380.130 553.675 2380.410 554.045 ;
        RECT 2287.280 553.365 2287.420 553.530 ;
        RECT 1270.610 552.995 1270.890 553.365 ;
        RECT 1296.830 552.995 1297.110 553.365 ;
        RECT 1296.840 552.850 1297.100 552.995 ;
        RECT 1338.240 552.850 1338.500 553.170 ;
        RECT 1675.870 552.995 1676.150 553.365 ;
        RECT 2089.410 552.995 2089.690 553.365 ;
        RECT 2090.790 552.995 2091.070 553.365 ;
        RECT 2186.010 552.995 2186.290 553.365 ;
        RECT 2187.390 552.995 2187.670 553.365 ;
        RECT 2287.210 552.995 2287.490 553.365 ;
        RECT 2089.420 552.850 2089.680 552.995 ;
        RECT 2090.800 552.850 2091.060 552.995 ;
        RECT 2186.020 552.850 2186.280 552.995 ;
        RECT 2187.400 552.850 2187.660 552.995 ;
        RECT 1338.300 552.685 1338.440 552.850 ;
        RECT 1338.230 552.315 1338.510 552.685 ;
        RECT 2359.500 552.005 2359.640 553.675 ;
        RECT 2380.200 553.250 2380.340 553.675 ;
        RECT 2381.050 553.250 2381.330 553.365 ;
        RECT 2380.200 553.110 2381.330 553.250 ;
        RECT 2381.050 552.995 2381.330 553.110 ;
        RECT 2439.080 552.685 2439.220 554.355 ;
        RECT 2439.010 552.315 2439.290 552.685 ;
        RECT 2359.430 551.635 2359.710 552.005 ;
      LAYER via2 ;
        RECT 1218.170 2896.320 1218.450 2896.600 ;
        RECT 1628.030 555.080 1628.310 555.360 ;
        RECT 2439.010 554.400 2439.290 554.680 ;
        RECT 1242.090 553.720 1242.370 554.000 ;
        RECT 1531.430 553.720 1531.710 554.000 ;
        RECT 1579.730 553.720 1580.010 554.000 ;
        RECT 1628.030 553.720 1628.310 554.000 ;
        RECT 1675.870 553.720 1676.150 554.000 ;
        RECT 2282.610 553.720 2282.890 554.000 ;
        RECT 2359.430 553.720 2359.710 554.000 ;
        RECT 2380.130 553.720 2380.410 554.000 ;
        RECT 1270.610 553.040 1270.890 553.320 ;
        RECT 1296.830 553.040 1297.110 553.320 ;
        RECT 1675.870 553.040 1676.150 553.320 ;
        RECT 2089.410 553.040 2089.690 553.320 ;
        RECT 2090.790 553.040 2091.070 553.320 ;
        RECT 2186.010 553.040 2186.290 553.320 ;
        RECT 2187.390 553.040 2187.670 553.320 ;
        RECT 2287.210 553.040 2287.490 553.320 ;
        RECT 1338.230 552.360 1338.510 552.640 ;
        RECT 2381.050 553.040 2381.330 553.320 ;
        RECT 2439.010 552.360 2439.290 552.640 ;
        RECT 2359.430 551.680 2359.710 551.960 ;
      LAYER met3 ;
        RECT 1218.145 2896.610 1218.475 2896.625 ;
        RECT 1220.190 2896.610 1220.570 2896.620 ;
        RECT 1218.145 2896.310 1220.570 2896.610 ;
        RECT 1218.145 2896.295 1218.475 2896.310 ;
        RECT 1220.190 2896.300 1220.570 2896.310 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2916.710 557.110 2924.800 557.410 ;
        RECT 1483.310 555.370 1483.690 555.380 ;
        RECT 1524.710 555.370 1525.090 555.380 ;
        RECT 1483.310 555.070 1525.090 555.370 ;
        RECT 1483.310 555.060 1483.690 555.070 ;
        RECT 1524.710 555.060 1525.090 555.070 ;
        RECT 1579.910 555.370 1580.290 555.380 ;
        RECT 1628.005 555.370 1628.335 555.385 ;
        RECT 1579.910 555.070 1628.335 555.370 ;
        RECT 1579.910 555.060 1580.290 555.070 ;
        RECT 1628.005 555.055 1628.335 555.070 ;
        RECT 1628.670 554.380 1629.050 554.700 ;
        RECT 2027.030 554.690 2027.410 554.700 ;
        RECT 2438.985 554.690 2439.315 554.705 ;
        RECT 1683.910 554.390 1709.050 554.690 ;
        RECT 1220.190 554.010 1220.570 554.020 ;
        RECT 1242.065 554.010 1242.395 554.025 ;
        RECT 1220.190 553.710 1242.395 554.010 ;
        RECT 1220.190 553.700 1220.570 553.710 ;
        RECT 1242.065 553.695 1242.395 553.710 ;
        RECT 1483.310 553.700 1483.690 554.020 ;
        RECT 1524.710 554.010 1525.090 554.020 ;
        RECT 1531.405 554.010 1531.735 554.025 ;
        RECT 1524.710 553.710 1531.735 554.010 ;
        RECT 1524.710 553.700 1525.090 553.710 ;
        RECT 1270.585 553.330 1270.915 553.345 ;
        RECT 1296.805 553.330 1297.135 553.345 ;
        RECT 1270.585 553.030 1297.135 553.330 ;
        RECT 1270.585 553.015 1270.915 553.030 ;
        RECT 1296.805 553.015 1297.135 553.030 ;
        RECT 1428.110 553.330 1428.490 553.340 ;
        RECT 1483.350 553.330 1483.650 553.700 ;
        RECT 1531.405 553.695 1531.735 553.710 ;
        RECT 1579.705 554.020 1580.035 554.025 ;
        RECT 1579.705 554.010 1580.290 554.020 ;
        RECT 1628.005 554.010 1628.335 554.025 ;
        RECT 1628.710 554.010 1629.010 554.380 ;
        RECT 1579.705 553.710 1580.670 554.010 ;
        RECT 1628.005 553.710 1629.010 554.010 ;
        RECT 1675.845 554.010 1676.175 554.025 ;
        RECT 1683.910 554.010 1684.210 554.390 ;
        RECT 1675.845 553.710 1684.210 554.010 ;
        RECT 1579.705 553.700 1580.290 553.710 ;
        RECT 1579.705 553.695 1580.035 553.700 ;
        RECT 1628.005 553.695 1628.335 553.710 ;
        RECT 1675.845 553.695 1676.175 553.710 ;
        RECT 1428.110 553.030 1483.650 553.330 ;
        RECT 1628.670 553.330 1629.050 553.340 ;
        RECT 1675.845 553.330 1676.175 553.345 ;
        RECT 1628.670 553.030 1676.175 553.330 ;
        RECT 1428.110 553.020 1428.490 553.030 ;
        RECT 1628.670 553.020 1629.050 553.030 ;
        RECT 1675.845 553.015 1676.175 553.030 ;
        RECT 1338.205 552.650 1338.535 552.665 ;
        RECT 1386.710 552.650 1387.090 552.660 ;
        RECT 1338.205 552.350 1387.090 552.650 ;
        RECT 1708.750 552.650 1709.050 554.390 ;
        RECT 1993.030 554.390 2027.410 554.690 ;
        RECT 1848.590 553.710 1897.650 554.010 ;
        RECT 1786.910 553.330 1787.290 553.340 ;
        RECT 1752.910 553.030 1787.290 553.330 ;
        RECT 1752.910 552.650 1753.210 553.030 ;
        RECT 1786.910 553.020 1787.290 553.030 ;
        RECT 1708.750 552.350 1753.210 552.650 ;
        RECT 1787.830 552.650 1788.210 552.660 ;
        RECT 1848.590 552.650 1848.890 553.710 ;
        RECT 1787.830 552.350 1848.890 552.650 ;
        RECT 1897.350 552.650 1897.650 553.710 ;
        RECT 1993.030 553.330 1993.330 554.390 ;
        RECT 2027.030 554.380 2027.410 554.390 ;
        RECT 2415.310 554.390 2439.315 554.690 ;
        RECT 2282.585 554.010 2282.915 554.025 ;
        RECT 2235.910 553.710 2282.915 554.010 ;
        RECT 2089.385 553.330 2089.715 553.345 ;
        RECT 1946.110 553.030 1993.330 553.330 ;
        RECT 2042.710 553.030 2089.715 553.330 ;
        RECT 1946.110 552.650 1946.410 553.030 ;
        RECT 1897.350 552.350 1946.410 552.650 ;
        RECT 2027.950 552.650 2028.330 552.660 ;
        RECT 2042.710 552.650 2043.010 553.030 ;
        RECT 2089.385 553.015 2089.715 553.030 ;
        RECT 2090.765 553.330 2091.095 553.345 ;
        RECT 2185.985 553.330 2186.315 553.345 ;
        RECT 2090.765 553.030 2124.890 553.330 ;
        RECT 2090.765 553.015 2091.095 553.030 ;
        RECT 2027.950 552.350 2043.010 552.650 ;
        RECT 2124.590 552.650 2124.890 553.030 ;
        RECT 2139.310 553.030 2186.315 553.330 ;
        RECT 2139.310 552.650 2139.610 553.030 ;
        RECT 2185.985 553.015 2186.315 553.030 ;
        RECT 2187.365 553.330 2187.695 553.345 ;
        RECT 2187.365 553.030 2221.490 553.330 ;
        RECT 2187.365 553.015 2187.695 553.030 ;
        RECT 2124.590 552.350 2139.610 552.650 ;
        RECT 2221.190 552.650 2221.490 553.030 ;
        RECT 2235.910 552.650 2236.210 553.710 ;
        RECT 2282.585 553.695 2282.915 553.710 ;
        RECT 2359.405 554.010 2359.735 554.025 ;
        RECT 2380.105 554.010 2380.435 554.025 ;
        RECT 2359.405 553.710 2380.435 554.010 ;
        RECT 2359.405 553.695 2359.735 553.710 ;
        RECT 2380.105 553.695 2380.435 553.710 ;
        RECT 2287.185 553.330 2287.515 553.345 ;
        RECT 2311.310 553.330 2311.690 553.340 ;
        RECT 2287.185 553.030 2311.690 553.330 ;
        RECT 2287.185 553.015 2287.515 553.030 ;
        RECT 2311.310 553.020 2311.690 553.030 ;
        RECT 2381.025 553.330 2381.355 553.345 ;
        RECT 2415.310 553.330 2415.610 554.390 ;
        RECT 2438.985 554.375 2439.315 554.390 ;
        RECT 2463.110 554.010 2463.490 554.020 ;
        RECT 2463.110 553.710 2546.250 554.010 ;
        RECT 2463.110 553.700 2463.490 553.710 ;
        RECT 2381.025 553.030 2415.610 553.330 ;
        RECT 2545.950 553.330 2546.250 553.710 ;
        RECT 2594.710 553.710 2642.850 554.010 ;
        RECT 2545.950 553.030 2594.090 553.330 ;
        RECT 2381.025 553.015 2381.355 553.030 ;
        RECT 2221.190 552.350 2236.210 552.650 ;
        RECT 2438.985 552.650 2439.315 552.665 ;
        RECT 2463.110 552.650 2463.490 552.660 ;
        RECT 2438.985 552.350 2463.490 552.650 ;
        RECT 2593.790 552.650 2594.090 553.030 ;
        RECT 2594.710 552.650 2595.010 553.710 ;
        RECT 2642.550 553.330 2642.850 553.710 ;
        RECT 2691.310 553.710 2739.450 554.010 ;
        RECT 2642.550 553.030 2690.690 553.330 ;
        RECT 2593.790 552.350 2595.010 552.650 ;
        RECT 2690.390 552.650 2690.690 553.030 ;
        RECT 2691.310 552.650 2691.610 553.710 ;
        RECT 2739.150 553.330 2739.450 553.710 ;
        RECT 2787.910 553.710 2836.050 554.010 ;
        RECT 2739.150 553.030 2787.290 553.330 ;
        RECT 2690.390 552.350 2691.610 552.650 ;
        RECT 2786.990 552.650 2787.290 553.030 ;
        RECT 2787.910 552.650 2788.210 553.710 ;
        RECT 2835.750 553.330 2836.050 553.710 ;
        RECT 2916.710 553.330 2917.010 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
        RECT 2835.750 553.030 2883.890 553.330 ;
        RECT 2786.990 552.350 2788.210 552.650 ;
        RECT 2883.590 552.650 2883.890 553.030 ;
        RECT 2884.510 553.030 2917.010 553.330 ;
        RECT 2884.510 552.650 2884.810 553.030 ;
        RECT 2883.590 552.350 2884.810 552.650 ;
        RECT 1338.205 552.335 1338.535 552.350 ;
        RECT 1386.710 552.340 1387.090 552.350 ;
        RECT 1787.830 552.340 1788.210 552.350 ;
        RECT 2027.950 552.340 2028.330 552.350 ;
        RECT 2438.985 552.335 2439.315 552.350 ;
        RECT 2463.110 552.340 2463.490 552.350 ;
        RECT 2311.310 551.970 2311.690 551.980 ;
        RECT 2359.405 551.970 2359.735 551.985 ;
        RECT 2311.310 551.670 2359.735 551.970 ;
        RECT 2311.310 551.660 2311.690 551.670 ;
        RECT 2359.405 551.655 2359.735 551.670 ;
        RECT 1386.710 551.290 1387.090 551.300 ;
        RECT 1428.110 551.290 1428.490 551.300 ;
        RECT 1386.710 550.990 1428.490 551.290 ;
        RECT 1386.710 550.980 1387.090 550.990 ;
        RECT 1428.110 550.980 1428.490 550.990 ;
      LAYER via3 ;
        RECT 1220.220 2896.300 1220.540 2896.620 ;
        RECT 1483.340 555.060 1483.660 555.380 ;
        RECT 1524.740 555.060 1525.060 555.380 ;
        RECT 1579.940 555.060 1580.260 555.380 ;
        RECT 1628.700 554.380 1629.020 554.700 ;
        RECT 1220.220 553.700 1220.540 554.020 ;
        RECT 1483.340 553.700 1483.660 554.020 ;
        RECT 1524.740 553.700 1525.060 554.020 ;
        RECT 1428.140 553.020 1428.460 553.340 ;
        RECT 1579.940 553.700 1580.260 554.020 ;
        RECT 1628.700 553.020 1629.020 553.340 ;
        RECT 1386.740 552.340 1387.060 552.660 ;
        RECT 1786.940 553.020 1787.260 553.340 ;
        RECT 1787.860 552.340 1788.180 552.660 ;
        RECT 2027.060 554.380 2027.380 554.700 ;
        RECT 2027.980 552.340 2028.300 552.660 ;
        RECT 2311.340 553.020 2311.660 553.340 ;
        RECT 2463.140 553.700 2463.460 554.020 ;
        RECT 2463.140 552.340 2463.460 552.660 ;
        RECT 2311.340 551.660 2311.660 551.980 ;
        RECT 1386.740 550.980 1387.060 551.300 ;
        RECT 1428.140 550.980 1428.460 551.300 ;
      LAYER met4 ;
        RECT 1220.215 2896.295 1220.545 2896.625 ;
        RECT 1220.230 554.025 1220.530 2896.295 ;
        RECT 1483.335 555.055 1483.665 555.385 ;
        RECT 1524.735 555.055 1525.065 555.385 ;
        RECT 1579.935 555.055 1580.265 555.385 ;
        RECT 1483.350 554.025 1483.650 555.055 ;
        RECT 1524.750 554.025 1525.050 555.055 ;
        RECT 1579.950 554.025 1580.250 555.055 ;
        RECT 1628.695 554.375 1629.025 554.705 ;
        RECT 2027.055 554.375 2027.385 554.705 ;
        RECT 1220.215 553.695 1220.545 554.025 ;
        RECT 1483.335 553.695 1483.665 554.025 ;
        RECT 1524.735 553.695 1525.065 554.025 ;
        RECT 1579.935 553.695 1580.265 554.025 ;
        RECT 1628.710 553.345 1629.010 554.375 ;
        RECT 1428.135 553.015 1428.465 553.345 ;
        RECT 1628.695 553.015 1629.025 553.345 ;
        RECT 1786.935 553.015 1787.265 553.345 ;
        RECT 1386.735 552.335 1387.065 552.665 ;
        RECT 1386.750 551.305 1387.050 552.335 ;
        RECT 1428.150 551.305 1428.450 553.015 ;
        RECT 1786.950 552.650 1787.250 553.015 ;
        RECT 1787.855 552.650 1788.185 552.665 ;
        RECT 1786.950 552.350 1788.185 552.650 ;
        RECT 2027.070 552.650 2027.370 554.375 ;
        RECT 2463.135 553.695 2463.465 554.025 ;
        RECT 2311.335 553.015 2311.665 553.345 ;
        RECT 2027.975 552.650 2028.305 552.665 ;
        RECT 2027.070 552.350 2028.305 552.650 ;
        RECT 1787.855 552.335 1788.185 552.350 ;
        RECT 2027.975 552.335 2028.305 552.350 ;
        RECT 2311.350 551.985 2311.650 553.015 ;
        RECT 2463.150 552.665 2463.450 553.695 ;
        RECT 2463.135 552.335 2463.465 552.665 ;
        RECT 2311.335 551.655 2311.665 551.985 ;
        RECT 1386.735 550.975 1387.065 551.305 ;
        RECT 1428.135 550.975 1428.465 551.305 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2101.370 2914.635 2101.650 2915.005 ;
        RECT 2101.440 2900.000 2101.580 2914.635 ;
        RECT 2101.305 2896.000 2101.585 2900.000 ;
      LAYER via2 ;
        RECT 2101.370 2914.680 2101.650 2914.960 ;
      LAYER met3 ;
        RECT 1239.510 2914.970 1239.890 2914.980 ;
        RECT 2101.345 2914.970 2101.675 2914.985 ;
        RECT 1239.510 2914.670 2101.675 2914.970 ;
        RECT 1239.510 2914.660 1239.890 2914.670 ;
        RECT 2101.345 2914.655 2101.675 2914.670 ;
        RECT 1239.510 1690.290 1239.890 1690.300 ;
        RECT 3.070 1689.990 1239.890 1690.290 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 3.070 1687.570 3.370 1689.990 ;
        RECT 1239.510 1689.980 1239.890 1689.990 ;
        RECT -4.800 1687.270 3.370 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
      LAYER via3 ;
        RECT 1239.540 2914.660 1239.860 2914.980 ;
        RECT 1239.540 1689.980 1239.860 1690.300 ;
      LAYER met4 ;
        RECT 1239.535 2914.655 1239.865 2914.985 ;
        RECT 1239.550 1690.305 1239.850 2914.655 ;
        RECT 1239.535 1689.975 1239.865 1690.305 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.850 2899.760 20.170 2899.820 ;
        RECT 2132.170 2899.760 2132.490 2899.820 ;
        RECT 19.850 2899.620 2132.490 2899.760 ;
        RECT 19.850 2899.560 20.170 2899.620 ;
        RECT 2132.170 2899.560 2132.490 2899.620 ;
      LAYER via ;
        RECT 19.880 2899.560 20.140 2899.820 ;
        RECT 2132.200 2899.560 2132.460 2899.820 ;
      LAYER met2 ;
        RECT 2133.045 2899.930 2133.325 2900.000 ;
        RECT 2132.260 2899.850 2133.325 2899.930 ;
        RECT 19.880 2899.530 20.140 2899.850 ;
        RECT 2132.200 2899.790 2133.325 2899.850 ;
        RECT 2132.200 2899.530 2132.460 2899.790 ;
        RECT 19.940 1472.045 20.080 2899.530 ;
        RECT 2133.045 2896.000 2133.325 2899.790 ;
        RECT 19.870 1471.675 20.150 1472.045 ;
      LAYER via2 ;
        RECT 19.870 1471.720 20.150 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 19.845 1472.010 20.175 1472.025 ;
        RECT -4.800 1471.710 20.175 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 19.845 1471.695 20.175 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2164.850 2913.955 2165.130 2914.325 ;
        RECT 2164.920 2900.000 2165.060 2913.955 ;
        RECT 2164.785 2896.000 2165.065 2900.000 ;
        RECT 15.730 1262.235 16.010 1262.605 ;
        RECT 15.800 1256.485 15.940 1262.235 ;
        RECT 15.730 1256.115 16.010 1256.485 ;
      LAYER via2 ;
        RECT 2164.850 2914.000 2165.130 2914.280 ;
        RECT 15.730 1262.280 16.010 1262.560 ;
        RECT 15.730 1256.160 16.010 1256.440 ;
      LAYER met3 ;
        RECT 1238.590 2914.290 1238.970 2914.300 ;
        RECT 2164.825 2914.290 2165.155 2914.305 ;
        RECT 1238.590 2913.990 2165.155 2914.290 ;
        RECT 1238.590 2913.980 1238.970 2913.990 ;
        RECT 2164.825 2913.975 2165.155 2913.990 ;
        RECT 15.705 1262.570 16.035 1262.585 ;
        RECT 1238.590 1262.570 1238.970 1262.580 ;
        RECT 15.705 1262.270 1238.970 1262.570 ;
        RECT 15.705 1262.255 16.035 1262.270 ;
        RECT 1238.590 1262.260 1238.970 1262.270 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 15.705 1256.450 16.035 1256.465 ;
        RECT -4.800 1256.150 16.035 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 15.705 1256.135 16.035 1256.150 ;
      LAYER via3 ;
        RECT 1238.620 2913.980 1238.940 2914.300 ;
        RECT 1238.620 1262.260 1238.940 1262.580 ;
      LAYER met4 ;
        RECT 1238.615 2913.975 1238.945 2914.305 ;
        RECT 1238.630 1262.585 1238.930 2913.975 ;
        RECT 1238.615 1262.255 1238.945 1262.585 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 18.930 2899.420 19.250 2899.480 ;
        RECT 2194.270 2899.420 2194.590 2899.480 ;
        RECT 18.930 2899.280 2194.590 2899.420 ;
        RECT 18.930 2899.220 19.250 2899.280 ;
        RECT 2194.270 2899.220 2194.590 2899.280 ;
      LAYER via ;
        RECT 18.960 2899.220 19.220 2899.480 ;
        RECT 2194.300 2899.220 2194.560 2899.480 ;
      LAYER met2 ;
        RECT 18.960 2899.190 19.220 2899.510 ;
        RECT 2194.300 2899.250 2194.560 2899.510 ;
        RECT 2196.065 2899.250 2196.345 2900.000 ;
        RECT 2194.300 2899.190 2196.345 2899.250 ;
        RECT 19.020 1040.925 19.160 2899.190 ;
        RECT 2194.360 2899.110 2196.345 2899.190 ;
        RECT 2196.065 2896.000 2196.345 2899.110 ;
        RECT 18.950 1040.555 19.230 1040.925 ;
      LAYER via2 ;
        RECT 18.950 1040.600 19.230 1040.880 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 18.925 1040.890 19.255 1040.905 ;
        RECT -4.800 1040.590 19.255 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 18.925 1040.575 19.255 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2227.870 2913.275 2228.150 2913.645 ;
        RECT 2227.940 2900.000 2228.080 2913.275 ;
        RECT 2227.805 2896.000 2228.085 2900.000 ;
      LAYER via2 ;
        RECT 2227.870 2913.320 2228.150 2913.600 ;
      LAYER met3 ;
        RECT 1237.670 2913.610 1238.050 2913.620 ;
        RECT 2227.845 2913.610 2228.175 2913.625 ;
        RECT 1237.670 2913.310 2228.175 2913.610 ;
        RECT 1237.670 2913.300 1238.050 2913.310 ;
        RECT 2227.845 2913.295 2228.175 2913.310 ;
        RECT 1237.670 828.050 1238.050 828.060 ;
        RECT 3.070 827.750 1238.050 828.050 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 3.070 825.330 3.370 827.750 ;
        RECT 1237.670 827.740 1238.050 827.750 ;
        RECT -4.800 825.030 3.370 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
      LAYER via3 ;
        RECT 1237.700 2913.300 1238.020 2913.620 ;
        RECT 1237.700 827.740 1238.020 828.060 ;
      LAYER met4 ;
        RECT 1237.695 2913.295 1238.025 2913.625 ;
        RECT 1237.710 828.065 1238.010 2913.295 ;
        RECT 1237.695 827.735 1238.025 828.065 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.910 2899.080 25.230 2899.140 ;
        RECT 2257.750 2899.080 2258.070 2899.140 ;
        RECT 24.910 2898.940 2258.070 2899.080 ;
        RECT 24.910 2898.880 25.230 2898.940 ;
        RECT 2257.750 2898.880 2258.070 2898.940 ;
        RECT 13.870 611.560 14.190 611.620 ;
        RECT 24.910 611.560 25.230 611.620 ;
        RECT 13.870 611.420 25.230 611.560 ;
        RECT 13.870 611.360 14.190 611.420 ;
        RECT 24.910 611.360 25.230 611.420 ;
      LAYER via ;
        RECT 24.940 2898.880 25.200 2899.140 ;
        RECT 2257.780 2898.880 2258.040 2899.140 ;
        RECT 13.900 611.360 14.160 611.620 ;
        RECT 24.940 611.360 25.200 611.620 ;
      LAYER met2 ;
        RECT 2259.545 2899.250 2259.825 2900.000 ;
        RECT 2257.840 2899.170 2259.825 2899.250 ;
        RECT 24.940 2898.850 25.200 2899.170 ;
        RECT 2257.780 2899.110 2259.825 2899.170 ;
        RECT 2257.780 2898.850 2258.040 2899.110 ;
        RECT 25.000 611.650 25.140 2898.850 ;
        RECT 2259.545 2896.000 2259.825 2899.110 ;
        RECT 13.900 611.330 14.160 611.650 ;
        RECT 24.940 611.330 25.200 611.650 ;
        RECT 13.960 610.485 14.100 611.330 ;
        RECT 13.890 610.115 14.170 610.485 ;
      LAYER via2 ;
        RECT 13.890 610.160 14.170 610.440 ;
      LAYER met3 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 13.865 610.450 14.195 610.465 ;
        RECT -4.800 610.150 14.195 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 13.865 610.135 14.195 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 24.450 2898.740 24.770 2898.800 ;
        RECT 2291.330 2898.740 2291.650 2898.800 ;
        RECT 24.450 2898.600 2291.650 2898.740 ;
        RECT 24.450 2898.540 24.770 2898.600 ;
        RECT 2291.330 2898.540 2291.650 2898.600 ;
        RECT 13.870 399.060 14.190 399.120 ;
        RECT 24.450 399.060 24.770 399.120 ;
        RECT 13.870 398.920 24.770 399.060 ;
        RECT 13.870 398.860 14.190 398.920 ;
        RECT 24.450 398.860 24.770 398.920 ;
      LAYER via ;
        RECT 24.480 2898.540 24.740 2898.800 ;
        RECT 2291.360 2898.540 2291.620 2898.800 ;
        RECT 13.900 398.860 14.160 399.120 ;
        RECT 24.480 398.860 24.740 399.120 ;
      LAYER met2 ;
        RECT 24.480 2898.510 24.740 2898.830 ;
        RECT 2290.825 2898.570 2291.105 2900.000 ;
        RECT 2291.360 2898.570 2291.620 2898.830 ;
        RECT 2290.825 2898.510 2291.620 2898.570 ;
        RECT 24.540 399.150 24.680 2898.510 ;
        RECT 2290.825 2898.430 2291.560 2898.510 ;
        RECT 2290.825 2896.000 2291.105 2898.430 ;
        RECT 13.900 398.830 14.160 399.150 ;
        RECT 24.480 398.830 24.740 399.150 ;
        RECT 13.960 394.925 14.100 398.830 ;
        RECT 13.890 394.555 14.170 394.925 ;
      LAYER via2 ;
        RECT 13.890 394.600 14.170 394.880 ;
      LAYER met3 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 13.865 394.890 14.195 394.905 ;
        RECT -4.800 394.590 14.195 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 13.865 394.575 14.195 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 30.890 2898.400 31.210 2898.460 ;
        RECT 2321.230 2898.400 2321.550 2898.460 ;
        RECT 30.890 2898.260 2321.550 2898.400 ;
        RECT 30.890 2898.200 31.210 2898.260 ;
        RECT 2321.230 2898.200 2321.550 2898.260 ;
        RECT 15.710 179.420 16.030 179.480 ;
        RECT 30.890 179.420 31.210 179.480 ;
        RECT 15.710 179.280 31.210 179.420 ;
        RECT 15.710 179.220 16.030 179.280 ;
        RECT 30.890 179.220 31.210 179.280 ;
      LAYER via ;
        RECT 30.920 2898.200 31.180 2898.460 ;
        RECT 2321.260 2898.200 2321.520 2898.460 ;
        RECT 15.740 179.220 16.000 179.480 ;
        RECT 30.920 179.220 31.180 179.480 ;
      LAYER met2 ;
        RECT 2322.565 2898.570 2322.845 2900.000 ;
        RECT 2321.320 2898.490 2322.845 2898.570 ;
        RECT 30.920 2898.170 31.180 2898.490 ;
        RECT 2321.260 2898.430 2322.845 2898.490 ;
        RECT 2321.260 2898.170 2321.520 2898.430 ;
        RECT 30.980 179.510 31.120 2898.170 ;
        RECT 2322.565 2896.000 2322.845 2898.430 ;
        RECT 15.740 179.365 16.000 179.510 ;
        RECT 15.730 178.995 16.010 179.365 ;
        RECT 30.920 179.190 31.180 179.510 ;
      LAYER via2 ;
        RECT 15.730 179.040 16.010 179.320 ;
      LAYER met3 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 15.705 179.330 16.035 179.345 ;
        RECT -4.800 179.030 16.035 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 15.705 179.015 16.035 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1891.130 788.700 1891.450 788.760 ;
        RECT 1931.610 788.700 1931.930 788.760 ;
        RECT 1891.130 788.560 1931.930 788.700 ;
        RECT 1891.130 788.500 1891.450 788.560 ;
        RECT 1931.610 788.500 1931.930 788.560 ;
        RECT 1531.870 787.680 1532.190 787.740 ;
        RECT 1579.710 787.680 1580.030 787.740 ;
        RECT 1531.870 787.540 1580.030 787.680 ;
        RECT 1531.870 787.480 1532.190 787.540 ;
        RECT 1579.710 787.480 1580.030 787.540 ;
        RECT 1683.670 787.680 1683.990 787.740 ;
        RECT 1731.510 787.680 1731.830 787.740 ;
        RECT 1683.670 787.540 1731.830 787.680 ;
        RECT 1683.670 787.480 1683.990 787.540 ;
        RECT 1731.510 787.480 1731.830 787.540 ;
        RECT 2089.390 787.680 2089.710 787.740 ;
        RECT 2090.770 787.680 2091.090 787.740 ;
        RECT 2089.390 787.540 2091.090 787.680 ;
        RECT 2089.390 787.480 2089.710 787.540 ;
        RECT 2090.770 787.480 2091.090 787.540 ;
        RECT 2185.990 787.680 2186.310 787.740 ;
        RECT 2187.370 787.680 2187.690 787.740 ;
        RECT 2185.990 787.540 2187.690 787.680 ;
        RECT 2185.990 787.480 2186.310 787.540 ;
        RECT 2187.370 787.480 2187.690 787.540 ;
      LAYER via ;
        RECT 1891.160 788.500 1891.420 788.760 ;
        RECT 1931.640 788.500 1931.900 788.760 ;
        RECT 1531.900 787.480 1532.160 787.740 ;
        RECT 1579.740 787.480 1580.000 787.740 ;
        RECT 1683.700 787.480 1683.960 787.740 ;
        RECT 1731.540 787.480 1731.800 787.740 ;
        RECT 2089.420 787.480 2089.680 787.740 ;
        RECT 2090.800 787.480 2091.060 787.740 ;
        RECT 2186.020 787.480 2186.280 787.740 ;
        RECT 2187.400 787.480 2187.660 787.740 ;
      LAYER met2 ;
        RECT 1247.610 2896.530 1247.890 2896.645 ;
        RECT 1248.465 2896.530 1248.745 2900.000 ;
        RECT 1247.610 2896.390 1248.745 2896.530 ;
        RECT 1247.610 2896.275 1247.890 2896.390 ;
        RECT 1248.465 2896.000 1248.745 2896.390 ;
        RECT 1891.160 788.645 1891.420 788.790 ;
        RECT 1931.640 788.645 1931.900 788.790 ;
        RECT 1586.630 788.275 1586.910 788.645 ;
        RECT 1891.150 788.275 1891.430 788.645 ;
        RECT 1931.630 788.275 1931.910 788.645 ;
        RECT 1531.890 787.595 1532.170 787.965 ;
        RECT 1531.900 787.450 1532.160 787.595 ;
        RECT 1579.740 787.450 1580.000 787.770 ;
        RECT 1579.800 787.285 1579.940 787.450 ;
        RECT 1586.700 787.285 1586.840 788.275 ;
        RECT 1683.690 787.595 1683.970 787.965 ;
        RECT 1800.530 787.850 1800.810 787.965 ;
        RECT 1801.450 787.850 1801.730 787.965 ;
        RECT 1683.700 787.450 1683.960 787.595 ;
        RECT 1731.540 787.450 1731.800 787.770 ;
        RECT 1800.530 787.710 1801.730 787.850 ;
        RECT 1800.530 787.595 1800.810 787.710 ;
        RECT 1801.450 787.595 1801.730 787.710 ;
        RECT 2089.410 787.595 2089.690 787.965 ;
        RECT 2090.790 787.595 2091.070 787.965 ;
        RECT 2186.010 787.595 2186.290 787.965 ;
        RECT 2187.390 787.595 2187.670 787.965 ;
        RECT 2089.420 787.450 2089.680 787.595 ;
        RECT 2090.800 787.450 2091.060 787.595 ;
        RECT 2186.020 787.450 2186.280 787.595 ;
        RECT 2187.400 787.450 2187.660 787.595 ;
        RECT 1731.600 787.285 1731.740 787.450 ;
        RECT 1579.730 786.915 1580.010 787.285 ;
        RECT 1586.630 786.915 1586.910 787.285 ;
        RECT 1731.530 786.915 1731.810 787.285 ;
      LAYER via2 ;
        RECT 1247.610 2896.320 1247.890 2896.600 ;
        RECT 1586.630 788.320 1586.910 788.600 ;
        RECT 1891.150 788.320 1891.430 788.600 ;
        RECT 1931.630 788.320 1931.910 788.600 ;
        RECT 1531.890 787.640 1532.170 787.920 ;
        RECT 1683.690 787.640 1683.970 787.920 ;
        RECT 1800.530 787.640 1800.810 787.920 ;
        RECT 1801.450 787.640 1801.730 787.920 ;
        RECT 2089.410 787.640 2089.690 787.920 ;
        RECT 2090.790 787.640 2091.070 787.920 ;
        RECT 2186.010 787.640 2186.290 787.920 ;
        RECT 2187.390 787.640 2187.670 787.920 ;
        RECT 1579.730 786.960 1580.010 787.240 ;
        RECT 1586.630 786.960 1586.910 787.240 ;
        RECT 1731.530 786.960 1731.810 787.240 ;
      LAYER met3 ;
        RECT 1245.030 2896.610 1245.410 2896.620 ;
        RECT 1247.585 2896.610 1247.915 2896.625 ;
        RECT 1245.030 2896.310 1247.915 2896.610 ;
        RECT 1245.030 2896.300 1245.410 2896.310 ;
        RECT 1247.585 2896.295 1247.915 2896.310 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2916.710 791.710 2924.800 792.010 ;
        RECT 2027.030 789.290 2027.410 789.300 ;
        RECT 1993.030 788.990 2027.410 789.290 ;
        RECT 1586.605 788.610 1586.935 788.625 ;
        RECT 1891.125 788.610 1891.455 788.625 ;
        RECT 1586.605 788.310 1652.930 788.610 ;
        RECT 1586.605 788.295 1586.935 788.310 ;
        RECT 1245.030 787.930 1245.410 787.940 ;
        RECT 1531.865 787.930 1532.195 787.945 ;
        RECT 1245.030 787.630 1270.210 787.930 ;
        RECT 1245.030 787.620 1245.410 787.630 ;
        RECT 1269.910 787.250 1270.210 787.630 ;
        RECT 1376.630 787.630 1532.195 787.930 ;
        RECT 1652.630 787.930 1652.930 788.310 ;
        RECT 1849.510 788.310 1891.455 788.610 ;
        RECT 1683.665 787.930 1683.995 787.945 ;
        RECT 1800.505 787.930 1800.835 787.945 ;
        RECT 1652.630 787.630 1683.995 787.930 ;
        RECT 1376.630 787.250 1376.930 787.630 ;
        RECT 1531.865 787.615 1532.195 787.630 ;
        RECT 1683.665 787.615 1683.995 787.630 ;
        RECT 1752.910 787.630 1800.835 787.930 ;
        RECT 1269.910 786.950 1376.930 787.250 ;
        RECT 1579.705 787.250 1580.035 787.265 ;
        RECT 1586.605 787.250 1586.935 787.265 ;
        RECT 1579.705 786.950 1586.935 787.250 ;
        RECT 1579.705 786.935 1580.035 786.950 ;
        RECT 1586.605 786.935 1586.935 786.950 ;
        RECT 1731.505 787.250 1731.835 787.265 ;
        RECT 1752.910 787.250 1753.210 787.630 ;
        RECT 1800.505 787.615 1800.835 787.630 ;
        RECT 1801.425 787.930 1801.755 787.945 ;
        RECT 1801.425 787.630 1848.890 787.930 ;
        RECT 1801.425 787.615 1801.755 787.630 ;
        RECT 1731.505 786.950 1753.210 787.250 ;
        RECT 1848.590 787.250 1848.890 787.630 ;
        RECT 1849.510 787.250 1849.810 788.310 ;
        RECT 1891.125 788.295 1891.455 788.310 ;
        RECT 1931.605 788.610 1931.935 788.625 ;
        RECT 1931.605 788.310 1945.490 788.610 ;
        RECT 1931.605 788.295 1931.935 788.310 ;
        RECT 1848.590 786.950 1849.810 787.250 ;
        RECT 1945.190 787.250 1945.490 788.310 ;
        RECT 1993.030 787.930 1993.330 788.990 ;
        RECT 2027.030 788.980 2027.410 788.990 ;
        RECT 2352.750 788.310 2400.890 788.610 ;
        RECT 2089.385 787.930 2089.715 787.945 ;
        RECT 1946.110 787.630 1993.330 787.930 ;
        RECT 2042.710 787.630 2089.715 787.930 ;
        RECT 1946.110 787.250 1946.410 787.630 ;
        RECT 1945.190 786.950 1946.410 787.250 ;
        RECT 2027.950 787.250 2028.330 787.260 ;
        RECT 2042.710 787.250 2043.010 787.630 ;
        RECT 2089.385 787.615 2089.715 787.630 ;
        RECT 2090.765 787.930 2091.095 787.945 ;
        RECT 2185.985 787.930 2186.315 787.945 ;
        RECT 2090.765 787.630 2124.890 787.930 ;
        RECT 2090.765 787.615 2091.095 787.630 ;
        RECT 2027.950 786.950 2043.010 787.250 ;
        RECT 2124.590 787.250 2124.890 787.630 ;
        RECT 2139.310 787.630 2186.315 787.930 ;
        RECT 2139.310 787.250 2139.610 787.630 ;
        RECT 2185.985 787.615 2186.315 787.630 ;
        RECT 2187.365 787.930 2187.695 787.945 ;
        RECT 2187.365 787.630 2221.490 787.930 ;
        RECT 2187.365 787.615 2187.695 787.630 ;
        RECT 2124.590 786.950 2139.610 787.250 ;
        RECT 2221.190 787.250 2221.490 787.630 ;
        RECT 2235.910 787.630 2318.090 787.930 ;
        RECT 2235.910 787.250 2236.210 787.630 ;
        RECT 2221.190 786.950 2236.210 787.250 ;
        RECT 2317.790 787.250 2318.090 787.630 ;
        RECT 2352.750 787.250 2353.050 788.310 ;
        RECT 2317.790 786.950 2353.050 787.250 ;
        RECT 2400.590 787.250 2400.890 788.310 ;
        RECT 2401.510 788.310 2449.650 788.610 ;
        RECT 2401.510 787.250 2401.810 788.310 ;
        RECT 2449.350 787.930 2449.650 788.310 ;
        RECT 2498.110 788.310 2546.250 788.610 ;
        RECT 2449.350 787.630 2497.490 787.930 ;
        RECT 2400.590 786.950 2401.810 787.250 ;
        RECT 2497.190 787.250 2497.490 787.630 ;
        RECT 2498.110 787.250 2498.410 788.310 ;
        RECT 2545.950 787.930 2546.250 788.310 ;
        RECT 2594.710 788.310 2642.850 788.610 ;
        RECT 2545.950 787.630 2594.090 787.930 ;
        RECT 2497.190 786.950 2498.410 787.250 ;
        RECT 2593.790 787.250 2594.090 787.630 ;
        RECT 2594.710 787.250 2595.010 788.310 ;
        RECT 2642.550 787.930 2642.850 788.310 ;
        RECT 2691.310 788.310 2739.450 788.610 ;
        RECT 2642.550 787.630 2690.690 787.930 ;
        RECT 2593.790 786.950 2595.010 787.250 ;
        RECT 2690.390 787.250 2690.690 787.630 ;
        RECT 2691.310 787.250 2691.610 788.310 ;
        RECT 2739.150 787.930 2739.450 788.310 ;
        RECT 2787.910 788.310 2836.050 788.610 ;
        RECT 2739.150 787.630 2787.290 787.930 ;
        RECT 2690.390 786.950 2691.610 787.250 ;
        RECT 2786.990 787.250 2787.290 787.630 ;
        RECT 2787.910 787.250 2788.210 788.310 ;
        RECT 2835.750 787.930 2836.050 788.310 ;
        RECT 2916.710 787.930 2917.010 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
        RECT 2835.750 787.630 2883.890 787.930 ;
        RECT 2786.990 786.950 2788.210 787.250 ;
        RECT 2883.590 787.250 2883.890 787.630 ;
        RECT 2884.510 787.630 2917.010 787.930 ;
        RECT 2884.510 787.250 2884.810 787.630 ;
        RECT 2883.590 786.950 2884.810 787.250 ;
        RECT 1731.505 786.935 1731.835 786.950 ;
        RECT 2027.950 786.940 2028.330 786.950 ;
      LAYER via3 ;
        RECT 1245.060 2896.300 1245.380 2896.620 ;
        RECT 1245.060 787.620 1245.380 787.940 ;
        RECT 2027.060 788.980 2027.380 789.300 ;
        RECT 2027.980 786.940 2028.300 787.260 ;
      LAYER met4 ;
        RECT 1245.055 2896.295 1245.385 2896.625 ;
        RECT 1245.070 787.945 1245.370 2896.295 ;
        RECT 2027.055 788.975 2027.385 789.305 ;
        RECT 1245.055 787.615 1245.385 787.945 ;
        RECT 2027.070 787.250 2027.370 788.975 ;
        RECT 2027.975 787.250 2028.305 787.265 ;
        RECT 2027.070 786.950 2028.305 787.250 ;
        RECT 2027.975 786.935 2028.305 786.950 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1280.250 2917.440 1280.570 2917.500 ;
        RECT 2902.210 2917.440 2902.530 2917.500 ;
        RECT 1280.250 2917.300 2902.530 2917.440 ;
        RECT 1280.250 2917.240 1280.570 2917.300 ;
        RECT 2902.210 2917.240 2902.530 2917.300 ;
      LAYER via ;
        RECT 1280.280 2917.240 1280.540 2917.500 ;
        RECT 2902.240 2917.240 2902.500 2917.500 ;
      LAYER met2 ;
        RECT 1280.280 2917.210 1280.540 2917.530 ;
        RECT 2902.240 2917.210 2902.500 2917.530 ;
        RECT 1280.340 2900.000 1280.480 2917.210 ;
        RECT 1280.205 2896.000 1280.485 2900.000 ;
        RECT 2902.300 1026.645 2902.440 2917.210 ;
        RECT 2902.230 1026.275 2902.510 1026.645 ;
      LAYER via2 ;
        RECT 2902.230 1026.320 2902.510 1026.600 ;
      LAYER met3 ;
        RECT 2902.205 1026.610 2902.535 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2902.205 1026.310 2924.800 1026.610 ;
        RECT 2902.205 1026.295 2902.535 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.990 2917.780 1312.310 2917.840 ;
        RECT 2903.590 2917.780 2903.910 2917.840 ;
        RECT 1311.990 2917.640 2903.910 2917.780 ;
        RECT 1311.990 2917.580 1312.310 2917.640 ;
        RECT 2903.590 2917.580 2903.910 2917.640 ;
      LAYER via ;
        RECT 1312.020 2917.580 1312.280 2917.840 ;
        RECT 2903.620 2917.580 2903.880 2917.840 ;
      LAYER met2 ;
        RECT 1312.020 2917.550 1312.280 2917.870 ;
        RECT 2903.620 2917.550 2903.880 2917.870 ;
        RECT 1312.080 2900.000 1312.220 2917.550 ;
        RECT 1311.945 2896.000 1312.225 2900.000 ;
        RECT 2903.680 1261.245 2903.820 2917.550 ;
        RECT 2903.610 1260.875 2903.890 1261.245 ;
      LAYER via2 ;
        RECT 2903.610 1260.920 2903.890 1261.200 ;
      LAYER met3 ;
        RECT 2903.585 1261.210 2903.915 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2903.585 1260.910 2924.800 1261.210 ;
        RECT 2903.585 1260.895 2903.915 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1343.270 2901.460 1343.590 2901.520 ;
        RECT 2349.290 2901.460 2349.610 2901.520 ;
        RECT 1343.270 2901.320 2349.610 2901.460 ;
        RECT 1343.270 2901.260 1343.590 2901.320 ;
        RECT 2349.290 2901.260 2349.610 2901.320 ;
        RECT 2349.290 1497.260 2349.610 1497.320 ;
        RECT 2900.830 1497.260 2901.150 1497.320 ;
        RECT 2349.290 1497.120 2901.150 1497.260 ;
        RECT 2349.290 1497.060 2349.610 1497.120 ;
        RECT 2900.830 1497.060 2901.150 1497.120 ;
      LAYER via ;
        RECT 1343.300 2901.260 1343.560 2901.520 ;
        RECT 2349.320 2901.260 2349.580 2901.520 ;
        RECT 2349.320 1497.060 2349.580 1497.320 ;
        RECT 2900.860 1497.060 2901.120 1497.320 ;
      LAYER met2 ;
        RECT 1343.300 2901.230 1343.560 2901.550 ;
        RECT 2349.320 2901.230 2349.580 2901.550 ;
        RECT 1343.360 2900.000 1343.500 2901.230 ;
        RECT 1343.225 2896.000 1343.505 2900.000 ;
        RECT 2349.380 1497.350 2349.520 2901.230 ;
        RECT 2349.320 1497.030 2349.580 1497.350 ;
        RECT 2900.860 1497.030 2901.120 1497.350 ;
        RECT 2900.920 1495.845 2901.060 1497.030 ;
        RECT 2900.850 1495.475 2901.130 1495.845 ;
      LAYER via2 ;
        RECT 2900.850 1495.520 2901.130 1495.800 ;
      LAYER met3 ;
        RECT 2900.825 1495.810 2901.155 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2900.825 1495.510 2924.800 1495.810 ;
        RECT 2900.825 1495.495 2901.155 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1375.010 2905.880 1375.330 2905.940 ;
        RECT 2350.210 2905.880 2350.530 2905.940 ;
        RECT 1375.010 2905.740 2350.530 2905.880 ;
        RECT 1375.010 2905.680 1375.330 2905.740 ;
        RECT 2350.210 2905.680 2350.530 2905.740 ;
        RECT 2350.210 1731.860 2350.530 1731.920 ;
        RECT 2898.990 1731.860 2899.310 1731.920 ;
        RECT 2350.210 1731.720 2899.310 1731.860 ;
        RECT 2350.210 1731.660 2350.530 1731.720 ;
        RECT 2898.990 1731.660 2899.310 1731.720 ;
      LAYER via ;
        RECT 1375.040 2905.680 1375.300 2905.940 ;
        RECT 2350.240 2905.680 2350.500 2905.940 ;
        RECT 2350.240 1731.660 2350.500 1731.920 ;
        RECT 2899.020 1731.660 2899.280 1731.920 ;
      LAYER met2 ;
        RECT 1375.040 2905.650 1375.300 2905.970 ;
        RECT 2350.240 2905.650 2350.500 2905.970 ;
        RECT 1375.100 2900.000 1375.240 2905.650 ;
        RECT 1374.965 2896.000 1375.245 2900.000 ;
        RECT 2350.300 1731.950 2350.440 2905.650 ;
        RECT 2350.240 1731.630 2350.500 1731.950 ;
        RECT 2899.020 1731.630 2899.280 1731.950 ;
        RECT 2899.080 1730.445 2899.220 1731.630 ;
        RECT 2899.010 1730.075 2899.290 1730.445 ;
      LAYER via2 ;
        RECT 2899.010 1730.120 2899.290 1730.400 ;
      LAYER met3 ;
        RECT 2898.985 1730.410 2899.315 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2898.985 1730.110 2924.800 1730.410 ;
        RECT 2898.985 1730.095 2899.315 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1406.750 2906.220 1407.070 2906.280 ;
        RECT 2350.670 2906.220 2350.990 2906.280 ;
        RECT 1406.750 2906.080 2350.990 2906.220 ;
        RECT 1406.750 2906.020 1407.070 2906.080 ;
        RECT 2350.670 2906.020 2350.990 2906.080 ;
        RECT 2350.670 1966.460 2350.990 1966.520 ;
        RECT 2899.450 1966.460 2899.770 1966.520 ;
        RECT 2350.670 1966.320 2899.770 1966.460 ;
        RECT 2350.670 1966.260 2350.990 1966.320 ;
        RECT 2899.450 1966.260 2899.770 1966.320 ;
      LAYER via ;
        RECT 1406.780 2906.020 1407.040 2906.280 ;
        RECT 2350.700 2906.020 2350.960 2906.280 ;
        RECT 2350.700 1966.260 2350.960 1966.520 ;
        RECT 2899.480 1966.260 2899.740 1966.520 ;
      LAYER met2 ;
        RECT 1406.780 2905.990 1407.040 2906.310 ;
        RECT 2350.700 2905.990 2350.960 2906.310 ;
        RECT 1406.840 2900.000 1406.980 2905.990 ;
        RECT 1406.705 2896.000 1406.985 2900.000 ;
        RECT 2350.760 1966.550 2350.900 2905.990 ;
        RECT 2350.700 1966.230 2350.960 1966.550 ;
        RECT 2899.480 1966.230 2899.740 1966.550 ;
        RECT 2899.540 1965.045 2899.680 1966.230 ;
        RECT 2899.470 1964.675 2899.750 1965.045 ;
      LAYER via2 ;
        RECT 2899.470 1964.720 2899.750 1965.000 ;
      LAYER met3 ;
        RECT 2899.445 1965.010 2899.775 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2899.445 1964.710 2924.800 1965.010 ;
        RECT 2899.445 1964.695 2899.775 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1438.030 2906.900 1438.350 2906.960 ;
        RECT 2352.050 2906.900 2352.370 2906.960 ;
        RECT 1438.030 2906.760 2352.370 2906.900 ;
        RECT 1438.030 2906.700 1438.350 2906.760 ;
        RECT 2352.050 2906.700 2352.370 2906.760 ;
        RECT 2352.050 2201.060 2352.370 2201.120 ;
        RECT 2899.450 2201.060 2899.770 2201.120 ;
        RECT 2352.050 2200.920 2899.770 2201.060 ;
        RECT 2352.050 2200.860 2352.370 2200.920 ;
        RECT 2899.450 2200.860 2899.770 2200.920 ;
      LAYER via ;
        RECT 1438.060 2906.700 1438.320 2906.960 ;
        RECT 2352.080 2906.700 2352.340 2906.960 ;
        RECT 2352.080 2200.860 2352.340 2201.120 ;
        RECT 2899.480 2200.860 2899.740 2201.120 ;
      LAYER met2 ;
        RECT 1438.060 2906.670 1438.320 2906.990 ;
        RECT 2352.080 2906.670 2352.340 2906.990 ;
        RECT 1438.120 2900.000 1438.260 2906.670 ;
        RECT 1437.985 2896.000 1438.265 2900.000 ;
        RECT 2352.140 2201.150 2352.280 2906.670 ;
        RECT 2352.080 2200.830 2352.340 2201.150 ;
        RECT 2899.480 2200.830 2899.740 2201.150 ;
        RECT 2899.540 2199.645 2899.680 2200.830 ;
        RECT 2899.470 2199.275 2899.750 2199.645 ;
      LAYER via2 ;
        RECT 2899.470 2199.320 2899.750 2199.600 ;
      LAYER met3 ;
        RECT 2899.445 2199.610 2899.775 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2899.445 2199.310 2924.800 2199.610 ;
        RECT 2899.445 2199.295 2899.775 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2185.990 201.180 2186.310 201.240 ;
        RECT 2187.830 201.180 2188.150 201.240 ;
        RECT 2185.990 201.040 2188.150 201.180 ;
        RECT 2185.990 200.980 2186.310 201.040 ;
        RECT 2187.830 200.980 2188.150 201.040 ;
        RECT 2282.590 201.180 2282.910 201.240 ;
        RECT 2284.430 201.180 2284.750 201.240 ;
        RECT 2282.590 201.040 2284.750 201.180 ;
        RECT 2282.590 200.980 2282.910 201.040 ;
        RECT 2284.430 200.980 2284.750 201.040 ;
        RECT 2089.390 200.840 2089.710 200.900 ;
        RECT 2090.770 200.840 2091.090 200.900 ;
        RECT 2089.390 200.700 2091.090 200.840 ;
        RECT 2089.390 200.640 2089.710 200.700 ;
        RECT 2090.770 200.640 2091.090 200.700 ;
      LAYER via ;
        RECT 2186.020 200.980 2186.280 201.240 ;
        RECT 2187.860 200.980 2188.120 201.240 ;
        RECT 2282.620 200.980 2282.880 201.240 ;
        RECT 2284.460 200.980 2284.720 201.240 ;
        RECT 2089.420 200.640 2089.680 200.900 ;
        RECT 2090.800 200.640 2091.060 200.900 ;
      LAYER met2 ;
        RECT 1164.285 2896.530 1164.565 2900.000 ;
        RECT 1164.810 2896.530 1165.090 2896.645 ;
        RECT 1164.285 2896.390 1165.090 2896.530 ;
        RECT 1164.285 2896.000 1164.565 2896.390 ;
        RECT 1164.810 2896.275 1165.090 2896.390 ;
        RECT 2186.020 201.125 2186.280 201.270 ;
        RECT 2187.860 201.125 2188.120 201.270 ;
        RECT 2282.620 201.125 2282.880 201.270 ;
        RECT 2284.460 201.125 2284.720 201.270 ;
        RECT 1352.030 200.755 1352.310 201.125 ;
        RECT 1800.530 201.010 1800.810 201.125 ;
        RECT 1801.450 201.010 1801.730 201.125 ;
        RECT 1800.530 200.870 1801.730 201.010 ;
        RECT 1800.530 200.755 1800.810 200.870 ;
        RECT 1801.450 200.755 1801.730 200.870 ;
        RECT 2089.410 200.755 2089.690 201.125 ;
        RECT 2090.790 200.755 2091.070 201.125 ;
        RECT 2186.010 200.755 2186.290 201.125 ;
        RECT 2187.850 200.755 2188.130 201.125 ;
        RECT 2282.610 200.755 2282.890 201.125 ;
        RECT 2284.450 200.755 2284.730 201.125 ;
        RECT 1352.100 200.445 1352.240 200.755 ;
        RECT 2089.420 200.610 2089.680 200.755 ;
        RECT 2090.800 200.610 2091.060 200.755 ;
        RECT 1352.030 200.075 1352.310 200.445 ;
      LAYER via2 ;
        RECT 1164.810 2896.320 1165.090 2896.600 ;
        RECT 1352.030 200.800 1352.310 201.080 ;
        RECT 1800.530 200.800 1800.810 201.080 ;
        RECT 1801.450 200.800 1801.730 201.080 ;
        RECT 2089.410 200.800 2089.690 201.080 ;
        RECT 2090.790 200.800 2091.070 201.080 ;
        RECT 2186.010 200.800 2186.290 201.080 ;
        RECT 2187.850 200.800 2188.130 201.080 ;
        RECT 2282.610 200.800 2282.890 201.080 ;
        RECT 2284.450 200.800 2284.730 201.080 ;
        RECT 1352.030 200.120 1352.310 200.400 ;
      LAYER met3 ;
        RECT 1164.785 2896.620 1165.115 2896.625 ;
        RECT 1164.785 2896.610 1165.370 2896.620 ;
        RECT 1164.785 2896.310 1165.570 2896.610 ;
        RECT 1164.785 2896.300 1165.370 2896.310 ;
        RECT 1164.785 2896.295 1165.115 2896.300 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2916.710 204.870 2924.800 205.170 ;
        RECT 1980.150 202.150 2028.290 202.450 ;
        RECT 1352.710 201.470 1377.850 201.770 ;
        RECT 1352.005 201.090 1352.335 201.105 ;
        RECT 1352.710 201.090 1353.010 201.470 ;
        RECT 1173.310 200.790 1270.210 201.090 ;
        RECT 1164.990 200.410 1165.370 200.420 ;
        RECT 1173.310 200.410 1173.610 200.790 ;
        RECT 1164.990 200.110 1173.610 200.410 ;
        RECT 1269.910 200.410 1270.210 200.790 ;
        RECT 1352.005 200.790 1353.010 201.090 ;
        RECT 1377.550 201.090 1377.850 201.470 ;
        RECT 1655.390 201.470 1704.450 201.770 ;
        RECT 1377.550 200.790 1560.010 201.090 ;
        RECT 1352.005 200.775 1352.335 200.790 ;
        RECT 1352.005 200.410 1352.335 200.425 ;
        RECT 1269.910 200.110 1352.335 200.410 ;
        RECT 1559.710 200.410 1560.010 200.790 ;
        RECT 1655.390 200.410 1655.690 201.470 ;
        RECT 1559.710 200.110 1655.690 200.410 ;
        RECT 1704.150 200.410 1704.450 201.470 ;
        RECT 1849.510 201.470 1949.170 201.770 ;
        RECT 1800.505 201.090 1800.835 201.105 ;
        RECT 1752.910 200.790 1800.835 201.090 ;
        RECT 1752.910 200.410 1753.210 200.790 ;
        RECT 1800.505 200.775 1800.835 200.790 ;
        RECT 1801.425 201.090 1801.755 201.105 ;
        RECT 1801.425 200.790 1848.890 201.090 ;
        RECT 1801.425 200.775 1801.755 200.790 ;
        RECT 1704.150 200.110 1753.210 200.410 ;
        RECT 1848.590 200.410 1848.890 200.790 ;
        RECT 1849.510 200.410 1849.810 201.470 ;
        RECT 1948.870 201.090 1949.170 201.470 ;
        RECT 1980.150 201.090 1980.450 202.150 ;
        RECT 2027.990 201.780 2028.290 202.150 ;
        RECT 2027.950 201.460 2028.330 201.780 ;
        RECT 2352.750 201.470 2400.890 201.770 ;
        RECT 2089.385 201.090 2089.715 201.105 ;
        RECT 1948.870 200.790 1980.450 201.090 ;
        RECT 2042.710 200.790 2089.715 201.090 ;
        RECT 1848.590 200.110 1849.810 200.410 ;
        RECT 2027.950 200.410 2028.330 200.420 ;
        RECT 2042.710 200.410 2043.010 200.790 ;
        RECT 2089.385 200.775 2089.715 200.790 ;
        RECT 2090.765 201.090 2091.095 201.105 ;
        RECT 2185.985 201.090 2186.315 201.105 ;
        RECT 2090.765 200.790 2124.890 201.090 ;
        RECT 2090.765 200.775 2091.095 200.790 ;
        RECT 2027.950 200.110 2043.010 200.410 ;
        RECT 2124.590 200.410 2124.890 200.790 ;
        RECT 2139.310 200.790 2186.315 201.090 ;
        RECT 2139.310 200.410 2139.610 200.790 ;
        RECT 2185.985 200.775 2186.315 200.790 ;
        RECT 2187.825 201.090 2188.155 201.105 ;
        RECT 2282.585 201.090 2282.915 201.105 ;
        RECT 2187.825 200.790 2221.490 201.090 ;
        RECT 2187.825 200.775 2188.155 200.790 ;
        RECT 2124.590 200.110 2139.610 200.410 ;
        RECT 2221.190 200.410 2221.490 200.790 ;
        RECT 2235.910 200.790 2282.915 201.090 ;
        RECT 2235.910 200.410 2236.210 200.790 ;
        RECT 2282.585 200.775 2282.915 200.790 ;
        RECT 2284.425 201.090 2284.755 201.105 ;
        RECT 2284.425 200.790 2331.890 201.090 ;
        RECT 2284.425 200.775 2284.755 200.790 ;
        RECT 2221.190 200.110 2236.210 200.410 ;
        RECT 2331.590 200.410 2331.890 200.790 ;
        RECT 2352.750 200.410 2353.050 201.470 ;
        RECT 2331.590 200.110 2353.050 200.410 ;
        RECT 2400.590 200.410 2400.890 201.470 ;
        RECT 2401.510 201.470 2449.650 201.770 ;
        RECT 2401.510 200.410 2401.810 201.470 ;
        RECT 2449.350 201.090 2449.650 201.470 ;
        RECT 2498.110 201.470 2546.250 201.770 ;
        RECT 2449.350 200.790 2497.490 201.090 ;
        RECT 2400.590 200.110 2401.810 200.410 ;
        RECT 2497.190 200.410 2497.490 200.790 ;
        RECT 2498.110 200.410 2498.410 201.470 ;
        RECT 2545.950 201.090 2546.250 201.470 ;
        RECT 2594.710 201.470 2642.850 201.770 ;
        RECT 2545.950 200.790 2594.090 201.090 ;
        RECT 2497.190 200.110 2498.410 200.410 ;
        RECT 2593.790 200.410 2594.090 200.790 ;
        RECT 2594.710 200.410 2595.010 201.470 ;
        RECT 2642.550 201.090 2642.850 201.470 ;
        RECT 2691.310 201.470 2739.450 201.770 ;
        RECT 2642.550 200.790 2690.690 201.090 ;
        RECT 2593.790 200.110 2595.010 200.410 ;
        RECT 2690.390 200.410 2690.690 200.790 ;
        RECT 2691.310 200.410 2691.610 201.470 ;
        RECT 2739.150 201.090 2739.450 201.470 ;
        RECT 2787.910 201.470 2836.050 201.770 ;
        RECT 2739.150 200.790 2787.290 201.090 ;
        RECT 2690.390 200.110 2691.610 200.410 ;
        RECT 2786.990 200.410 2787.290 200.790 ;
        RECT 2787.910 200.410 2788.210 201.470 ;
        RECT 2835.750 201.090 2836.050 201.470 ;
        RECT 2916.710 201.090 2917.010 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
        RECT 2835.750 200.790 2883.890 201.090 ;
        RECT 2786.990 200.110 2788.210 200.410 ;
        RECT 2883.590 200.410 2883.890 200.790 ;
        RECT 2884.510 200.790 2917.010 201.090 ;
        RECT 2884.510 200.410 2884.810 200.790 ;
        RECT 2883.590 200.110 2884.810 200.410 ;
        RECT 1164.990 200.100 1165.370 200.110 ;
        RECT 1352.005 200.095 1352.335 200.110 ;
        RECT 2027.950 200.100 2028.330 200.110 ;
      LAYER via3 ;
        RECT 1165.020 2896.300 1165.340 2896.620 ;
        RECT 1165.020 200.100 1165.340 200.420 ;
        RECT 2027.980 201.460 2028.300 201.780 ;
        RECT 2027.980 200.100 2028.300 200.420 ;
      LAYER met4 ;
        RECT 1165.015 2896.295 1165.345 2896.625 ;
        RECT 1165.030 200.425 1165.330 2896.295 ;
        RECT 2027.975 201.455 2028.305 201.785 ;
        RECT 2027.990 200.425 2028.290 201.455 ;
        RECT 1165.015 200.095 1165.345 200.425 ;
        RECT 2027.975 200.095 2028.305 200.425 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1480.350 2907.580 1480.670 2907.640 ;
        RECT 2348.370 2907.580 2348.690 2907.640 ;
        RECT 1480.350 2907.440 2348.690 2907.580 ;
        RECT 1480.350 2907.380 1480.670 2907.440 ;
        RECT 2348.370 2907.380 2348.690 2907.440 ;
        RECT 2348.370 2552.960 2348.690 2553.020 ;
        RECT 2898.990 2552.960 2899.310 2553.020 ;
        RECT 2348.370 2552.820 2899.310 2552.960 ;
        RECT 2348.370 2552.760 2348.690 2552.820 ;
        RECT 2898.990 2552.760 2899.310 2552.820 ;
      LAYER via ;
        RECT 1480.380 2907.380 1480.640 2907.640 ;
        RECT 2348.400 2907.380 2348.660 2907.640 ;
        RECT 2348.400 2552.760 2348.660 2553.020 ;
        RECT 2899.020 2552.760 2899.280 2553.020 ;
      LAYER met2 ;
        RECT 1480.380 2907.350 1480.640 2907.670 ;
        RECT 2348.400 2907.350 2348.660 2907.670 ;
        RECT 1480.440 2900.000 1480.580 2907.350 ;
        RECT 1480.305 2896.000 1480.585 2900.000 ;
        RECT 2348.460 2553.050 2348.600 2907.350 ;
        RECT 2348.400 2552.730 2348.660 2553.050 ;
        RECT 2899.020 2552.730 2899.280 2553.050 ;
        RECT 2899.080 2551.885 2899.220 2552.730 ;
        RECT 2899.010 2551.515 2899.290 2551.885 ;
      LAYER via2 ;
        RECT 2899.010 2551.560 2899.290 2551.840 ;
      LAYER met3 ;
        RECT 2898.985 2551.850 2899.315 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2898.985 2551.550 2924.800 2551.850 ;
        RECT 2898.985 2551.535 2899.315 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1512.090 2907.920 1512.410 2907.980 ;
        RECT 2347.910 2907.920 2348.230 2907.980 ;
        RECT 1512.090 2907.780 2348.230 2907.920 ;
        RECT 1512.090 2907.720 1512.410 2907.780 ;
        RECT 2347.910 2907.720 2348.230 2907.780 ;
        RECT 2347.910 2787.560 2348.230 2787.620 ;
        RECT 2898.990 2787.560 2899.310 2787.620 ;
        RECT 2347.910 2787.420 2899.310 2787.560 ;
        RECT 2347.910 2787.360 2348.230 2787.420 ;
        RECT 2898.990 2787.360 2899.310 2787.420 ;
      LAYER via ;
        RECT 1512.120 2907.720 1512.380 2907.980 ;
        RECT 2347.940 2907.720 2348.200 2907.980 ;
        RECT 2347.940 2787.360 2348.200 2787.620 ;
        RECT 2899.020 2787.360 2899.280 2787.620 ;
      LAYER met2 ;
        RECT 1512.120 2907.690 1512.380 2908.010 ;
        RECT 2347.940 2907.690 2348.200 2908.010 ;
        RECT 1512.180 2900.000 1512.320 2907.690 ;
        RECT 1512.045 2896.000 1512.325 2900.000 ;
        RECT 2348.000 2787.650 2348.140 2907.690 ;
        RECT 2347.940 2787.330 2348.200 2787.650 ;
        RECT 2899.020 2787.330 2899.280 2787.650 ;
        RECT 2899.080 2786.485 2899.220 2787.330 ;
        RECT 2899.010 2786.115 2899.290 2786.485 ;
      LAYER via2 ;
        RECT 2899.010 2786.160 2899.290 2786.440 ;
      LAYER met3 ;
        RECT 2898.985 2786.450 2899.315 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2898.985 2786.150 2924.800 2786.450 ;
        RECT 2898.985 2786.135 2899.315 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1545.210 3015.700 1545.530 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 1545.210 3015.560 2901.150 3015.700 ;
        RECT 1545.210 3015.500 1545.530 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 1545.240 3015.500 1545.500 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 1545.240 3015.470 1545.500 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 1543.325 2899.930 1543.605 2900.000 ;
        RECT 1545.300 2899.930 1545.440 3015.470 ;
        RECT 1543.325 2899.790 1545.440 2899.930 ;
        RECT 1543.325 2896.000 1543.605 2899.790 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1579.710 3250.300 1580.030 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 1579.710 3250.160 2901.150 3250.300 ;
        RECT 1579.710 3250.100 1580.030 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
      LAYER via ;
        RECT 1579.740 3250.100 1580.000 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 1579.740 3250.070 1580.000 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 1575.065 2899.250 1575.345 2900.000 ;
        RECT 1579.800 2899.250 1579.940 3250.070 ;
        RECT 1575.065 2899.110 1579.940 2899.250 ;
        RECT 1575.065 2896.000 1575.345 2899.110 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1607.310 3484.900 1607.630 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1607.310 3484.760 2901.150 3484.900 ;
        RECT 1607.310 3484.700 1607.630 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
      LAYER via ;
        RECT 1607.340 3484.700 1607.600 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1607.340 3484.670 1607.600 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1606.805 2899.930 1607.085 2900.000 ;
        RECT 1607.400 2899.930 1607.540 3484.670 ;
        RECT 1606.805 2899.790 1607.540 2899.930 ;
        RECT 1606.805 2896.000 1607.085 2899.790 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1641.810 3504.280 1642.130 3504.340 ;
        RECT 2635.870 3504.280 2636.190 3504.340 ;
        RECT 1641.810 3504.140 2636.190 3504.280 ;
        RECT 1641.810 3504.080 1642.130 3504.140 ;
        RECT 2635.870 3504.080 2636.190 3504.140 ;
      LAYER via ;
        RECT 1641.840 3504.080 1642.100 3504.340 ;
        RECT 2635.900 3504.080 2636.160 3504.340 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3504.370 2636.100 3517.600 ;
        RECT 1641.840 3504.050 1642.100 3504.370 ;
        RECT 2635.900 3504.050 2636.160 3504.370 ;
        RECT 1638.085 2899.250 1638.365 2900.000 ;
        RECT 1641.900 2899.250 1642.040 3504.050 ;
        RECT 1638.085 2899.110 1642.040 2899.250 ;
        RECT 1638.085 2896.000 1638.365 2899.110 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1676.310 3500.540 1676.630 3500.600 ;
        RECT 2311.570 3500.540 2311.890 3500.600 ;
        RECT 1676.310 3500.400 2311.890 3500.540 ;
        RECT 1676.310 3500.340 1676.630 3500.400 ;
        RECT 2311.570 3500.340 2311.890 3500.400 ;
      LAYER via ;
        RECT 1676.340 3500.340 1676.600 3500.600 ;
        RECT 2311.600 3500.340 2311.860 3500.600 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3500.630 2311.800 3517.600 ;
        RECT 1676.340 3500.310 1676.600 3500.630 ;
        RECT 2311.600 3500.310 2311.860 3500.630 ;
        RECT 1676.400 2900.610 1676.540 3500.310 ;
        RECT 1672.260 2900.470 1676.540 2900.610 ;
        RECT 1669.825 2899.250 1670.105 2900.000 ;
        RECT 1672.260 2899.250 1672.400 2900.470 ;
        RECT 1669.825 2899.110 1672.400 2899.250 ;
        RECT 1669.825 2896.000 1670.105 2899.110 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1703.910 3498.840 1704.230 3498.900 ;
        RECT 1987.270 3498.840 1987.590 3498.900 ;
        RECT 1703.910 3498.700 1987.590 3498.840 ;
        RECT 1703.910 3498.640 1704.230 3498.700 ;
        RECT 1987.270 3498.640 1987.590 3498.700 ;
      LAYER via ;
        RECT 1703.940 3498.640 1704.200 3498.900 ;
        RECT 1987.300 3498.640 1987.560 3498.900 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3498.930 1987.500 3517.600 ;
        RECT 1703.940 3498.610 1704.200 3498.930 ;
        RECT 1987.300 3498.610 1987.560 3498.930 ;
        RECT 1701.565 2899.930 1701.845 2900.000 ;
        RECT 1704.000 2899.930 1704.140 3498.610 ;
        RECT 1701.565 2899.790 1704.140 2899.930 ;
        RECT 1701.565 2896.000 1701.845 2899.790 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1662.510 3498.500 1662.830 3498.560 ;
        RECT 1731.970 3498.500 1732.290 3498.560 ;
        RECT 1662.510 3498.360 1732.290 3498.500 ;
        RECT 1662.510 3498.300 1662.830 3498.360 ;
        RECT 1731.970 3498.300 1732.290 3498.360 ;
      LAYER via ;
        RECT 1662.540 3498.300 1662.800 3498.560 ;
        RECT 1732.000 3498.300 1732.260 3498.560 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3498.590 1662.740 3517.600 ;
        RECT 1662.540 3498.270 1662.800 3498.590 ;
        RECT 1732.000 3498.270 1732.260 3498.590 ;
        RECT 1732.060 2899.930 1732.200 3498.270 ;
        RECT 1732.845 2899.930 1733.125 2900.000 ;
        RECT 1732.060 2899.790 1733.125 2899.930 ;
        RECT 1732.845 2896.000 1733.125 2899.790 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1338.210 3499.860 1338.530 3499.920 ;
        RECT 1759.570 3499.860 1759.890 3499.920 ;
        RECT 1338.210 3499.720 1759.890 3499.860 ;
        RECT 1338.210 3499.660 1338.530 3499.720 ;
        RECT 1759.570 3499.660 1759.890 3499.720 ;
      LAYER via ;
        RECT 1338.240 3499.660 1338.500 3499.920 ;
        RECT 1759.600 3499.660 1759.860 3499.920 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3499.950 1338.440 3517.600 ;
        RECT 1338.240 3499.630 1338.500 3499.950 ;
        RECT 1759.600 3499.630 1759.860 3499.950 ;
        RECT 1759.660 2899.250 1759.800 3499.630 ;
        RECT 1764.585 2899.250 1764.865 2900.000 ;
        RECT 1759.660 2899.110 1764.865 2899.250 ;
        RECT 1764.585 2896.000 1764.865 2899.110 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2089.390 435.780 2089.710 435.840 ;
        RECT 2093.070 435.780 2093.390 435.840 ;
        RECT 2089.390 435.640 2093.390 435.780 ;
        RECT 2089.390 435.580 2089.710 435.640 ;
        RECT 2093.070 435.580 2093.390 435.640 ;
        RECT 2270.170 435.780 2270.490 435.840 ;
        RECT 2317.090 435.780 2317.410 435.840 ;
        RECT 2270.170 435.640 2317.410 435.780 ;
        RECT 2270.170 435.580 2270.490 435.640 ;
        RECT 2317.090 435.580 2317.410 435.640 ;
        RECT 2318.470 435.780 2318.790 435.840 ;
        RECT 2339.630 435.780 2339.950 435.840 ;
        RECT 2318.470 435.640 2339.950 435.780 ;
        RECT 2318.470 435.580 2318.790 435.640 ;
        RECT 2339.630 435.580 2339.950 435.640 ;
        RECT 2473.030 435.780 2473.350 435.840 ;
        RECT 2511.210 435.780 2511.530 435.840 ;
        RECT 2473.030 435.640 2511.530 435.780 ;
        RECT 2473.030 435.580 2473.350 435.640 ;
        RECT 2511.210 435.580 2511.530 435.640 ;
        RECT 1683.670 435.440 1683.990 435.500 ;
        RECT 1731.510 435.440 1731.830 435.500 ;
        RECT 1683.670 435.300 1731.830 435.440 ;
        RECT 1683.670 435.240 1683.990 435.300 ;
        RECT 1731.510 435.240 1731.830 435.300 ;
        RECT 1895.270 435.440 1895.590 435.500 ;
        RECT 1931.150 435.440 1931.470 435.500 ;
        RECT 1895.270 435.300 1931.470 435.440 ;
        RECT 1895.270 435.240 1895.590 435.300 ;
        RECT 1931.150 435.240 1931.470 435.300 ;
        RECT 1980.370 435.440 1980.690 435.500 ;
        RECT 2027.750 435.440 2028.070 435.500 ;
        RECT 1980.370 435.300 2028.070 435.440 ;
        RECT 1980.370 435.240 1980.690 435.300 ;
        RECT 2027.750 435.240 2028.070 435.300 ;
        RECT 2185.990 435.440 2186.310 435.500 ;
        RECT 2187.370 435.440 2187.690 435.500 ;
        RECT 2185.990 435.300 2187.690 435.440 ;
        RECT 2185.990 435.240 2186.310 435.300 ;
        RECT 2187.370 435.240 2187.690 435.300 ;
      LAYER via ;
        RECT 2089.420 435.580 2089.680 435.840 ;
        RECT 2093.100 435.580 2093.360 435.840 ;
        RECT 2270.200 435.580 2270.460 435.840 ;
        RECT 2317.120 435.580 2317.380 435.840 ;
        RECT 2318.500 435.580 2318.760 435.840 ;
        RECT 2339.660 435.580 2339.920 435.840 ;
        RECT 2473.060 435.580 2473.320 435.840 ;
        RECT 2511.240 435.580 2511.500 435.840 ;
        RECT 1683.700 435.240 1683.960 435.500 ;
        RECT 1731.540 435.240 1731.800 435.500 ;
        RECT 1895.300 435.240 1895.560 435.500 ;
        RECT 1931.180 435.240 1931.440 435.500 ;
        RECT 1980.400 435.240 1980.660 435.500 ;
        RECT 2027.780 435.240 2028.040 435.500 ;
        RECT 2186.020 435.240 2186.280 435.500 ;
        RECT 2187.400 435.240 2187.660 435.500 ;
      LAYER met2 ;
        RECT 1196.025 2896.530 1196.305 2900.000 ;
        RECT 1197.010 2896.530 1197.290 2896.645 ;
        RECT 1196.025 2896.390 1197.290 2896.530 ;
        RECT 1196.025 2896.000 1196.305 2896.390 ;
        RECT 1197.010 2896.275 1197.290 2896.390 ;
        RECT 1659.310 436.715 1659.590 437.085 ;
        RECT 2456.030 436.715 2456.310 437.085 ;
        RECT 1431.150 436.035 1431.430 436.405 ;
        RECT 1365.370 435.610 1365.650 435.725 ;
        RECT 1366.290 435.610 1366.570 435.725 ;
        RECT 1365.370 435.470 1366.570 435.610 ;
        RECT 1365.370 435.355 1365.650 435.470 ;
        RECT 1366.290 435.355 1366.570 435.470 ;
        RECT 1431.220 435.045 1431.360 436.035 ;
        RECT 1659.380 435.725 1659.520 436.715 ;
        RECT 2270.190 436.035 2270.470 436.405 ;
        RECT 2339.650 436.035 2339.930 436.405 ;
        RECT 2380.130 436.035 2380.410 436.405 ;
        RECT 2270.260 435.870 2270.400 436.035 ;
        RECT 2089.420 435.725 2089.680 435.870 ;
        RECT 2093.100 435.725 2093.360 435.870 ;
        RECT 1659.310 435.355 1659.590 435.725 ;
        RECT 1683.690 435.355 1683.970 435.725 ;
        RECT 1683.700 435.210 1683.960 435.355 ;
        RECT 1731.540 435.210 1731.800 435.530 ;
        RECT 1895.290 435.355 1895.570 435.725 ;
        RECT 1895.300 435.210 1895.560 435.355 ;
        RECT 1931.180 435.210 1931.440 435.530 ;
        RECT 1980.390 435.355 1980.670 435.725 ;
        RECT 1980.400 435.210 1980.660 435.355 ;
        RECT 2027.780 435.210 2028.040 435.530 ;
        RECT 2089.410 435.355 2089.690 435.725 ;
        RECT 2093.090 435.355 2093.370 435.725 ;
        RECT 2186.010 435.355 2186.290 435.725 ;
        RECT 2187.390 435.355 2187.670 435.725 ;
        RECT 2270.200 435.550 2270.460 435.870 ;
        RECT 2317.110 435.525 2317.390 435.895 ;
        RECT 2339.720 435.870 2339.860 436.035 ;
        RECT 2318.500 435.725 2318.760 435.870 ;
        RECT 2318.490 435.355 2318.770 435.725 ;
        RECT 2339.660 435.550 2339.920 435.870 ;
        RECT 2380.200 435.610 2380.340 436.035 ;
        RECT 2381.050 435.610 2381.330 435.725 ;
        RECT 2380.200 435.470 2381.330 435.610 ;
        RECT 2381.050 435.355 2381.330 435.470 ;
        RECT 2186.020 435.210 2186.280 435.355 ;
        RECT 2187.400 435.210 2187.660 435.355 ;
        RECT 1731.600 435.045 1731.740 435.210 ;
        RECT 1431.150 434.675 1431.430 435.045 ;
        RECT 1731.530 434.675 1731.810 435.045 ;
        RECT 1931.240 434.930 1931.380 435.210 ;
        RECT 2027.840 435.045 2027.980 435.210 ;
        RECT 2456.100 435.045 2456.240 436.715 ;
        RECT 2511.230 436.035 2511.510 436.405 ;
        RECT 2511.300 435.870 2511.440 436.035 ;
        RECT 2473.060 435.550 2473.320 435.870 ;
        RECT 2511.240 435.550 2511.500 435.870 ;
        RECT 2473.120 435.045 2473.260 435.550 ;
        RECT 1931.630 434.930 1931.910 435.045 ;
        RECT 1931.240 434.790 1931.910 434.930 ;
        RECT 1931.630 434.675 1931.910 434.790 ;
        RECT 2027.770 434.675 2028.050 435.045 ;
        RECT 2456.030 434.675 2456.310 435.045 ;
        RECT 2473.050 434.675 2473.330 435.045 ;
      LAYER via2 ;
        RECT 1197.010 2896.320 1197.290 2896.600 ;
        RECT 1659.310 436.760 1659.590 437.040 ;
        RECT 2456.030 436.760 2456.310 437.040 ;
        RECT 1431.150 436.080 1431.430 436.360 ;
        RECT 1365.370 435.400 1365.650 435.680 ;
        RECT 1366.290 435.400 1366.570 435.680 ;
        RECT 2270.190 436.080 2270.470 436.360 ;
        RECT 2339.650 436.080 2339.930 436.360 ;
        RECT 2380.130 436.080 2380.410 436.360 ;
        RECT 1659.310 435.400 1659.590 435.680 ;
        RECT 1683.690 435.400 1683.970 435.680 ;
        RECT 1895.290 435.400 1895.570 435.680 ;
        RECT 1980.390 435.400 1980.670 435.680 ;
        RECT 2089.410 435.400 2089.690 435.680 ;
        RECT 2093.090 435.400 2093.370 435.680 ;
        RECT 2186.010 435.400 2186.290 435.680 ;
        RECT 2187.390 435.400 2187.670 435.680 ;
        RECT 2317.110 435.570 2317.390 435.850 ;
        RECT 2318.490 435.400 2318.770 435.680 ;
        RECT 2381.050 435.400 2381.330 435.680 ;
        RECT 1431.150 434.720 1431.430 435.000 ;
        RECT 1731.530 434.720 1731.810 435.000 ;
        RECT 2511.230 436.080 2511.510 436.360 ;
        RECT 1931.630 434.720 1931.910 435.000 ;
        RECT 2027.770 434.720 2028.050 435.000 ;
        RECT 2456.030 434.720 2456.310 435.000 ;
        RECT 2473.050 434.720 2473.330 435.000 ;
      LAYER met3 ;
        RECT 1196.985 2896.610 1197.315 2896.625 ;
        RECT 1199.950 2896.610 1200.330 2896.620 ;
        RECT 1196.985 2896.310 1200.330 2896.610 ;
        RECT 1196.985 2896.295 1197.315 2896.310 ;
        RECT 1199.950 2896.300 1200.330 2896.310 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2916.710 439.470 2924.800 439.770 ;
        RECT 1497.110 437.050 1497.490 437.060 ;
        RECT 1659.285 437.050 1659.615 437.065 ;
        RECT 1497.110 436.750 1510.330 437.050 ;
        RECT 1497.110 436.740 1497.490 436.750 ;
        RECT 1199.950 436.370 1200.330 436.380 ;
        RECT 1431.125 436.370 1431.455 436.385 ;
        RECT 1199.950 436.070 1249.050 436.370 ;
        RECT 1199.950 436.060 1200.330 436.070 ;
        RECT 1248.750 435.690 1249.050 436.070 ;
        RECT 1369.270 436.070 1431.455 436.370 ;
        RECT 1365.345 435.690 1365.675 435.705 ;
        RECT 1248.750 435.390 1365.675 435.690 ;
        RECT 1365.345 435.375 1365.675 435.390 ;
        RECT 1366.265 435.690 1366.595 435.705 ;
        RECT 1369.270 435.690 1369.570 436.070 ;
        RECT 1431.125 436.055 1431.455 436.070 ;
        RECT 1497.110 435.690 1497.490 435.700 ;
        RECT 1366.265 435.390 1369.570 435.690 ;
        RECT 1447.470 435.390 1497.490 435.690 ;
        RECT 1510.030 435.690 1510.330 436.750 ;
        RECT 1611.230 436.750 1659.615 437.050 ;
        RECT 1611.230 435.690 1611.530 436.750 ;
        RECT 1659.285 436.735 1659.615 436.750 ;
        RECT 2407.910 437.050 2408.290 437.060 ;
        RECT 2456.005 437.050 2456.335 437.065 ;
        RECT 2407.910 436.750 2456.335 437.050 ;
        RECT 2407.910 436.740 2408.290 436.750 ;
        RECT 2456.005 436.735 2456.335 436.750 ;
        RECT 2270.165 436.370 2270.495 436.385 ;
        RECT 2235.910 436.070 2270.495 436.370 ;
        RECT 1510.030 435.390 1559.090 435.690 ;
        RECT 1366.265 435.375 1366.595 435.390 ;
        RECT 1431.125 435.010 1431.455 435.025 ;
        RECT 1447.470 435.010 1447.770 435.390 ;
        RECT 1497.110 435.380 1497.490 435.390 ;
        RECT 1431.125 434.710 1447.770 435.010 ;
        RECT 1558.790 435.010 1559.090 435.390 ;
        RECT 1559.710 435.390 1611.530 435.690 ;
        RECT 1659.285 435.690 1659.615 435.705 ;
        RECT 1683.665 435.690 1683.995 435.705 ;
        RECT 1895.265 435.690 1895.595 435.705 ;
        RECT 1980.365 435.690 1980.695 435.705 ;
        RECT 2089.385 435.690 2089.715 435.705 ;
        RECT 1659.285 435.390 1683.995 435.690 ;
        RECT 1559.710 435.010 1560.010 435.390 ;
        RECT 1659.285 435.375 1659.615 435.390 ;
        RECT 1683.665 435.375 1683.995 435.390 ;
        RECT 1752.910 435.390 1801.050 435.690 ;
        RECT 1558.790 434.710 1560.010 435.010 ;
        RECT 1731.505 435.010 1731.835 435.025 ;
        RECT 1752.910 435.010 1753.210 435.390 ;
        RECT 1731.505 434.710 1753.210 435.010 ;
        RECT 1800.750 435.010 1801.050 435.390 ;
        RECT 1849.510 435.390 1895.595 435.690 ;
        RECT 1849.510 435.010 1849.810 435.390 ;
        RECT 1895.265 435.375 1895.595 435.390 ;
        RECT 1946.110 435.390 1980.695 435.690 ;
        RECT 1800.750 434.710 1849.810 435.010 ;
        RECT 1931.605 435.010 1931.935 435.025 ;
        RECT 1946.110 435.010 1946.410 435.390 ;
        RECT 1980.365 435.375 1980.695 435.390 ;
        RECT 2042.710 435.390 2089.715 435.690 ;
        RECT 1931.605 434.710 1946.410 435.010 ;
        RECT 2027.745 435.010 2028.075 435.025 ;
        RECT 2042.710 435.010 2043.010 435.390 ;
        RECT 2089.385 435.375 2089.715 435.390 ;
        RECT 2093.065 435.690 2093.395 435.705 ;
        RECT 2185.985 435.690 2186.315 435.705 ;
        RECT 2093.065 435.390 2124.890 435.690 ;
        RECT 2093.065 435.375 2093.395 435.390 ;
        RECT 2027.745 434.710 2043.010 435.010 ;
        RECT 2124.590 435.010 2124.890 435.390 ;
        RECT 2139.310 435.390 2186.315 435.690 ;
        RECT 2139.310 435.010 2139.610 435.390 ;
        RECT 2185.985 435.375 2186.315 435.390 ;
        RECT 2187.365 435.690 2187.695 435.705 ;
        RECT 2187.365 435.390 2221.490 435.690 ;
        RECT 2187.365 435.375 2187.695 435.390 ;
        RECT 2124.590 434.710 2139.610 435.010 ;
        RECT 2221.190 435.010 2221.490 435.390 ;
        RECT 2235.910 435.010 2236.210 436.070 ;
        RECT 2270.165 436.055 2270.495 436.070 ;
        RECT 2339.625 436.370 2339.955 436.385 ;
        RECT 2380.105 436.370 2380.435 436.385 ;
        RECT 2339.625 436.070 2380.435 436.370 ;
        RECT 2339.625 436.055 2339.955 436.070 ;
        RECT 2380.105 436.055 2380.435 436.070 ;
        RECT 2511.205 436.370 2511.535 436.385 ;
        RECT 2511.205 436.070 2546.250 436.370 ;
        RECT 2511.205 436.055 2511.535 436.070 ;
        RECT 2317.085 435.860 2317.415 435.875 ;
        RECT 2317.085 435.690 2318.090 435.860 ;
        RECT 2318.465 435.690 2318.795 435.705 ;
        RECT 2317.085 435.560 2318.795 435.690 ;
        RECT 2317.085 435.545 2317.415 435.560 ;
        RECT 2317.790 435.390 2318.795 435.560 ;
        RECT 2318.465 435.375 2318.795 435.390 ;
        RECT 2381.025 435.690 2381.355 435.705 ;
        RECT 2407.910 435.690 2408.290 435.700 ;
        RECT 2381.025 435.390 2408.290 435.690 ;
        RECT 2545.950 435.690 2546.250 436.070 ;
        RECT 2594.710 436.070 2642.850 436.370 ;
        RECT 2545.950 435.390 2594.090 435.690 ;
        RECT 2381.025 435.375 2381.355 435.390 ;
        RECT 2407.910 435.380 2408.290 435.390 ;
        RECT 2221.190 434.710 2236.210 435.010 ;
        RECT 2456.005 435.010 2456.335 435.025 ;
        RECT 2473.025 435.010 2473.355 435.025 ;
        RECT 2456.005 434.710 2473.355 435.010 ;
        RECT 2593.790 435.010 2594.090 435.390 ;
        RECT 2594.710 435.010 2595.010 436.070 ;
        RECT 2642.550 435.690 2642.850 436.070 ;
        RECT 2691.310 436.070 2739.450 436.370 ;
        RECT 2642.550 435.390 2690.690 435.690 ;
        RECT 2593.790 434.710 2595.010 435.010 ;
        RECT 2690.390 435.010 2690.690 435.390 ;
        RECT 2691.310 435.010 2691.610 436.070 ;
        RECT 2739.150 435.690 2739.450 436.070 ;
        RECT 2787.910 436.070 2836.050 436.370 ;
        RECT 2739.150 435.390 2787.290 435.690 ;
        RECT 2690.390 434.710 2691.610 435.010 ;
        RECT 2786.990 435.010 2787.290 435.390 ;
        RECT 2787.910 435.010 2788.210 436.070 ;
        RECT 2835.750 435.690 2836.050 436.070 ;
        RECT 2916.710 435.690 2917.010 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
        RECT 2835.750 435.390 2883.890 435.690 ;
        RECT 2786.990 434.710 2788.210 435.010 ;
        RECT 2883.590 435.010 2883.890 435.390 ;
        RECT 2884.510 435.390 2917.010 435.690 ;
        RECT 2884.510 435.010 2884.810 435.390 ;
        RECT 2883.590 434.710 2884.810 435.010 ;
        RECT 1431.125 434.695 1431.455 434.710 ;
        RECT 1731.505 434.695 1731.835 434.710 ;
        RECT 1931.605 434.695 1931.935 434.710 ;
        RECT 2027.745 434.695 2028.075 434.710 ;
        RECT 2456.005 434.695 2456.335 434.710 ;
        RECT 2473.025 434.695 2473.355 434.710 ;
      LAYER via3 ;
        RECT 1199.980 2896.300 1200.300 2896.620 ;
        RECT 1497.140 436.740 1497.460 437.060 ;
        RECT 1199.980 436.060 1200.300 436.380 ;
        RECT 1497.140 435.380 1497.460 435.700 ;
        RECT 2407.940 436.740 2408.260 437.060 ;
        RECT 2407.940 435.380 2408.260 435.700 ;
      LAYER met4 ;
        RECT 1199.975 2896.295 1200.305 2896.625 ;
        RECT 1199.990 436.385 1200.290 2896.295 ;
        RECT 1497.135 436.735 1497.465 437.065 ;
        RECT 2407.935 436.735 2408.265 437.065 ;
        RECT 1199.975 436.055 1200.305 436.385 ;
        RECT 1497.150 435.705 1497.450 436.735 ;
        RECT 2407.950 435.705 2408.250 436.735 ;
        RECT 1497.135 435.375 1497.465 435.705 ;
        RECT 2407.935 435.375 2408.265 435.705 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3504.960 1014.230 3505.020 ;
        RECT 1794.070 3504.960 1794.390 3505.020 ;
        RECT 1013.910 3504.820 1794.390 3504.960 ;
        RECT 1013.910 3504.760 1014.230 3504.820 ;
        RECT 1794.070 3504.760 1794.390 3504.820 ;
      LAYER via ;
        RECT 1013.940 3504.760 1014.200 3505.020 ;
        RECT 1794.100 3504.760 1794.360 3505.020 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3505.050 1014.140 3517.600 ;
        RECT 1013.940 3504.730 1014.200 3505.050 ;
        RECT 1794.100 3504.730 1794.360 3505.050 ;
        RECT 1794.160 2899.250 1794.300 3504.730 ;
        RECT 1796.325 2899.250 1796.605 2900.000 ;
        RECT 1794.160 2899.110 1796.605 2899.250 ;
        RECT 1796.325 2896.000 1796.605 2899.110 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3503.260 689.470 3503.320 ;
        RECT 1821.670 3503.260 1821.990 3503.320 ;
        RECT 689.150 3503.120 1821.990 3503.260 ;
        RECT 689.150 3503.060 689.470 3503.120 ;
        RECT 1821.670 3503.060 1821.990 3503.120 ;
      LAYER via ;
        RECT 689.180 3503.060 689.440 3503.320 ;
        RECT 1821.700 3503.060 1821.960 3503.320 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3503.350 689.380 3517.600 ;
        RECT 689.180 3503.030 689.440 3503.350 ;
        RECT 1821.700 3503.030 1821.960 3503.350 ;
        RECT 1821.760 2900.610 1821.900 3503.030 ;
        RECT 1821.760 2900.470 1826.040 2900.610 ;
        RECT 1825.900 2899.930 1826.040 2900.470 ;
        RECT 1827.605 2899.930 1827.885 2900.000 ;
        RECT 1825.900 2899.790 1827.885 2899.930 ;
        RECT 1827.605 2896.000 1827.885 2899.790 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3502.240 365.170 3502.300 ;
        RECT 1856.170 3502.240 1856.490 3502.300 ;
        RECT 364.850 3502.100 1856.490 3502.240 ;
        RECT 364.850 3502.040 365.170 3502.100 ;
        RECT 1856.170 3502.040 1856.490 3502.100 ;
      LAYER via ;
        RECT 364.880 3502.040 365.140 3502.300 ;
        RECT 1856.200 3502.040 1856.460 3502.300 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3502.330 365.080 3517.600 ;
        RECT 364.880 3502.010 365.140 3502.330 ;
        RECT 1856.200 3502.010 1856.460 3502.330 ;
        RECT 1856.260 2899.250 1856.400 3502.010 ;
        RECT 1859.345 2899.250 1859.625 2900.000 ;
        RECT 1856.260 2899.110 1859.625 2899.250 ;
        RECT 1859.345 2896.000 1859.625 2899.110 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3501.845 40.780 3517.600 ;
        RECT 40.570 3501.475 40.850 3501.845 ;
        RECT 1890.690 3501.475 1890.970 3501.845 ;
        RECT 1890.760 2899.930 1890.900 3501.475 ;
        RECT 1891.085 2899.930 1891.365 2900.000 ;
        RECT 1890.760 2899.790 1891.365 2899.930 ;
        RECT 1891.085 2896.000 1891.365 2899.790 ;
      LAYER via2 ;
        RECT 40.570 3501.520 40.850 3501.800 ;
        RECT 1890.690 3501.520 1890.970 3501.800 ;
      LAYER met3 ;
        RECT 40.545 3501.810 40.875 3501.825 ;
        RECT 1890.665 3501.810 1890.995 3501.825 ;
        RECT 40.545 3501.510 1890.995 3501.810 ;
        RECT 40.545 3501.495 40.875 3501.510 ;
        RECT 1890.665 3501.495 1890.995 3501.510 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 3263.900 15.570 3263.960 ;
        RECT 1918.270 3263.900 1918.590 3263.960 ;
        RECT 15.250 3263.760 1918.590 3263.900 ;
        RECT 15.250 3263.700 15.570 3263.760 ;
        RECT 1918.270 3263.700 1918.590 3263.760 ;
      LAYER via ;
        RECT 15.280 3263.700 15.540 3263.960 ;
        RECT 1918.300 3263.700 1918.560 3263.960 ;
      LAYER met2 ;
        RECT 15.270 3267.555 15.550 3267.925 ;
        RECT 15.340 3263.990 15.480 3267.555 ;
        RECT 15.280 3263.670 15.540 3263.990 ;
        RECT 1918.300 3263.670 1918.560 3263.990 ;
        RECT 1918.360 2899.250 1918.500 3263.670 ;
        RECT 1922.365 2899.250 1922.645 2900.000 ;
        RECT 1918.360 2899.110 1922.645 2899.250 ;
        RECT 1922.365 2896.000 1922.645 2899.110 ;
      LAYER via2 ;
        RECT 15.270 3267.600 15.550 3267.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 15.245 3267.890 15.575 3267.905 ;
        RECT -4.800 3267.590 15.575 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 15.245 3267.575 15.575 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.170 2974.220 16.490 2974.280 ;
        RECT 1952.770 2974.220 1953.090 2974.280 ;
        RECT 16.170 2974.080 1953.090 2974.220 ;
        RECT 16.170 2974.020 16.490 2974.080 ;
        RECT 1952.770 2974.020 1953.090 2974.080 ;
      LAYER via ;
        RECT 16.200 2974.020 16.460 2974.280 ;
        RECT 1952.800 2974.020 1953.060 2974.280 ;
      LAYER met2 ;
        RECT 16.190 2979.915 16.470 2980.285 ;
        RECT 16.260 2974.310 16.400 2979.915 ;
        RECT 16.200 2973.990 16.460 2974.310 ;
        RECT 1952.800 2973.990 1953.060 2974.310 ;
        RECT 1952.860 2899.930 1953.000 2973.990 ;
        RECT 1954.105 2899.930 1954.385 2900.000 ;
        RECT 1952.860 2899.790 1954.385 2899.930 ;
        RECT 1954.105 2896.000 1954.385 2899.790 ;
      LAYER via2 ;
        RECT 16.190 2979.960 16.470 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 16.165 2980.250 16.495 2980.265 ;
        RECT -4.800 2979.950 16.495 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 16.165 2979.935 16.495 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1983.665 2892.805 1983.835 2896.715 ;
      LAYER mcon ;
        RECT 1983.665 2896.545 1983.835 2896.715 ;
      LAYER met1 ;
        RECT 1983.590 2896.700 1983.910 2896.760 ;
        RECT 1983.395 2896.560 1983.910 2896.700 ;
        RECT 1983.590 2896.500 1983.910 2896.560 ;
        RECT 32.730 2892.960 33.050 2893.020 ;
        RECT 1983.605 2892.960 1983.895 2893.005 ;
        RECT 32.730 2892.820 1983.895 2892.960 ;
        RECT 32.730 2892.760 33.050 2892.820 ;
        RECT 1983.605 2892.775 1983.895 2892.820 ;
        RECT 15.250 2695.420 15.570 2695.480 ;
        RECT 32.730 2695.420 33.050 2695.480 ;
        RECT 15.250 2695.280 33.050 2695.420 ;
        RECT 15.250 2695.220 15.570 2695.280 ;
        RECT 32.730 2695.220 33.050 2695.280 ;
      LAYER via ;
        RECT 1983.620 2896.500 1983.880 2896.760 ;
        RECT 32.760 2892.760 33.020 2893.020 ;
        RECT 15.280 2695.220 15.540 2695.480 ;
        RECT 32.760 2695.220 33.020 2695.480 ;
      LAYER met2 ;
        RECT 1983.620 2896.530 1983.880 2896.790 ;
        RECT 1985.385 2896.530 1985.665 2900.000 ;
        RECT 1983.620 2896.470 1985.665 2896.530 ;
        RECT 1983.680 2896.390 1985.665 2896.470 ;
        RECT 1985.385 2896.000 1985.665 2896.390 ;
        RECT 32.760 2892.730 33.020 2893.050 ;
        RECT 32.820 2695.510 32.960 2892.730 ;
        RECT 15.280 2695.190 15.540 2695.510 ;
        RECT 32.760 2695.190 33.020 2695.510 ;
        RECT 15.340 2693.325 15.480 2695.190 ;
        RECT 15.270 2692.955 15.550 2693.325 ;
      LAYER via2 ;
        RECT 15.270 2693.000 15.550 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 15.245 2693.290 15.575 2693.305 ;
        RECT -4.800 2692.990 15.575 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 15.245 2692.975 15.575 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 31.810 2916.420 32.130 2916.480 ;
        RECT 2017.170 2916.420 2017.490 2916.480 ;
        RECT 31.810 2916.280 2017.490 2916.420 ;
        RECT 31.810 2916.220 32.130 2916.280 ;
        RECT 2017.170 2916.220 2017.490 2916.280 ;
        RECT 15.710 2406.420 16.030 2406.480 ;
        RECT 31.810 2406.420 32.130 2406.480 ;
        RECT 15.710 2406.280 32.130 2406.420 ;
        RECT 15.710 2406.220 16.030 2406.280 ;
        RECT 31.810 2406.220 32.130 2406.280 ;
      LAYER via ;
        RECT 31.840 2916.220 32.100 2916.480 ;
        RECT 2017.200 2916.220 2017.460 2916.480 ;
        RECT 15.740 2406.220 16.000 2406.480 ;
        RECT 31.840 2406.220 32.100 2406.480 ;
      LAYER met2 ;
        RECT 31.840 2916.190 32.100 2916.510 ;
        RECT 2017.200 2916.190 2017.460 2916.510 ;
        RECT 31.900 2406.510 32.040 2916.190 ;
        RECT 2017.260 2900.000 2017.400 2916.190 ;
        RECT 2017.125 2896.000 2017.405 2900.000 ;
        RECT 15.740 2406.190 16.000 2406.510 ;
        RECT 31.840 2406.190 32.100 2406.510 ;
        RECT 15.800 2405.685 15.940 2406.190 ;
        RECT 15.730 2405.315 16.010 2405.685 ;
      LAYER via2 ;
        RECT 15.730 2405.360 16.010 2405.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 15.705 2405.650 16.035 2405.665 ;
        RECT -4.800 2405.350 16.035 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 15.705 2405.335 16.035 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.750 2915.740 27.070 2915.800 ;
        RECT 2048.910 2915.740 2049.230 2915.800 ;
        RECT 26.750 2915.600 2049.230 2915.740 ;
        RECT 26.750 2915.540 27.070 2915.600 ;
        RECT 2048.910 2915.540 2049.230 2915.600 ;
        RECT 13.870 2124.220 14.190 2124.280 ;
        RECT 26.750 2124.220 27.070 2124.280 ;
        RECT 13.870 2124.080 27.070 2124.220 ;
        RECT 13.870 2124.020 14.190 2124.080 ;
        RECT 26.750 2124.020 27.070 2124.080 ;
      LAYER via ;
        RECT 26.780 2915.540 27.040 2915.800 ;
        RECT 2048.940 2915.540 2049.200 2915.800 ;
        RECT 13.900 2124.020 14.160 2124.280 ;
        RECT 26.780 2124.020 27.040 2124.280 ;
      LAYER met2 ;
        RECT 26.780 2915.510 27.040 2915.830 ;
        RECT 2048.940 2915.510 2049.200 2915.830 ;
        RECT 26.840 2124.310 26.980 2915.510 ;
        RECT 2049.000 2900.000 2049.140 2915.510 ;
        RECT 2048.865 2896.000 2049.145 2900.000 ;
        RECT 13.900 2123.990 14.160 2124.310 ;
        RECT 26.780 2123.990 27.040 2124.310 ;
        RECT 13.960 2118.725 14.100 2123.990 ;
        RECT 13.890 2118.355 14.170 2118.725 ;
      LAYER via2 ;
        RECT 13.890 2118.400 14.170 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 13.865 2118.690 14.195 2118.705 ;
        RECT -4.800 2118.390 14.195 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 13.865 2118.375 14.195 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2078.425 2892.465 2078.595 2896.715 ;
      LAYER mcon ;
        RECT 2078.425 2896.545 2078.595 2896.715 ;
      LAYER met1 ;
        RECT 2078.350 2896.700 2078.670 2896.760 ;
        RECT 2078.155 2896.560 2078.670 2896.700 ;
        RECT 2078.350 2896.500 2078.670 2896.560 ;
        RECT 16.630 2892.620 16.950 2892.680 ;
        RECT 2078.365 2892.620 2078.655 2892.665 ;
        RECT 16.630 2892.480 2078.655 2892.620 ;
        RECT 16.630 2892.420 16.950 2892.480 ;
        RECT 2078.365 2892.435 2078.655 2892.480 ;
      LAYER via ;
        RECT 2078.380 2896.500 2078.640 2896.760 ;
        RECT 16.660 2892.420 16.920 2892.680 ;
      LAYER met2 ;
        RECT 2078.380 2896.530 2078.640 2896.790 ;
        RECT 2080.145 2896.530 2080.425 2900.000 ;
        RECT 2078.380 2896.470 2080.425 2896.530 ;
        RECT 2078.440 2896.390 2080.425 2896.470 ;
        RECT 2080.145 2896.000 2080.425 2896.390 ;
        RECT 16.660 2892.390 16.920 2892.710 ;
        RECT 16.720 1831.085 16.860 2892.390 ;
        RECT 16.650 1830.715 16.930 1831.085 ;
      LAYER via2 ;
        RECT 16.650 1830.760 16.930 1831.040 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 16.625 1831.050 16.955 1831.065 ;
        RECT -4.800 1830.750 16.955 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 16.625 1830.735 16.955 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1891.130 671.060 1891.450 671.120 ;
        RECT 1931.610 671.060 1931.930 671.120 ;
        RECT 1891.130 670.920 1931.930 671.060 ;
        RECT 1891.130 670.860 1891.450 670.920 ;
        RECT 1931.610 670.860 1931.930 670.920 ;
        RECT 2282.590 670.720 2282.910 670.780 ;
        RECT 2287.190 670.720 2287.510 670.780 ;
        RECT 2282.590 670.580 2287.510 670.720 ;
        RECT 2282.590 670.520 2282.910 670.580 ;
        RECT 2287.190 670.520 2287.510 670.580 ;
        RECT 1545.210 670.380 1545.530 670.440 ;
        RECT 1579.710 670.380 1580.030 670.440 ;
        RECT 1545.210 670.240 1580.030 670.380 ;
        RECT 1545.210 670.180 1545.530 670.240 ;
        RECT 1579.710 670.180 1580.030 670.240 ;
        RECT 2185.990 670.380 2186.310 670.440 ;
        RECT 2187.830 670.380 2188.150 670.440 ;
        RECT 2185.990 670.240 2188.150 670.380 ;
        RECT 2185.990 670.180 2186.310 670.240 ;
        RECT 2187.830 670.180 2188.150 670.240 ;
        RECT 2377.810 670.380 2378.130 670.440 ;
        RECT 2414.610 670.380 2414.930 670.440 ;
        RECT 2377.810 670.240 2414.930 670.380 ;
        RECT 2377.810 670.180 2378.130 670.240 ;
        RECT 2414.610 670.180 2414.930 670.240 ;
        RECT 2089.390 670.040 2089.710 670.100 ;
        RECT 2090.770 670.040 2091.090 670.100 ;
        RECT 2089.390 669.900 2091.090 670.040 ;
        RECT 2089.390 669.840 2089.710 669.900 ;
        RECT 2090.770 669.840 2091.090 669.900 ;
      LAYER via ;
        RECT 1891.160 670.860 1891.420 671.120 ;
        RECT 1931.640 670.860 1931.900 671.120 ;
        RECT 2282.620 670.520 2282.880 670.780 ;
        RECT 2287.220 670.520 2287.480 670.780 ;
        RECT 1545.240 670.180 1545.500 670.440 ;
        RECT 1579.740 670.180 1580.000 670.440 ;
        RECT 2186.020 670.180 2186.280 670.440 ;
        RECT 2187.860 670.180 2188.120 670.440 ;
        RECT 2377.840 670.180 2378.100 670.440 ;
        RECT 2414.640 670.180 2414.900 670.440 ;
        RECT 2089.420 669.840 2089.680 670.100 ;
        RECT 2090.800 669.840 2091.060 670.100 ;
      LAYER met2 ;
        RECT 1226.910 2896.530 1227.190 2896.645 ;
        RECT 1227.765 2896.530 1228.045 2900.000 ;
        RECT 1226.910 2896.390 1228.045 2896.530 ;
        RECT 1226.910 2896.275 1227.190 2896.390 ;
        RECT 1227.765 2896.000 1228.045 2896.390 ;
        RECT 1338.230 672.675 1338.510 673.045 ;
        RECT 1338.300 671.685 1338.440 672.675 ;
        RECT 1338.230 671.315 1338.510 671.685 ;
        RECT 1351.570 671.570 1351.850 671.685 ;
        RECT 1352.490 671.570 1352.770 671.685 ;
        RECT 1351.570 671.430 1352.770 671.570 ;
        RECT 1351.570 671.315 1351.850 671.430 ;
        RECT 1352.490 671.315 1352.770 671.430 ;
        RECT 2439.010 671.315 2439.290 671.685 ;
        RECT 1891.160 671.005 1891.420 671.150 ;
        RECT 1931.640 671.005 1931.900 671.150 ;
        RECT 1434.830 670.635 1435.110 671.005 ;
        RECT 1579.730 670.635 1580.010 671.005 ;
        RECT 1642.290 670.635 1642.570 671.005 ;
        RECT 1891.150 670.635 1891.430 671.005 ;
        RECT 1931.630 670.635 1931.910 671.005 ;
        RECT 2282.610 670.635 2282.890 671.005 ;
        RECT 1434.900 668.965 1435.040 670.635 ;
        RECT 1579.800 670.470 1579.940 670.635 ;
        RECT 1545.240 670.325 1545.500 670.470 ;
        RECT 1459.210 669.955 1459.490 670.325 ;
        RECT 1545.230 669.955 1545.510 670.325 ;
        RECT 1579.740 670.150 1580.000 670.470 ;
        RECT 1459.280 668.965 1459.420 669.955 ;
        RECT 1642.360 669.645 1642.500 670.635 ;
        RECT 2282.620 670.490 2282.880 670.635 ;
        RECT 2287.220 670.490 2287.480 670.810 ;
        RECT 2186.020 670.325 2186.280 670.470 ;
        RECT 2187.860 670.325 2188.120 670.470 ;
        RECT 2287.280 670.325 2287.420 670.490 ;
        RECT 2377.840 670.325 2378.100 670.470 ;
        RECT 2414.640 670.325 2414.900 670.470 ;
        RECT 1800.530 670.210 1800.810 670.325 ;
        RECT 1801.450 670.210 1801.730 670.325 ;
        RECT 1800.530 670.070 1801.730 670.210 ;
        RECT 1800.530 669.955 1800.810 670.070 ;
        RECT 1801.450 669.955 1801.730 670.070 ;
        RECT 2089.410 669.955 2089.690 670.325 ;
        RECT 2090.790 669.955 2091.070 670.325 ;
        RECT 2186.010 669.955 2186.290 670.325 ;
        RECT 2187.850 669.955 2188.130 670.325 ;
        RECT 2287.210 669.955 2287.490 670.325 ;
        RECT 2377.830 669.955 2378.110 670.325 ;
        RECT 2414.630 669.955 2414.910 670.325 ;
        RECT 2089.420 669.810 2089.680 669.955 ;
        RECT 2090.800 669.810 2091.060 669.955 ;
        RECT 2439.080 669.645 2439.220 671.315 ;
        RECT 1642.290 669.275 1642.570 669.645 ;
        RECT 2439.010 669.275 2439.290 669.645 ;
        RECT 1434.830 668.595 1435.110 668.965 ;
        RECT 1459.210 668.595 1459.490 668.965 ;
      LAYER via2 ;
        RECT 1226.910 2896.320 1227.190 2896.600 ;
        RECT 1338.230 672.720 1338.510 673.000 ;
        RECT 1338.230 671.360 1338.510 671.640 ;
        RECT 1351.570 671.360 1351.850 671.640 ;
        RECT 1352.490 671.360 1352.770 671.640 ;
        RECT 2439.010 671.360 2439.290 671.640 ;
        RECT 1434.830 670.680 1435.110 670.960 ;
        RECT 1579.730 670.680 1580.010 670.960 ;
        RECT 1642.290 670.680 1642.570 670.960 ;
        RECT 1891.150 670.680 1891.430 670.960 ;
        RECT 1931.630 670.680 1931.910 670.960 ;
        RECT 2282.610 670.680 2282.890 670.960 ;
        RECT 1459.210 670.000 1459.490 670.280 ;
        RECT 1545.230 670.000 1545.510 670.280 ;
        RECT 1800.530 670.000 1800.810 670.280 ;
        RECT 1801.450 670.000 1801.730 670.280 ;
        RECT 2089.410 670.000 2089.690 670.280 ;
        RECT 2090.790 670.000 2091.070 670.280 ;
        RECT 2186.010 670.000 2186.290 670.280 ;
        RECT 2187.850 670.000 2188.130 670.280 ;
        RECT 2287.210 670.000 2287.490 670.280 ;
        RECT 2377.830 670.000 2378.110 670.280 ;
        RECT 2414.630 670.000 2414.910 670.280 ;
        RECT 1642.290 669.320 1642.570 669.600 ;
        RECT 2439.010 669.320 2439.290 669.600 ;
        RECT 1434.830 668.640 1435.110 668.920 ;
        RECT 1459.210 668.640 1459.490 668.920 ;
      LAYER met3 ;
        RECT 1226.885 2896.620 1227.215 2896.625 ;
        RECT 1226.630 2896.610 1227.215 2896.620 ;
        RECT 1226.430 2896.310 1227.215 2896.610 ;
        RECT 1226.630 2896.300 1227.215 2896.310 ;
        RECT 1226.885 2896.295 1227.215 2896.300 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2916.710 674.070 2924.800 674.370 ;
        RECT 1290.110 673.010 1290.490 673.020 ;
        RECT 1338.205 673.010 1338.535 673.025 ;
        RECT 1290.110 672.710 1338.535 673.010 ;
        RECT 1290.110 672.700 1290.490 672.710 ;
        RECT 1338.205 672.695 1338.535 672.710 ;
        RECT 1338.205 671.650 1338.535 671.665 ;
        RECT 1351.545 671.650 1351.875 671.665 ;
        RECT 1338.205 671.350 1351.875 671.650 ;
        RECT 1338.205 671.335 1338.535 671.350 ;
        RECT 1351.545 671.335 1351.875 671.350 ;
        RECT 1352.465 671.650 1352.795 671.665 ;
        RECT 2438.985 671.650 2439.315 671.665 ;
        RECT 1352.465 671.350 1363.130 671.650 ;
        RECT 1352.465 671.335 1352.795 671.350 ;
        RECT 1226.630 670.970 1227.010 670.980 ;
        RECT 1290.110 670.970 1290.490 670.980 ;
        RECT 1226.630 670.670 1290.490 670.970 ;
        RECT 1362.830 670.970 1363.130 671.350 ;
        RECT 1980.150 671.350 2028.290 671.650 ;
        RECT 1434.805 670.970 1435.135 670.985 ;
        RECT 1362.830 670.670 1435.135 670.970 ;
        RECT 1226.630 670.660 1227.010 670.670 ;
        RECT 1290.110 670.660 1290.490 670.670 ;
        RECT 1434.805 670.655 1435.135 670.670 ;
        RECT 1579.705 670.970 1580.035 670.985 ;
        RECT 1642.265 670.970 1642.595 670.985 ;
        RECT 1891.125 670.970 1891.455 670.985 ;
        RECT 1579.705 670.670 1617.970 670.970 ;
        RECT 1579.705 670.655 1580.035 670.670 ;
        RECT 1459.185 670.290 1459.515 670.305 ;
        RECT 1545.205 670.290 1545.535 670.305 ;
        RECT 1459.185 669.990 1545.535 670.290 ;
        RECT 1459.185 669.975 1459.515 669.990 ;
        RECT 1545.205 669.975 1545.535 669.990 ;
        RECT 1617.670 669.610 1617.970 670.670 ;
        RECT 1642.265 670.670 1704.450 670.970 ;
        RECT 1642.265 670.655 1642.595 670.670 ;
        RECT 1642.265 669.610 1642.595 669.625 ;
        RECT 1617.670 669.310 1642.595 669.610 ;
        RECT 1704.150 669.610 1704.450 670.670 ;
        RECT 1849.510 670.670 1891.455 670.970 ;
        RECT 1800.505 670.290 1800.835 670.305 ;
        RECT 1752.910 669.990 1800.835 670.290 ;
        RECT 1752.910 669.610 1753.210 669.990 ;
        RECT 1800.505 669.975 1800.835 669.990 ;
        RECT 1801.425 670.290 1801.755 670.305 ;
        RECT 1801.425 669.990 1848.890 670.290 ;
        RECT 1801.425 669.975 1801.755 669.990 ;
        RECT 1704.150 669.310 1753.210 669.610 ;
        RECT 1848.590 669.610 1848.890 669.990 ;
        RECT 1849.510 669.610 1849.810 670.670 ;
        RECT 1891.125 670.655 1891.455 670.670 ;
        RECT 1931.605 670.970 1931.935 670.985 ;
        RECT 1931.605 670.670 1945.490 670.970 ;
        RECT 1931.605 670.655 1931.935 670.670 ;
        RECT 1848.590 669.310 1849.810 669.610 ;
        RECT 1945.190 669.610 1945.490 670.670 ;
        RECT 1980.150 670.290 1980.450 671.350 ;
        RECT 2027.990 670.980 2028.290 671.350 ;
        RECT 2415.310 671.350 2439.315 671.650 ;
        RECT 2027.950 670.660 2028.330 670.980 ;
        RECT 2282.585 670.970 2282.915 670.985 ;
        RECT 2235.910 670.670 2282.915 670.970 ;
        RECT 2089.385 670.290 2089.715 670.305 ;
        RECT 1946.110 669.990 1980.450 670.290 ;
        RECT 2042.710 669.990 2089.715 670.290 ;
        RECT 1946.110 669.610 1946.410 669.990 ;
        RECT 1945.190 669.310 1946.410 669.610 ;
        RECT 2027.950 669.610 2028.330 669.620 ;
        RECT 2042.710 669.610 2043.010 669.990 ;
        RECT 2089.385 669.975 2089.715 669.990 ;
        RECT 2090.765 670.290 2091.095 670.305 ;
        RECT 2185.985 670.290 2186.315 670.305 ;
        RECT 2090.765 669.990 2124.890 670.290 ;
        RECT 2090.765 669.975 2091.095 669.990 ;
        RECT 2027.950 669.310 2043.010 669.610 ;
        RECT 2124.590 669.610 2124.890 669.990 ;
        RECT 2139.310 669.990 2186.315 670.290 ;
        RECT 2139.310 669.610 2139.610 669.990 ;
        RECT 2185.985 669.975 2186.315 669.990 ;
        RECT 2187.825 670.290 2188.155 670.305 ;
        RECT 2187.825 669.990 2221.490 670.290 ;
        RECT 2187.825 669.975 2188.155 669.990 ;
        RECT 2124.590 669.310 2139.610 669.610 ;
        RECT 2221.190 669.610 2221.490 669.990 ;
        RECT 2235.910 669.610 2236.210 670.670 ;
        RECT 2282.585 670.655 2282.915 670.670 ;
        RECT 2287.185 670.290 2287.515 670.305 ;
        RECT 2377.805 670.290 2378.135 670.305 ;
        RECT 2287.185 669.990 2378.135 670.290 ;
        RECT 2287.185 669.975 2287.515 669.990 ;
        RECT 2377.805 669.975 2378.135 669.990 ;
        RECT 2414.605 670.290 2414.935 670.305 ;
        RECT 2415.310 670.290 2415.610 671.350 ;
        RECT 2438.985 671.335 2439.315 671.350 ;
        RECT 2463.110 670.970 2463.490 670.980 ;
        RECT 2463.110 670.670 2546.250 670.970 ;
        RECT 2463.110 670.660 2463.490 670.670 ;
        RECT 2414.605 669.990 2415.610 670.290 ;
        RECT 2545.950 670.290 2546.250 670.670 ;
        RECT 2594.710 670.670 2642.850 670.970 ;
        RECT 2545.950 669.990 2594.090 670.290 ;
        RECT 2414.605 669.975 2414.935 669.990 ;
        RECT 2221.190 669.310 2236.210 669.610 ;
        RECT 2438.985 669.610 2439.315 669.625 ;
        RECT 2463.110 669.610 2463.490 669.620 ;
        RECT 2438.985 669.310 2463.490 669.610 ;
        RECT 2593.790 669.610 2594.090 669.990 ;
        RECT 2594.710 669.610 2595.010 670.670 ;
        RECT 2642.550 670.290 2642.850 670.670 ;
        RECT 2691.310 670.670 2739.450 670.970 ;
        RECT 2642.550 669.990 2690.690 670.290 ;
        RECT 2593.790 669.310 2595.010 669.610 ;
        RECT 2690.390 669.610 2690.690 669.990 ;
        RECT 2691.310 669.610 2691.610 670.670 ;
        RECT 2739.150 670.290 2739.450 670.670 ;
        RECT 2787.910 670.670 2836.050 670.970 ;
        RECT 2739.150 669.990 2787.290 670.290 ;
        RECT 2690.390 669.310 2691.610 669.610 ;
        RECT 2786.990 669.610 2787.290 669.990 ;
        RECT 2787.910 669.610 2788.210 670.670 ;
        RECT 2835.750 670.290 2836.050 670.670 ;
        RECT 2916.710 670.290 2917.010 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
        RECT 2835.750 669.990 2883.890 670.290 ;
        RECT 2786.990 669.310 2788.210 669.610 ;
        RECT 2883.590 669.610 2883.890 669.990 ;
        RECT 2884.510 669.990 2917.010 670.290 ;
        RECT 2884.510 669.610 2884.810 669.990 ;
        RECT 2883.590 669.310 2884.810 669.610 ;
        RECT 1642.265 669.295 1642.595 669.310 ;
        RECT 2027.950 669.300 2028.330 669.310 ;
        RECT 2438.985 669.295 2439.315 669.310 ;
        RECT 2463.110 669.300 2463.490 669.310 ;
        RECT 1434.805 668.930 1435.135 668.945 ;
        RECT 1459.185 668.930 1459.515 668.945 ;
        RECT 1434.805 668.630 1459.515 668.930 ;
        RECT 1434.805 668.615 1435.135 668.630 ;
        RECT 1459.185 668.615 1459.515 668.630 ;
      LAYER via3 ;
        RECT 1226.660 2896.300 1226.980 2896.620 ;
        RECT 1290.140 672.700 1290.460 673.020 ;
        RECT 1226.660 670.660 1226.980 670.980 ;
        RECT 1290.140 670.660 1290.460 670.980 ;
        RECT 2027.980 670.660 2028.300 670.980 ;
        RECT 2027.980 669.300 2028.300 669.620 ;
        RECT 2463.140 670.660 2463.460 670.980 ;
        RECT 2463.140 669.300 2463.460 669.620 ;
      LAYER met4 ;
        RECT 1226.655 2896.295 1226.985 2896.625 ;
        RECT 1226.670 670.985 1226.970 2896.295 ;
        RECT 1290.135 672.695 1290.465 673.025 ;
        RECT 1290.150 670.985 1290.450 672.695 ;
        RECT 1226.655 670.655 1226.985 670.985 ;
        RECT 1290.135 670.655 1290.465 670.985 ;
        RECT 2027.975 670.655 2028.305 670.985 ;
        RECT 2463.135 670.655 2463.465 670.985 ;
        RECT 2027.990 669.625 2028.290 670.655 ;
        RECT 2463.150 669.625 2463.450 670.655 ;
        RECT 2027.975 669.295 2028.305 669.625 ;
        RECT 2463.135 669.295 2463.465 669.625 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 20.310 2913.700 20.630 2913.760 ;
        RECT 2111.930 2913.700 2112.250 2913.760 ;
        RECT 20.310 2913.560 2112.250 2913.700 ;
        RECT 20.310 2913.500 20.630 2913.560 ;
        RECT 2111.930 2913.500 2112.250 2913.560 ;
      LAYER via ;
        RECT 20.340 2913.500 20.600 2913.760 ;
        RECT 2111.960 2913.500 2112.220 2913.760 ;
      LAYER met2 ;
        RECT 20.340 2913.470 20.600 2913.790 ;
        RECT 2111.960 2913.470 2112.220 2913.790 ;
        RECT 20.400 1544.125 20.540 2913.470 ;
        RECT 2112.020 2900.000 2112.160 2913.470 ;
        RECT 2111.885 2896.000 2112.165 2900.000 ;
        RECT 20.330 1543.755 20.610 1544.125 ;
      LAYER via2 ;
        RECT 20.330 1543.800 20.610 1544.080 ;
      LAYER met3 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 20.305 1544.090 20.635 1544.105 ;
        RECT -4.800 1543.790 20.635 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 20.305 1543.775 20.635 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2141.905 2892.125 2142.075 2896.715 ;
      LAYER mcon ;
        RECT 2141.905 2896.545 2142.075 2896.715 ;
      LAYER met1 ;
        RECT 2141.830 2896.700 2142.150 2896.760 ;
        RECT 2141.635 2896.560 2142.150 2896.700 ;
        RECT 2141.830 2896.500 2142.150 2896.560 ;
        RECT 19.390 2892.280 19.710 2892.340 ;
        RECT 2141.845 2892.280 2142.135 2892.325 ;
        RECT 19.390 2892.140 2142.135 2892.280 ;
        RECT 19.390 2892.080 19.710 2892.140 ;
        RECT 2141.845 2892.095 2142.135 2892.140 ;
      LAYER via ;
        RECT 2141.860 2896.500 2142.120 2896.760 ;
        RECT 19.420 2892.080 19.680 2892.340 ;
      LAYER met2 ;
        RECT 2141.860 2896.530 2142.120 2896.790 ;
        RECT 2143.625 2896.530 2143.905 2900.000 ;
        RECT 2141.860 2896.470 2143.905 2896.530 ;
        RECT 2141.920 2896.390 2143.905 2896.470 ;
        RECT 2143.625 2896.000 2143.905 2896.390 ;
        RECT 19.420 2892.050 19.680 2892.370 ;
        RECT 19.480 1328.565 19.620 2892.050 ;
        RECT 19.410 1328.195 19.690 1328.565 ;
      LAYER via2 ;
        RECT 19.410 1328.240 19.690 1328.520 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 19.385 1328.530 19.715 1328.545 ;
        RECT -4.800 1328.230 19.715 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 19.385 1328.215 19.715 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 25.830 2912.680 26.150 2912.740 ;
        RECT 2174.950 2912.680 2175.270 2912.740 ;
        RECT 25.830 2912.540 2175.270 2912.680 ;
        RECT 25.830 2912.480 26.150 2912.540 ;
        RECT 2174.950 2912.480 2175.270 2912.540 ;
        RECT 13.870 1115.440 14.190 1115.500 ;
        RECT 25.830 1115.440 26.150 1115.500 ;
        RECT 13.870 1115.300 26.150 1115.440 ;
        RECT 13.870 1115.240 14.190 1115.300 ;
        RECT 25.830 1115.240 26.150 1115.300 ;
      LAYER via ;
        RECT 25.860 2912.480 26.120 2912.740 ;
        RECT 2174.980 2912.480 2175.240 2912.740 ;
        RECT 13.900 1115.240 14.160 1115.500 ;
        RECT 25.860 1115.240 26.120 1115.500 ;
      LAYER met2 ;
        RECT 25.860 2912.450 26.120 2912.770 ;
        RECT 2174.980 2912.450 2175.240 2912.770 ;
        RECT 25.920 1115.530 26.060 2912.450 ;
        RECT 2175.040 2900.000 2175.180 2912.450 ;
        RECT 2174.905 2896.000 2175.185 2900.000 ;
        RECT 13.900 1115.210 14.160 1115.530 ;
        RECT 25.860 1115.210 26.120 1115.530 ;
        RECT 13.960 1113.005 14.100 1115.210 ;
        RECT 13.890 1112.635 14.170 1113.005 ;
      LAYER via2 ;
        RECT 13.890 1112.680 14.170 1112.960 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 13.865 1112.970 14.195 1112.985 ;
        RECT -4.800 1112.670 14.195 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 13.865 1112.655 14.195 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2205.385 2891.785 2205.555 2896.715 ;
      LAYER mcon ;
        RECT 2205.385 2896.545 2205.555 2896.715 ;
      LAYER met1 ;
        RECT 2205.310 2896.700 2205.630 2896.760 ;
        RECT 2205.115 2896.560 2205.630 2896.700 ;
        RECT 2205.310 2896.500 2205.630 2896.560 ;
        RECT 18.010 2891.940 18.330 2892.000 ;
        RECT 2205.325 2891.940 2205.615 2891.985 ;
        RECT 18.010 2891.800 2205.615 2891.940 ;
        RECT 18.010 2891.740 18.330 2891.800 ;
        RECT 2205.325 2891.755 2205.615 2891.800 ;
      LAYER via ;
        RECT 2205.340 2896.500 2205.600 2896.760 ;
        RECT 18.040 2891.740 18.300 2892.000 ;
      LAYER met2 ;
        RECT 2205.340 2896.530 2205.600 2896.790 ;
        RECT 2206.645 2896.530 2206.925 2900.000 ;
        RECT 2205.340 2896.470 2206.925 2896.530 ;
        RECT 2205.400 2896.390 2206.925 2896.470 ;
        RECT 2206.645 2896.000 2206.925 2896.390 ;
        RECT 18.040 2891.710 18.300 2892.030 ;
        RECT 18.100 897.445 18.240 2891.710 ;
        RECT 18.030 897.075 18.310 897.445 ;
      LAYER via2 ;
        RECT 18.030 897.120 18.310 897.400 ;
      LAYER met3 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 18.005 897.410 18.335 897.425 ;
        RECT -4.800 897.110 18.335 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 18.005 897.095 18.335 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 25.370 2912.000 25.690 2912.060 ;
        RECT 2238.430 2912.000 2238.750 2912.060 ;
        RECT 25.370 2911.860 2238.750 2912.000 ;
        RECT 25.370 2911.800 25.690 2911.860 ;
        RECT 2238.430 2911.800 2238.750 2911.860 ;
        RECT 13.870 682.620 14.190 682.680 ;
        RECT 25.370 682.620 25.690 682.680 ;
        RECT 13.870 682.480 25.690 682.620 ;
        RECT 13.870 682.420 14.190 682.480 ;
        RECT 25.370 682.420 25.690 682.480 ;
      LAYER via ;
        RECT 25.400 2911.800 25.660 2912.060 ;
        RECT 2238.460 2911.800 2238.720 2912.060 ;
        RECT 13.900 682.420 14.160 682.680 ;
        RECT 25.400 682.420 25.660 682.680 ;
      LAYER met2 ;
        RECT 25.400 2911.770 25.660 2912.090 ;
        RECT 2238.460 2911.770 2238.720 2912.090 ;
        RECT 25.460 682.710 25.600 2911.770 ;
        RECT 2238.520 2900.000 2238.660 2911.770 ;
        RECT 2238.385 2896.000 2238.665 2900.000 ;
        RECT 13.900 682.390 14.160 682.710 ;
        RECT 25.400 682.390 25.660 682.710 ;
        RECT 13.960 681.885 14.100 682.390 ;
        RECT 13.890 681.515 14.170 681.885 ;
      LAYER via2 ;
        RECT 13.890 681.560 14.170 681.840 ;
      LAYER met3 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 13.865 681.850 14.195 681.865 ;
        RECT -4.800 681.550 14.195 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 13.865 681.535 14.195 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2267.945 2891.445 2268.115 2896.715 ;
      LAYER mcon ;
        RECT 2267.945 2896.545 2268.115 2896.715 ;
      LAYER met1 ;
        RECT 2267.870 2896.700 2268.190 2896.760 ;
        RECT 2267.675 2896.560 2268.190 2896.700 ;
        RECT 2267.870 2896.500 2268.190 2896.560 ;
        RECT 17.090 2891.600 17.410 2891.660 ;
        RECT 2267.885 2891.600 2268.175 2891.645 ;
        RECT 17.090 2891.460 2268.175 2891.600 ;
        RECT 17.090 2891.400 17.410 2891.460 ;
        RECT 2267.885 2891.415 2268.175 2891.460 ;
      LAYER via ;
        RECT 2267.900 2896.500 2268.160 2896.760 ;
        RECT 17.120 2891.400 17.380 2891.660 ;
      LAYER met2 ;
        RECT 2267.900 2896.530 2268.160 2896.790 ;
        RECT 2269.665 2896.530 2269.945 2900.000 ;
        RECT 2267.900 2896.470 2269.945 2896.530 ;
        RECT 2267.960 2896.390 2269.945 2896.470 ;
        RECT 2269.665 2896.000 2269.945 2896.390 ;
        RECT 17.120 2891.370 17.380 2891.690 ;
        RECT 17.180 466.325 17.320 2891.370 ;
        RECT 17.110 465.955 17.390 466.325 ;
      LAYER via2 ;
        RECT 17.110 466.000 17.390 466.280 ;
      LAYER met3 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.085 466.290 17.415 466.305 ;
        RECT -4.800 465.990 17.415 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.085 465.975 17.415 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 13.870 252.520 14.190 252.580 ;
        RECT 23.990 252.520 24.310 252.580 ;
        RECT 13.870 252.380 24.310 252.520 ;
        RECT 13.870 252.320 14.190 252.380 ;
        RECT 23.990 252.320 24.310 252.380 ;
      LAYER via ;
        RECT 13.900 252.320 14.160 252.580 ;
        RECT 24.020 252.320 24.280 252.580 ;
      LAYER met2 ;
        RECT 24.010 2916.675 24.290 2917.045 ;
        RECT 2301.470 2916.675 2301.750 2917.045 ;
        RECT 24.080 252.610 24.220 2916.675 ;
        RECT 2301.540 2900.000 2301.680 2916.675 ;
        RECT 2301.405 2896.000 2301.685 2900.000 ;
        RECT 13.900 252.290 14.160 252.610 ;
        RECT 24.020 252.290 24.280 252.610 ;
        RECT 13.960 250.765 14.100 252.290 ;
        RECT 13.890 250.395 14.170 250.765 ;
      LAYER via2 ;
        RECT 24.010 2916.720 24.290 2917.000 ;
        RECT 2301.470 2916.720 2301.750 2917.000 ;
        RECT 13.890 250.440 14.170 250.720 ;
      LAYER met3 ;
        RECT 23.985 2917.010 24.315 2917.025 ;
        RECT 2301.445 2917.010 2301.775 2917.025 ;
        RECT 23.985 2916.710 2301.775 2917.010 ;
        RECT 23.985 2916.695 24.315 2916.710 ;
        RECT 2301.445 2916.695 2301.775 2916.710 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 13.865 250.730 14.195 250.745 ;
        RECT -4.800 250.430 14.195 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 13.865 250.415 14.195 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2332.290 2896.530 2332.570 2896.645 ;
        RECT 2333.145 2896.530 2333.425 2900.000 ;
        RECT 2332.290 2896.390 2333.425 2896.530 ;
        RECT 2332.290 2896.275 2332.570 2896.390 ;
        RECT 2333.145 2896.000 2333.425 2896.390 ;
        RECT 15.730 57.955 16.010 58.325 ;
        RECT 15.800 35.885 15.940 57.955 ;
        RECT 15.730 35.515 16.010 35.885 ;
      LAYER via2 ;
        RECT 2332.290 2896.320 2332.570 2896.600 ;
        RECT 15.730 58.000 16.010 58.280 ;
        RECT 15.730 35.560 16.010 35.840 ;
      LAYER met3 ;
        RECT 2332.265 2896.620 2332.595 2896.625 ;
        RECT 2332.265 2896.610 2332.850 2896.620 ;
        RECT 2332.265 2896.310 2333.050 2896.610 ;
        RECT 2332.265 2896.300 2332.850 2896.310 ;
        RECT 2332.265 2896.295 2332.595 2896.300 ;
        RECT 15.705 58.290 16.035 58.305 ;
        RECT 2332.470 58.290 2332.850 58.300 ;
        RECT 15.705 57.990 2332.850 58.290 ;
        RECT 15.705 57.975 16.035 57.990 ;
        RECT 2332.470 57.980 2332.850 57.990 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 15.705 35.850 16.035 35.865 ;
        RECT -4.800 35.550 16.035 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 15.705 35.535 16.035 35.550 ;
      LAYER via3 ;
        RECT 2332.500 2896.300 2332.820 2896.620 ;
        RECT 2332.500 57.980 2332.820 58.300 ;
      LAYER met4 ;
        RECT 2332.495 2896.295 2332.825 2896.625 ;
        RECT 2332.510 58.305 2332.810 2896.295 ;
        RECT 2332.495 57.975 2332.825 58.305 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1259.090 2917.100 1259.410 2917.160 ;
        RECT 2901.750 2917.100 2902.070 2917.160 ;
        RECT 1259.090 2916.960 2902.070 2917.100 ;
        RECT 1259.090 2916.900 1259.410 2916.960 ;
        RECT 2901.750 2916.900 2902.070 2916.960 ;
      LAYER via ;
        RECT 1259.120 2916.900 1259.380 2917.160 ;
        RECT 2901.780 2916.900 2902.040 2917.160 ;
      LAYER met2 ;
        RECT 1259.120 2916.870 1259.380 2917.190 ;
        RECT 2901.780 2916.870 2902.040 2917.190 ;
        RECT 1259.180 2900.000 1259.320 2916.870 ;
        RECT 1259.045 2896.000 1259.325 2900.000 ;
        RECT 2901.840 909.685 2901.980 2916.870 ;
        RECT 2901.770 909.315 2902.050 909.685 ;
      LAYER via2 ;
        RECT 2901.770 909.360 2902.050 909.640 ;
      LAYER met3 ;
        RECT 2901.745 909.650 2902.075 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2901.745 909.350 2924.800 909.650 ;
        RECT 2901.745 909.335 2902.075 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1290.830 2905.200 1291.150 2905.260 ;
        RECT 2903.130 2905.200 2903.450 2905.260 ;
        RECT 1290.830 2905.060 2903.450 2905.200 ;
        RECT 1290.830 2905.000 1291.150 2905.060 ;
        RECT 2903.130 2905.000 2903.450 2905.060 ;
      LAYER via ;
        RECT 1290.860 2905.000 1291.120 2905.260 ;
        RECT 2903.160 2905.000 2903.420 2905.260 ;
      LAYER met2 ;
        RECT 1290.860 2904.970 1291.120 2905.290 ;
        RECT 2903.160 2904.970 2903.420 2905.290 ;
        RECT 1290.920 2900.000 1291.060 2904.970 ;
        RECT 1290.785 2896.000 1291.065 2900.000 ;
        RECT 2903.220 1144.285 2903.360 2904.970 ;
        RECT 2903.150 1143.915 2903.430 1144.285 ;
      LAYER via2 ;
        RECT 2903.150 1143.960 2903.430 1144.240 ;
      LAYER met3 ;
        RECT 2903.125 1144.250 2903.455 1144.265 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2903.125 1143.950 2924.800 1144.250 ;
        RECT 2903.125 1143.935 2903.455 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1322.570 2905.540 1322.890 2905.600 ;
        RECT 2904.510 2905.540 2904.830 2905.600 ;
        RECT 1322.570 2905.400 2904.830 2905.540 ;
        RECT 1322.570 2905.340 1322.890 2905.400 ;
        RECT 2904.510 2905.340 2904.830 2905.400 ;
        RECT 2898.990 2835.840 2899.310 2835.900 ;
        RECT 2904.510 2835.840 2904.830 2835.900 ;
        RECT 2898.990 2835.700 2904.830 2835.840 ;
        RECT 2898.990 2835.640 2899.310 2835.700 ;
        RECT 2904.510 2835.640 2904.830 2835.700 ;
        RECT 2898.990 2788.240 2899.310 2788.300 ;
        RECT 2898.990 2788.100 2904.740 2788.240 ;
        RECT 2898.990 2788.040 2899.310 2788.100 ;
        RECT 2904.600 2787.960 2904.740 2788.100 ;
        RECT 2904.510 2787.700 2904.830 2787.960 ;
        RECT 2898.530 2739.280 2898.850 2739.340 ;
        RECT 2904.510 2739.280 2904.830 2739.340 ;
        RECT 2898.530 2739.140 2904.830 2739.280 ;
        RECT 2898.530 2739.080 2898.850 2739.140 ;
        RECT 2904.510 2739.080 2904.830 2739.140 ;
        RECT 2898.530 2691.340 2898.850 2691.400 ;
        RECT 2904.510 2691.340 2904.830 2691.400 ;
        RECT 2898.530 2691.200 2904.830 2691.340 ;
        RECT 2898.530 2691.140 2898.850 2691.200 ;
        RECT 2904.510 2691.140 2904.830 2691.200 ;
        RECT 2898.990 2642.720 2899.310 2642.780 ;
        RECT 2904.510 2642.720 2904.830 2642.780 ;
        RECT 2898.990 2642.580 2904.830 2642.720 ;
        RECT 2898.990 2642.520 2899.310 2642.580 ;
        RECT 2904.510 2642.520 2904.830 2642.580 ;
        RECT 2898.990 2594.780 2899.310 2594.840 ;
        RECT 2904.510 2594.780 2904.830 2594.840 ;
        RECT 2898.990 2594.640 2904.830 2594.780 ;
        RECT 2898.990 2594.580 2899.310 2594.640 ;
        RECT 2904.510 2594.580 2904.830 2594.640 ;
        RECT 2898.990 2546.160 2899.310 2546.220 ;
        RECT 2904.510 2546.160 2904.830 2546.220 ;
        RECT 2898.990 2546.020 2904.830 2546.160 ;
        RECT 2898.990 2545.960 2899.310 2546.020 ;
        RECT 2904.510 2545.960 2904.830 2546.020 ;
        RECT 2898.990 2498.220 2899.310 2498.280 ;
        RECT 2898.990 2498.080 2904.740 2498.220 ;
        RECT 2898.990 2498.020 2899.310 2498.080 ;
        RECT 2904.600 2497.940 2904.740 2498.080 ;
        RECT 2904.510 2497.680 2904.830 2497.940 ;
        RECT 2898.990 2449.260 2899.310 2449.320 ;
        RECT 2904.510 2449.260 2904.830 2449.320 ;
        RECT 2898.990 2449.120 2904.830 2449.260 ;
        RECT 2898.990 2449.060 2899.310 2449.120 ;
        RECT 2904.510 2449.060 2904.830 2449.120 ;
        RECT 2898.990 2401.320 2899.310 2401.380 ;
        RECT 2904.510 2401.320 2904.830 2401.380 ;
        RECT 2898.990 2401.180 2904.830 2401.320 ;
        RECT 2898.990 2401.120 2899.310 2401.180 ;
        RECT 2904.510 2401.120 2904.830 2401.180 ;
        RECT 2898.530 2352.700 2898.850 2352.760 ;
        RECT 2904.510 2352.700 2904.830 2352.760 ;
        RECT 2898.530 2352.560 2904.830 2352.700 ;
        RECT 2898.530 2352.500 2898.850 2352.560 ;
        RECT 2904.510 2352.500 2904.830 2352.560 ;
        RECT 2898.530 2304.760 2898.850 2304.820 ;
        RECT 2904.510 2304.760 2904.830 2304.820 ;
        RECT 2898.530 2304.620 2904.830 2304.760 ;
        RECT 2898.530 2304.560 2898.850 2304.620 ;
        RECT 2904.510 2304.560 2904.830 2304.620 ;
        RECT 2898.990 2063.020 2899.310 2063.080 ;
        RECT 2904.510 2063.020 2904.830 2063.080 ;
        RECT 2898.990 2062.880 2904.830 2063.020 ;
        RECT 2898.990 2062.820 2899.310 2062.880 ;
        RECT 2904.510 2062.820 2904.830 2062.880 ;
        RECT 2898.990 2015.080 2899.310 2015.140 ;
        RECT 2904.510 2015.080 2904.830 2015.140 ;
        RECT 2898.990 2014.940 2904.830 2015.080 ;
        RECT 2898.990 2014.880 2899.310 2014.940 ;
        RECT 2904.510 2014.880 2904.830 2014.940 ;
        RECT 2904.510 1966.460 2904.830 1966.520 ;
        RECT 2900.000 1966.320 2904.830 1966.460 ;
        RECT 2898.990 1966.120 2899.310 1966.180 ;
        RECT 2900.000 1966.120 2900.140 1966.320 ;
        RECT 2904.510 1966.260 2904.830 1966.320 ;
        RECT 2898.990 1965.980 2900.140 1966.120 ;
        RECT 2898.990 1965.920 2899.310 1965.980 ;
        RECT 2898.990 1921.580 2899.310 1921.640 ;
        RECT 2904.510 1921.580 2904.830 1921.640 ;
        RECT 2898.990 1921.440 2904.830 1921.580 ;
        RECT 2898.990 1921.380 2899.310 1921.440 ;
        RECT 2904.510 1921.380 2904.830 1921.440 ;
        RECT 2899.910 1806.320 2900.230 1806.380 ;
        RECT 2904.510 1806.320 2904.830 1806.380 ;
        RECT 2899.910 1806.180 2904.830 1806.320 ;
        RECT 2899.910 1806.120 2900.230 1806.180 ;
        RECT 2904.510 1806.120 2904.830 1806.180 ;
        RECT 2898.990 1800.880 2899.310 1800.940 ;
        RECT 2899.910 1800.880 2900.230 1800.940 ;
        RECT 2898.990 1800.740 2900.230 1800.880 ;
        RECT 2898.990 1800.680 2899.310 1800.740 ;
        RECT 2899.910 1800.680 2900.230 1800.740 ;
        RECT 2900.370 1725.400 2900.690 1725.460 ;
        RECT 2904.510 1725.400 2904.830 1725.460 ;
        RECT 2900.370 1725.260 2904.830 1725.400 ;
        RECT 2900.370 1725.200 2900.690 1725.260 ;
        RECT 2904.510 1725.200 2904.830 1725.260 ;
        RECT 2900.370 1724.720 2900.690 1724.780 ;
        RECT 2904.510 1724.720 2904.830 1724.780 ;
        RECT 2900.370 1724.580 2904.830 1724.720 ;
        RECT 2900.370 1724.520 2900.690 1724.580 ;
        RECT 2904.510 1724.520 2904.830 1724.580 ;
        RECT 2900.370 1677.120 2900.690 1677.180 ;
        RECT 2904.970 1677.120 2905.290 1677.180 ;
        RECT 2900.370 1676.980 2905.290 1677.120 ;
        RECT 2900.370 1676.920 2900.690 1676.980 ;
        RECT 2904.970 1676.920 2905.290 1676.980 ;
        RECT 2900.370 1676.440 2900.690 1676.500 ;
        RECT 2904.970 1676.440 2905.290 1676.500 ;
        RECT 2900.370 1676.300 2905.290 1676.440 ;
        RECT 2900.370 1676.240 2900.690 1676.300 ;
        RECT 2904.970 1676.240 2905.290 1676.300 ;
        RECT 2900.370 1628.500 2900.690 1628.560 ;
        RECT 2904.510 1628.500 2904.830 1628.560 ;
        RECT 2900.370 1628.360 2904.830 1628.500 ;
        RECT 2900.370 1628.300 2900.690 1628.360 ;
        RECT 2904.510 1628.300 2904.830 1628.360 ;
        RECT 2899.910 1580.560 2900.230 1580.620 ;
        RECT 2904.970 1580.560 2905.290 1580.620 ;
        RECT 2899.910 1580.420 2905.290 1580.560 ;
        RECT 2899.910 1580.360 2900.230 1580.420 ;
        RECT 2904.970 1580.360 2905.290 1580.420 ;
        RECT 2900.370 1579.880 2900.690 1579.940 ;
        RECT 2904.970 1579.880 2905.290 1579.940 ;
        RECT 2900.370 1579.740 2905.290 1579.880 ;
        RECT 2900.370 1579.680 2900.690 1579.740 ;
        RECT 2904.970 1579.680 2905.290 1579.740 ;
        RECT 2900.370 1531.940 2900.690 1532.000 ;
        RECT 2904.510 1531.940 2904.830 1532.000 ;
        RECT 2900.370 1531.800 2904.830 1531.940 ;
        RECT 2900.370 1531.740 2900.690 1531.800 ;
        RECT 2904.510 1531.740 2904.830 1531.800 ;
        RECT 2900.370 1484.000 2900.690 1484.060 ;
        RECT 2904.970 1484.000 2905.290 1484.060 ;
        RECT 2900.370 1483.860 2905.290 1484.000 ;
        RECT 2900.370 1483.800 2900.690 1483.860 ;
        RECT 2904.970 1483.800 2905.290 1483.860 ;
        RECT 2900.830 1483.320 2901.150 1483.380 ;
        RECT 2904.970 1483.320 2905.290 1483.380 ;
        RECT 2900.830 1483.180 2905.290 1483.320 ;
        RECT 2900.830 1483.120 2901.150 1483.180 ;
        RECT 2904.970 1483.120 2905.290 1483.180 ;
        RECT 2900.830 1435.380 2901.150 1435.440 ;
        RECT 2904.510 1435.380 2904.830 1435.440 ;
        RECT 2900.830 1435.240 2904.830 1435.380 ;
        RECT 2900.830 1435.180 2901.150 1435.240 ;
        RECT 2904.510 1435.180 2904.830 1435.240 ;
        RECT 2900.830 1386.760 2901.150 1386.820 ;
        RECT 2904.510 1386.760 2904.830 1386.820 ;
        RECT 2900.830 1386.620 2904.830 1386.760 ;
        RECT 2900.830 1386.560 2901.150 1386.620 ;
        RECT 2904.510 1386.560 2904.830 1386.620 ;
      LAYER via ;
        RECT 1322.600 2905.340 1322.860 2905.600 ;
        RECT 2904.540 2905.340 2904.800 2905.600 ;
        RECT 2899.020 2835.640 2899.280 2835.900 ;
        RECT 2904.540 2835.640 2904.800 2835.900 ;
        RECT 2899.020 2788.040 2899.280 2788.300 ;
        RECT 2904.540 2787.700 2904.800 2787.960 ;
        RECT 2898.560 2739.080 2898.820 2739.340 ;
        RECT 2904.540 2739.080 2904.800 2739.340 ;
        RECT 2898.560 2691.140 2898.820 2691.400 ;
        RECT 2904.540 2691.140 2904.800 2691.400 ;
        RECT 2899.020 2642.520 2899.280 2642.780 ;
        RECT 2904.540 2642.520 2904.800 2642.780 ;
        RECT 2899.020 2594.580 2899.280 2594.840 ;
        RECT 2904.540 2594.580 2904.800 2594.840 ;
        RECT 2899.020 2545.960 2899.280 2546.220 ;
        RECT 2904.540 2545.960 2904.800 2546.220 ;
        RECT 2899.020 2498.020 2899.280 2498.280 ;
        RECT 2904.540 2497.680 2904.800 2497.940 ;
        RECT 2899.020 2449.060 2899.280 2449.320 ;
        RECT 2904.540 2449.060 2904.800 2449.320 ;
        RECT 2899.020 2401.120 2899.280 2401.380 ;
        RECT 2904.540 2401.120 2904.800 2401.380 ;
        RECT 2898.560 2352.500 2898.820 2352.760 ;
        RECT 2904.540 2352.500 2904.800 2352.760 ;
        RECT 2898.560 2304.560 2898.820 2304.820 ;
        RECT 2904.540 2304.560 2904.800 2304.820 ;
        RECT 2899.020 2062.820 2899.280 2063.080 ;
        RECT 2904.540 2062.820 2904.800 2063.080 ;
        RECT 2899.020 2014.880 2899.280 2015.140 ;
        RECT 2904.540 2014.880 2904.800 2015.140 ;
        RECT 2899.020 1965.920 2899.280 1966.180 ;
        RECT 2904.540 1966.260 2904.800 1966.520 ;
        RECT 2899.020 1921.380 2899.280 1921.640 ;
        RECT 2904.540 1921.380 2904.800 1921.640 ;
        RECT 2899.940 1806.120 2900.200 1806.380 ;
        RECT 2904.540 1806.120 2904.800 1806.380 ;
        RECT 2899.020 1800.680 2899.280 1800.940 ;
        RECT 2899.940 1800.680 2900.200 1800.940 ;
        RECT 2900.400 1725.200 2900.660 1725.460 ;
        RECT 2904.540 1725.200 2904.800 1725.460 ;
        RECT 2900.400 1724.520 2900.660 1724.780 ;
        RECT 2904.540 1724.520 2904.800 1724.780 ;
        RECT 2900.400 1676.920 2900.660 1677.180 ;
        RECT 2905.000 1676.920 2905.260 1677.180 ;
        RECT 2900.400 1676.240 2900.660 1676.500 ;
        RECT 2905.000 1676.240 2905.260 1676.500 ;
        RECT 2900.400 1628.300 2900.660 1628.560 ;
        RECT 2904.540 1628.300 2904.800 1628.560 ;
        RECT 2899.940 1580.360 2900.200 1580.620 ;
        RECT 2905.000 1580.360 2905.260 1580.620 ;
        RECT 2900.400 1579.680 2900.660 1579.940 ;
        RECT 2905.000 1579.680 2905.260 1579.940 ;
        RECT 2900.400 1531.740 2900.660 1532.000 ;
        RECT 2904.540 1531.740 2904.800 1532.000 ;
        RECT 2900.400 1483.800 2900.660 1484.060 ;
        RECT 2905.000 1483.800 2905.260 1484.060 ;
        RECT 2900.860 1483.120 2901.120 1483.380 ;
        RECT 2905.000 1483.120 2905.260 1483.380 ;
        RECT 2900.860 1435.180 2901.120 1435.440 ;
        RECT 2904.540 1435.180 2904.800 1435.440 ;
        RECT 2900.860 1386.560 2901.120 1386.820 ;
        RECT 2904.540 1386.560 2904.800 1386.820 ;
      LAYER met2 ;
        RECT 1322.600 2905.310 1322.860 2905.630 ;
        RECT 2904.540 2905.310 2904.800 2905.630 ;
        RECT 1322.660 2900.000 1322.800 2905.310 ;
        RECT 1322.525 2896.000 1322.805 2900.000 ;
        RECT 2904.600 2835.930 2904.740 2905.310 ;
        RECT 2899.020 2835.610 2899.280 2835.930 ;
        RECT 2904.540 2835.610 2904.800 2835.930 ;
        RECT 2899.080 2788.330 2899.220 2835.610 ;
        RECT 2899.020 2788.010 2899.280 2788.330 ;
        RECT 2904.540 2787.670 2904.800 2787.990 ;
        RECT 2904.600 2739.370 2904.740 2787.670 ;
        RECT 2898.560 2739.050 2898.820 2739.370 ;
        RECT 2904.540 2739.050 2904.800 2739.370 ;
        RECT 2898.620 2691.430 2898.760 2739.050 ;
        RECT 2898.560 2691.110 2898.820 2691.430 ;
        RECT 2904.540 2691.110 2904.800 2691.430 ;
        RECT 2904.600 2642.810 2904.740 2691.110 ;
        RECT 2899.020 2642.490 2899.280 2642.810 ;
        RECT 2904.540 2642.490 2904.800 2642.810 ;
        RECT 2899.080 2594.870 2899.220 2642.490 ;
        RECT 2899.020 2594.550 2899.280 2594.870 ;
        RECT 2904.540 2594.550 2904.800 2594.870 ;
        RECT 2904.600 2546.250 2904.740 2594.550 ;
        RECT 2899.020 2545.930 2899.280 2546.250 ;
        RECT 2904.540 2545.930 2904.800 2546.250 ;
        RECT 2899.080 2498.310 2899.220 2545.930 ;
        RECT 2899.020 2497.990 2899.280 2498.310 ;
        RECT 2904.540 2497.650 2904.800 2497.970 ;
        RECT 2904.600 2449.350 2904.740 2497.650 ;
        RECT 2899.020 2449.030 2899.280 2449.350 ;
        RECT 2904.540 2449.030 2904.800 2449.350 ;
        RECT 2899.080 2401.410 2899.220 2449.030 ;
        RECT 2899.020 2401.090 2899.280 2401.410 ;
        RECT 2904.540 2401.090 2904.800 2401.410 ;
        RECT 2904.600 2352.790 2904.740 2401.090 ;
        RECT 2898.560 2352.470 2898.820 2352.790 ;
        RECT 2904.540 2352.470 2904.800 2352.790 ;
        RECT 2898.620 2304.850 2898.760 2352.470 ;
        RECT 2898.560 2304.530 2898.820 2304.850 ;
        RECT 2904.540 2304.530 2904.800 2304.850 ;
        RECT 2904.600 2063.110 2904.740 2304.530 ;
        RECT 2899.020 2062.790 2899.280 2063.110 ;
        RECT 2904.540 2062.790 2904.800 2063.110 ;
        RECT 2899.080 2015.170 2899.220 2062.790 ;
        RECT 2899.020 2014.850 2899.280 2015.170 ;
        RECT 2904.540 2014.850 2904.800 2015.170 ;
        RECT 2904.600 1966.550 2904.740 2014.850 ;
        RECT 2904.540 1966.230 2904.800 1966.550 ;
        RECT 2899.020 1965.890 2899.280 1966.210 ;
        RECT 2899.080 1921.670 2899.220 1965.890 ;
        RECT 2899.020 1921.350 2899.280 1921.670 ;
        RECT 2904.540 1921.350 2904.800 1921.670 ;
        RECT 2904.600 1806.410 2904.740 1921.350 ;
        RECT 2899.940 1806.090 2900.200 1806.410 ;
        RECT 2904.540 1806.090 2904.800 1806.410 ;
        RECT 2900.000 1800.970 2900.140 1806.090 ;
        RECT 2899.020 1800.650 2899.280 1800.970 ;
        RECT 2899.940 1800.650 2900.200 1800.970 ;
        RECT 2899.080 1788.130 2899.220 1800.650 ;
        RECT 2899.080 1787.990 2900.600 1788.130 ;
        RECT 2900.460 1725.490 2900.600 1787.990 ;
        RECT 2900.400 1725.170 2900.660 1725.490 ;
        RECT 2904.540 1725.170 2904.800 1725.490 ;
        RECT 2904.600 1724.810 2904.740 1725.170 ;
        RECT 2900.400 1724.490 2900.660 1724.810 ;
        RECT 2904.540 1724.490 2904.800 1724.810 ;
        RECT 2900.460 1677.210 2900.600 1724.490 ;
        RECT 2900.400 1676.890 2900.660 1677.210 ;
        RECT 2905.000 1676.890 2905.260 1677.210 ;
        RECT 2905.060 1676.530 2905.200 1676.890 ;
        RECT 2900.400 1676.210 2900.660 1676.530 ;
        RECT 2905.000 1676.210 2905.260 1676.530 ;
        RECT 2900.460 1628.590 2900.600 1676.210 ;
        RECT 2899.930 1628.075 2900.210 1628.445 ;
        RECT 2900.400 1628.270 2900.660 1628.590 ;
        RECT 2904.540 1628.445 2904.800 1628.590 ;
        RECT 2904.530 1628.075 2904.810 1628.445 ;
        RECT 2900.000 1580.650 2900.140 1628.075 ;
        RECT 2899.940 1580.330 2900.200 1580.650 ;
        RECT 2905.000 1580.330 2905.260 1580.650 ;
        RECT 2905.060 1579.970 2905.200 1580.330 ;
        RECT 2900.400 1579.650 2900.660 1579.970 ;
        RECT 2905.000 1579.650 2905.260 1579.970 ;
        RECT 2900.460 1532.030 2900.600 1579.650 ;
        RECT 2900.400 1531.885 2900.660 1532.030 ;
        RECT 2904.540 1531.885 2904.800 1532.030 ;
        RECT 2900.390 1531.515 2900.670 1531.885 ;
        RECT 2904.530 1531.515 2904.810 1531.885 ;
        RECT 2900.460 1484.090 2900.600 1531.515 ;
        RECT 2900.400 1483.770 2900.660 1484.090 ;
        RECT 2905.000 1483.770 2905.260 1484.090 ;
        RECT 2905.060 1483.410 2905.200 1483.770 ;
        RECT 2900.860 1483.090 2901.120 1483.410 ;
        RECT 2905.000 1483.090 2905.260 1483.410 ;
        RECT 2900.920 1435.470 2901.060 1483.090 ;
        RECT 2900.860 1435.150 2901.120 1435.470 ;
        RECT 2904.540 1435.150 2904.800 1435.470 ;
        RECT 2904.600 1386.850 2904.740 1435.150 ;
        RECT 2900.860 1386.530 2901.120 1386.850 ;
        RECT 2904.540 1386.530 2904.800 1386.850 ;
        RECT 2900.920 1378.885 2901.060 1386.530 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 2899.930 1628.120 2900.210 1628.400 ;
        RECT 2904.530 1628.120 2904.810 1628.400 ;
        RECT 2900.390 1531.560 2900.670 1531.840 ;
        RECT 2904.530 1531.560 2904.810 1531.840 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 2899.905 1628.410 2900.235 1628.425 ;
        RECT 2904.505 1628.410 2904.835 1628.425 ;
        RECT 2899.905 1628.110 2904.835 1628.410 ;
        RECT 2899.905 1628.095 2900.235 1628.110 ;
        RECT 2904.505 1628.095 2904.835 1628.110 ;
        RECT 2900.365 1531.850 2900.695 1531.865 ;
        RECT 2904.505 1531.850 2904.835 1531.865 ;
        RECT 2900.365 1531.550 2904.835 1531.850 ;
        RECT 2900.365 1531.535 2900.695 1531.550 ;
        RECT 2904.505 1531.535 2904.835 1531.550 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1355.690 2897.040 1356.010 2897.100 ;
        RECT 1355.690 2896.900 1411.120 2897.040 ;
        RECT 1355.690 2896.840 1356.010 2896.900 ;
        RECT 1410.980 2895.680 1411.120 2896.900 ;
        RECT 2349.750 2895.680 2350.070 2895.740 ;
        RECT 1410.980 2895.540 2350.070 2895.680 ;
        RECT 2349.750 2895.480 2350.070 2895.540 ;
        RECT 2349.750 1614.560 2350.070 1614.620 ;
        RECT 2900.370 1614.560 2900.690 1614.620 ;
        RECT 2349.750 1614.420 2900.690 1614.560 ;
        RECT 2349.750 1614.360 2350.070 1614.420 ;
        RECT 2900.370 1614.360 2900.690 1614.420 ;
      LAYER via ;
        RECT 1355.720 2896.840 1355.980 2897.100 ;
        RECT 2349.780 2895.480 2350.040 2895.740 ;
        RECT 2349.780 1614.360 2350.040 1614.620 ;
        RECT 2900.400 1614.360 2900.660 1614.620 ;
      LAYER met2 ;
        RECT 1353.805 2897.210 1354.085 2900.000 ;
        RECT 1353.805 2897.130 1355.920 2897.210 ;
        RECT 1353.805 2897.070 1355.980 2897.130 ;
        RECT 1353.805 2896.000 1354.085 2897.070 ;
        RECT 1355.720 2896.810 1355.980 2897.070 ;
        RECT 2349.780 2895.450 2350.040 2895.770 ;
        RECT 2349.840 1614.650 2349.980 2895.450 ;
        RECT 2349.780 1614.330 2350.040 1614.650 ;
        RECT 2900.400 1614.330 2900.660 1614.650 ;
        RECT 2900.460 1613.485 2900.600 1614.330 ;
        RECT 2900.390 1613.115 2900.670 1613.485 ;
      LAYER via2 ;
        RECT 2900.390 1613.160 2900.670 1613.440 ;
      LAYER met3 ;
        RECT 2900.365 1613.450 2900.695 1613.465 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2900.365 1613.150 2924.800 1613.450 ;
        RECT 2900.365 1613.135 2900.695 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1386.510 2896.500 1386.830 2896.760 ;
        RECT 1386.600 2894.660 1386.740 2896.500 ;
        RECT 2899.910 2894.660 2900.230 2894.720 ;
        RECT 1386.600 2894.520 2900.230 2894.660 ;
        RECT 2899.910 2894.460 2900.230 2894.520 ;
      LAYER via ;
        RECT 1386.540 2896.500 1386.800 2896.760 ;
        RECT 2899.940 2894.460 2900.200 2894.720 ;
      LAYER met2 ;
        RECT 1385.545 2896.530 1385.825 2900.000 ;
        RECT 1386.540 2896.530 1386.800 2896.790 ;
        RECT 1385.545 2896.470 1386.800 2896.530 ;
        RECT 1385.545 2896.390 1386.740 2896.470 ;
        RECT 1385.545 2896.000 1385.825 2896.390 ;
        RECT 2899.940 2894.430 2900.200 2894.750 ;
        RECT 2900.000 1848.085 2900.140 2894.430 ;
        RECT 2899.930 1847.715 2900.210 1848.085 ;
      LAYER via2 ;
        RECT 2899.930 1847.760 2900.210 1848.040 ;
      LAYER met3 ;
        RECT 2899.905 1848.050 2900.235 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2899.905 1847.750 2924.800 1848.050 ;
        RECT 2899.905 1847.735 2900.235 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1417.330 2906.560 1417.650 2906.620 ;
        RECT 2351.590 2906.560 2351.910 2906.620 ;
        RECT 1417.330 2906.420 2351.910 2906.560 ;
        RECT 1417.330 2906.360 1417.650 2906.420 ;
        RECT 2351.590 2906.360 2351.910 2906.420 ;
        RECT 2351.590 2083.760 2351.910 2083.820 ;
        RECT 2899.450 2083.760 2899.770 2083.820 ;
        RECT 2351.590 2083.620 2899.770 2083.760 ;
        RECT 2351.590 2083.560 2351.910 2083.620 ;
        RECT 2899.450 2083.560 2899.770 2083.620 ;
      LAYER via ;
        RECT 1417.360 2906.360 1417.620 2906.620 ;
        RECT 2351.620 2906.360 2351.880 2906.620 ;
        RECT 2351.620 2083.560 2351.880 2083.820 ;
        RECT 2899.480 2083.560 2899.740 2083.820 ;
      LAYER met2 ;
        RECT 1417.360 2906.330 1417.620 2906.650 ;
        RECT 2351.620 2906.330 2351.880 2906.650 ;
        RECT 1417.420 2900.000 1417.560 2906.330 ;
        RECT 1417.285 2896.000 1417.565 2900.000 ;
        RECT 2351.680 2083.850 2351.820 2906.330 ;
        RECT 2351.620 2083.530 2351.880 2083.850 ;
        RECT 2899.480 2083.530 2899.740 2083.850 ;
        RECT 2899.540 2082.685 2899.680 2083.530 ;
        RECT 2899.470 2082.315 2899.750 2082.685 ;
      LAYER via2 ;
        RECT 2899.470 2082.360 2899.750 2082.640 ;
      LAYER met3 ;
        RECT 2899.445 2082.650 2899.775 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2899.445 2082.350 2924.800 2082.650 ;
        RECT 2899.445 2082.335 2899.775 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1448.610 2907.240 1448.930 2907.300 ;
        RECT 2352.510 2907.240 2352.830 2907.300 ;
        RECT 1448.610 2907.100 2352.830 2907.240 ;
        RECT 1448.610 2907.040 1448.930 2907.100 ;
        RECT 2352.510 2907.040 2352.830 2907.100 ;
        RECT 2352.510 2318.360 2352.830 2318.420 ;
        RECT 2898.990 2318.360 2899.310 2318.420 ;
        RECT 2352.510 2318.220 2899.310 2318.360 ;
        RECT 2352.510 2318.160 2352.830 2318.220 ;
        RECT 2898.990 2318.160 2899.310 2318.220 ;
      LAYER via ;
        RECT 1448.640 2907.040 1448.900 2907.300 ;
        RECT 2352.540 2907.040 2352.800 2907.300 ;
        RECT 2352.540 2318.160 2352.800 2318.420 ;
        RECT 2899.020 2318.160 2899.280 2318.420 ;
      LAYER met2 ;
        RECT 1448.640 2907.010 1448.900 2907.330 ;
        RECT 2352.540 2907.010 2352.800 2907.330 ;
        RECT 1448.700 2900.000 1448.840 2907.010 ;
        RECT 1448.565 2896.000 1448.845 2900.000 ;
        RECT 2352.600 2318.450 2352.740 2907.010 ;
        RECT 2352.540 2318.130 2352.800 2318.450 ;
        RECT 2899.020 2318.130 2899.280 2318.450 ;
        RECT 2899.080 2317.285 2899.220 2318.130 ;
        RECT 2899.010 2316.915 2899.290 2317.285 ;
      LAYER via2 ;
        RECT 2899.010 2316.960 2899.290 2317.240 ;
      LAYER met3 ;
        RECT 2898.985 2317.250 2899.315 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2898.985 2316.950 2924.800 2317.250 ;
        RECT 2898.985 2316.935 2899.315 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1265.530 146.100 1265.850 146.160 ;
        RECT 1289.910 146.100 1290.230 146.160 ;
        RECT 1265.530 145.960 1290.230 146.100 ;
        RECT 1265.530 145.900 1265.850 145.960 ;
        RECT 1289.910 145.900 1290.230 145.960 ;
        RECT 2185.990 146.100 2186.310 146.160 ;
        RECT 2187.370 146.100 2187.690 146.160 ;
        RECT 2185.990 145.960 2187.690 146.100 ;
        RECT 2185.990 145.900 2186.310 145.960 ;
        RECT 2187.370 145.900 2187.690 145.960 ;
        RECT 2326.290 146.100 2326.610 146.160 ;
        RECT 2339.630 146.100 2339.950 146.160 ;
        RECT 2326.290 145.960 2339.950 146.100 ;
        RECT 2326.290 145.900 2326.610 145.960 ;
        RECT 2339.630 145.900 2339.950 145.960 ;
        RECT 2089.390 145.760 2089.710 145.820 ;
        RECT 2090.770 145.760 2091.090 145.820 ;
        RECT 2089.390 145.620 2091.090 145.760 ;
        RECT 2089.390 145.560 2089.710 145.620 ;
        RECT 2090.770 145.560 2091.090 145.620 ;
        RECT 2463.830 145.420 2464.150 145.480 ;
        RECT 2511.210 145.420 2511.530 145.480 ;
        RECT 2463.830 145.280 2511.530 145.420 ;
        RECT 2463.830 145.220 2464.150 145.280 ;
        RECT 2511.210 145.220 2511.530 145.280 ;
        RECT 1531.410 144.740 1531.730 144.800 ;
        RECT 1572.810 144.740 1573.130 144.800 ;
        RECT 1531.410 144.600 1573.130 144.740 ;
        RECT 1531.410 144.540 1531.730 144.600 ;
        RECT 1572.810 144.540 1573.130 144.600 ;
      LAYER via ;
        RECT 1265.560 145.900 1265.820 146.160 ;
        RECT 1289.940 145.900 1290.200 146.160 ;
        RECT 2186.020 145.900 2186.280 146.160 ;
        RECT 2187.400 145.900 2187.660 146.160 ;
        RECT 2326.320 145.900 2326.580 146.160 ;
        RECT 2339.660 145.900 2339.920 146.160 ;
        RECT 2089.420 145.560 2089.680 145.820 ;
        RECT 2090.800 145.560 2091.060 145.820 ;
        RECT 2463.860 145.220 2464.120 145.480 ;
        RECT 2511.240 145.220 2511.500 145.480 ;
        RECT 1531.440 144.540 1531.700 144.800 ;
        RECT 1572.840 144.540 1573.100 144.800 ;
      LAYER met2 ;
        RECT 1174.865 2896.530 1175.145 2900.000 ;
        RECT 1176.310 2896.530 1176.590 2896.645 ;
        RECT 1174.865 2896.390 1176.590 2896.530 ;
        RECT 1174.865 2896.000 1175.145 2896.390 ;
        RECT 1176.310 2896.275 1176.590 2896.390 ;
        RECT 2456.030 147.035 2456.310 147.405 ;
        RECT 1265.550 146.355 1265.830 146.725 ;
        RECT 1634.930 146.355 1635.210 146.725 ;
        RECT 1683.230 146.355 1683.510 146.725 ;
        RECT 2339.650 146.355 2339.930 146.725 ;
        RECT 2380.130 146.355 2380.410 146.725 ;
        RECT 1265.620 146.190 1265.760 146.355 ;
        RECT 1265.560 145.870 1265.820 146.190 ;
        RECT 1289.940 146.045 1290.200 146.190 ;
        RECT 1289.930 145.675 1290.210 146.045 ;
        RECT 1365.370 145.930 1365.650 146.045 ;
        RECT 1366.290 145.930 1366.570 146.045 ;
        RECT 1365.370 145.790 1366.570 145.930 ;
        RECT 1365.370 145.675 1365.650 145.790 ;
        RECT 1366.290 145.675 1366.570 145.790 ;
        RECT 1628.030 145.675 1628.310 146.045 ;
        RECT 1531.440 144.685 1531.700 144.830 ;
        RECT 1572.840 144.685 1573.100 144.830 ;
        RECT 1628.100 144.685 1628.240 145.675 ;
        RECT 1635.000 144.685 1635.140 146.355 ;
        RECT 1683.300 145.365 1683.440 146.355 ;
        RECT 2339.720 146.190 2339.860 146.355 ;
        RECT 2186.020 146.045 2186.280 146.190 ;
        RECT 2187.400 146.045 2187.660 146.190 ;
        RECT 2326.320 146.045 2326.580 146.190 ;
        RECT 1835.490 145.675 1835.770 146.045 ;
        RECT 2089.410 145.675 2089.690 146.045 ;
        RECT 2090.790 145.675 2091.070 146.045 ;
        RECT 2186.010 145.675 2186.290 146.045 ;
        RECT 2187.390 145.675 2187.670 146.045 ;
        RECT 2326.310 145.675 2326.590 146.045 ;
        RECT 2339.660 145.870 2339.920 146.190 ;
        RECT 2380.200 145.930 2380.340 146.355 ;
        RECT 2381.050 145.930 2381.330 146.045 ;
        RECT 2380.200 145.790 2381.330 145.930 ;
        RECT 2381.050 145.675 2381.330 145.790 ;
        RECT 1835.560 145.365 1835.700 145.675 ;
        RECT 2089.420 145.530 2089.680 145.675 ;
        RECT 2090.800 145.530 2091.060 145.675 ;
        RECT 2456.100 145.365 2456.240 147.035 ;
        RECT 2511.230 146.355 2511.510 146.725 ;
        RECT 2511.300 145.510 2511.440 146.355 ;
        RECT 2463.860 145.365 2464.120 145.510 ;
        RECT 1683.230 144.995 1683.510 145.365 ;
        RECT 1835.490 144.995 1835.770 145.365 ;
        RECT 2456.030 144.995 2456.310 145.365 ;
        RECT 2463.850 144.995 2464.130 145.365 ;
        RECT 2511.240 145.190 2511.500 145.510 ;
        RECT 1531.430 144.315 1531.710 144.685 ;
        RECT 1572.830 144.315 1573.110 144.685 ;
        RECT 1628.030 144.315 1628.310 144.685 ;
        RECT 1634.930 144.315 1635.210 144.685 ;
      LAYER via2 ;
        RECT 1176.310 2896.320 1176.590 2896.600 ;
        RECT 2456.030 147.080 2456.310 147.360 ;
        RECT 1265.550 146.400 1265.830 146.680 ;
        RECT 1634.930 146.400 1635.210 146.680 ;
        RECT 1683.230 146.400 1683.510 146.680 ;
        RECT 2339.650 146.400 2339.930 146.680 ;
        RECT 2380.130 146.400 2380.410 146.680 ;
        RECT 1289.930 145.720 1290.210 146.000 ;
        RECT 1365.370 145.720 1365.650 146.000 ;
        RECT 1366.290 145.720 1366.570 146.000 ;
        RECT 1628.030 145.720 1628.310 146.000 ;
        RECT 1835.490 145.720 1835.770 146.000 ;
        RECT 2089.410 145.720 2089.690 146.000 ;
        RECT 2090.790 145.720 2091.070 146.000 ;
        RECT 2186.010 145.720 2186.290 146.000 ;
        RECT 2187.390 145.720 2187.670 146.000 ;
        RECT 2326.310 145.720 2326.590 146.000 ;
        RECT 2381.050 145.720 2381.330 146.000 ;
        RECT 2511.230 146.400 2511.510 146.680 ;
        RECT 1683.230 145.040 1683.510 145.320 ;
        RECT 1835.490 145.040 1835.770 145.320 ;
        RECT 2456.030 145.040 2456.310 145.320 ;
        RECT 2463.850 145.040 2464.130 145.320 ;
        RECT 1531.430 144.360 1531.710 144.640 ;
        RECT 1572.830 144.360 1573.110 144.640 ;
        RECT 1628.030 144.360 1628.310 144.640 ;
        RECT 1634.930 144.360 1635.210 144.640 ;
      LAYER met3 ;
        RECT 1176.285 2896.610 1176.615 2896.625 ;
        RECT 1178.790 2896.610 1179.170 2896.620 ;
        RECT 1176.285 2896.310 1179.170 2896.610 ;
        RECT 1176.285 2896.295 1176.615 2896.310 ;
        RECT 1178.790 2896.300 1179.170 2896.310 ;
        RECT 2027.950 147.370 2028.330 147.380 ;
        RECT 1993.030 147.070 2028.330 147.370 ;
        RECT 1178.790 146.690 1179.170 146.700 ;
        RECT 1265.525 146.690 1265.855 146.705 ;
        RECT 1634.905 146.700 1635.235 146.705 ;
        RECT 1634.905 146.690 1635.490 146.700 ;
        RECT 1178.790 146.390 1265.855 146.690 ;
        RECT 1178.790 146.380 1179.170 146.390 ;
        RECT 1265.525 146.375 1265.855 146.390 ;
        RECT 1369.270 146.390 1394.410 146.690 ;
        RECT 1634.700 146.390 1635.490 146.690 ;
        RECT 1289.905 146.010 1290.235 146.025 ;
        RECT 1365.345 146.010 1365.675 146.025 ;
        RECT 1289.905 145.710 1365.675 146.010 ;
        RECT 1289.905 145.695 1290.235 145.710 ;
        RECT 1365.345 145.695 1365.675 145.710 ;
        RECT 1366.265 146.010 1366.595 146.025 ;
        RECT 1369.270 146.010 1369.570 146.390 ;
        RECT 1366.265 145.710 1369.570 146.010 ;
        RECT 1394.110 146.010 1394.410 146.390 ;
        RECT 1634.905 146.380 1635.490 146.390 ;
        RECT 1683.205 146.690 1683.535 146.705 ;
        RECT 1683.205 146.390 1704.450 146.690 ;
        RECT 1634.905 146.375 1635.235 146.380 ;
        RECT 1683.205 146.375 1683.535 146.390 ;
        RECT 1435.470 146.010 1435.850 146.020 ;
        RECT 1628.005 146.010 1628.335 146.025 ;
        RECT 1394.110 145.710 1435.850 146.010 ;
        RECT 1366.265 145.695 1366.595 145.710 ;
        RECT 1435.470 145.700 1435.850 145.710 ;
        RECT 1580.870 145.710 1628.335 146.010 ;
        RECT 1580.870 144.820 1581.170 145.710 ;
        RECT 1628.005 145.695 1628.335 145.710 ;
        RECT 1635.110 145.330 1635.490 145.340 ;
        RECT 1683.205 145.330 1683.535 145.345 ;
        RECT 1635.110 145.030 1683.535 145.330 ;
        RECT 1704.150 145.330 1704.450 146.390 ;
        RECT 1835.710 146.390 1897.650 146.690 ;
        RECT 1835.710 146.025 1836.010 146.390 ;
        RECT 1752.910 145.710 1811.170 146.010 ;
        RECT 1752.910 145.330 1753.210 145.710 ;
        RECT 1704.150 145.030 1753.210 145.330 ;
        RECT 1810.870 145.330 1811.170 145.710 ;
        RECT 1835.465 145.710 1836.010 146.025 ;
        RECT 1835.465 145.695 1835.795 145.710 ;
        RECT 1835.465 145.330 1835.795 145.345 ;
        RECT 1810.870 145.030 1835.795 145.330 ;
        RECT 1897.350 145.330 1897.650 146.390 ;
        RECT 1993.030 146.010 1993.330 147.070 ;
        RECT 2027.950 147.060 2028.330 147.070 ;
        RECT 2407.910 147.370 2408.290 147.380 ;
        RECT 2456.005 147.370 2456.335 147.385 ;
        RECT 2407.910 147.070 2456.335 147.370 ;
        RECT 2407.910 147.060 2408.290 147.070 ;
        RECT 2456.005 147.055 2456.335 147.070 ;
        RECT 2339.625 146.690 2339.955 146.705 ;
        RECT 2380.105 146.690 2380.435 146.705 ;
        RECT 2235.910 146.390 2318.090 146.690 ;
        RECT 2089.385 146.010 2089.715 146.025 ;
        RECT 1946.110 145.710 1993.330 146.010 ;
        RECT 2042.710 145.710 2089.715 146.010 ;
        RECT 1946.110 145.330 1946.410 145.710 ;
        RECT 1897.350 145.030 1946.410 145.330 ;
        RECT 2027.950 145.330 2028.330 145.340 ;
        RECT 2042.710 145.330 2043.010 145.710 ;
        RECT 2089.385 145.695 2089.715 145.710 ;
        RECT 2090.765 146.010 2091.095 146.025 ;
        RECT 2185.985 146.010 2186.315 146.025 ;
        RECT 2090.765 145.710 2124.890 146.010 ;
        RECT 2090.765 145.695 2091.095 145.710 ;
        RECT 2027.950 145.030 2043.010 145.330 ;
        RECT 2124.590 145.330 2124.890 145.710 ;
        RECT 2139.310 145.710 2186.315 146.010 ;
        RECT 2139.310 145.330 2139.610 145.710 ;
        RECT 2185.985 145.695 2186.315 145.710 ;
        RECT 2187.365 146.010 2187.695 146.025 ;
        RECT 2187.365 145.710 2221.490 146.010 ;
        RECT 2187.365 145.695 2187.695 145.710 ;
        RECT 2124.590 145.030 2139.610 145.330 ;
        RECT 2221.190 145.330 2221.490 145.710 ;
        RECT 2235.910 145.330 2236.210 146.390 ;
        RECT 2317.790 146.010 2318.090 146.390 ;
        RECT 2339.625 146.390 2380.435 146.690 ;
        RECT 2339.625 146.375 2339.955 146.390 ;
        RECT 2380.105 146.375 2380.435 146.390 ;
        RECT 2511.205 146.690 2511.535 146.705 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2511.205 146.390 2546.250 146.690 ;
        RECT 2511.205 146.375 2511.535 146.390 ;
        RECT 2326.285 146.010 2326.615 146.025 ;
        RECT 2317.790 145.710 2326.615 146.010 ;
        RECT 2326.285 145.695 2326.615 145.710 ;
        RECT 2381.025 146.010 2381.355 146.025 ;
        RECT 2407.910 146.010 2408.290 146.020 ;
        RECT 2381.025 145.710 2408.290 146.010 ;
        RECT 2545.950 146.010 2546.250 146.390 ;
        RECT 2594.710 146.390 2642.850 146.690 ;
        RECT 2545.950 145.710 2594.090 146.010 ;
        RECT 2381.025 145.695 2381.355 145.710 ;
        RECT 2407.910 145.700 2408.290 145.710 ;
        RECT 2221.190 145.030 2236.210 145.330 ;
        RECT 2456.005 145.330 2456.335 145.345 ;
        RECT 2463.825 145.330 2464.155 145.345 ;
        RECT 2456.005 145.030 2464.155 145.330 ;
        RECT 2593.790 145.330 2594.090 145.710 ;
        RECT 2594.710 145.330 2595.010 146.390 ;
        RECT 2642.550 146.010 2642.850 146.390 ;
        RECT 2691.310 146.390 2739.450 146.690 ;
        RECT 2642.550 145.710 2690.690 146.010 ;
        RECT 2593.790 145.030 2595.010 145.330 ;
        RECT 2690.390 145.330 2690.690 145.710 ;
        RECT 2691.310 145.330 2691.610 146.390 ;
        RECT 2739.150 146.010 2739.450 146.390 ;
        RECT 2787.910 146.390 2836.050 146.690 ;
        RECT 2739.150 145.710 2787.290 146.010 ;
        RECT 2690.390 145.030 2691.610 145.330 ;
        RECT 2786.990 145.330 2787.290 145.710 ;
        RECT 2787.910 145.330 2788.210 146.390 ;
        RECT 2835.750 146.010 2836.050 146.390 ;
        RECT 2916.710 146.390 2924.800 146.690 ;
        RECT 2916.710 146.010 2917.010 146.390 ;
        RECT 2835.750 145.710 2883.890 146.010 ;
        RECT 2786.990 145.030 2788.210 145.330 ;
        RECT 2883.590 145.330 2883.890 145.710 ;
        RECT 2884.510 145.710 2917.010 146.010 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
        RECT 2884.510 145.330 2884.810 145.710 ;
        RECT 2883.590 145.030 2884.810 145.330 ;
        RECT 1635.110 145.020 1635.490 145.030 ;
        RECT 1683.205 145.015 1683.535 145.030 ;
        RECT 1835.465 145.015 1835.795 145.030 ;
        RECT 2027.950 145.020 2028.330 145.030 ;
        RECT 2456.005 145.015 2456.335 145.030 ;
        RECT 2463.825 145.015 2464.155 145.030 ;
        RECT 1436.390 144.650 1436.770 144.660 ;
        RECT 1531.405 144.650 1531.735 144.665 ;
        RECT 1436.390 144.350 1531.735 144.650 ;
        RECT 1436.390 144.340 1436.770 144.350 ;
        RECT 1531.405 144.335 1531.735 144.350 ;
        RECT 1572.805 144.650 1573.135 144.665 ;
        RECT 1579.950 144.650 1581.170 144.820 ;
        RECT 1572.805 144.520 1581.170 144.650 ;
        RECT 1628.005 144.650 1628.335 144.665 ;
        RECT 1634.905 144.650 1635.235 144.665 ;
        RECT 1572.805 144.350 1580.250 144.520 ;
        RECT 1628.005 144.350 1635.235 144.650 ;
        RECT 1572.805 144.335 1573.135 144.350 ;
        RECT 1628.005 144.335 1628.335 144.350 ;
        RECT 1634.905 144.335 1635.235 144.350 ;
      LAYER via3 ;
        RECT 1178.820 2896.300 1179.140 2896.620 ;
        RECT 1178.820 146.380 1179.140 146.700 ;
        RECT 1635.140 146.380 1635.460 146.700 ;
        RECT 1435.500 145.700 1435.820 146.020 ;
        RECT 1635.140 145.020 1635.460 145.340 ;
        RECT 2027.980 147.060 2028.300 147.380 ;
        RECT 2407.940 147.060 2408.260 147.380 ;
        RECT 2027.980 145.020 2028.300 145.340 ;
        RECT 2407.940 145.700 2408.260 146.020 ;
        RECT 1436.420 144.340 1436.740 144.660 ;
      LAYER met4 ;
        RECT 1178.815 2896.295 1179.145 2896.625 ;
        RECT 1178.830 146.705 1179.130 2896.295 ;
        RECT 1435.510 147.750 1436.730 148.050 ;
        RECT 1178.815 146.375 1179.145 146.705 ;
        RECT 1435.510 146.025 1435.810 147.750 ;
        RECT 1435.495 145.695 1435.825 146.025 ;
        RECT 1436.430 144.665 1436.730 147.750 ;
        RECT 2027.975 147.055 2028.305 147.385 ;
        RECT 2407.935 147.055 2408.265 147.385 ;
        RECT 1635.135 146.375 1635.465 146.705 ;
        RECT 1635.150 145.345 1635.450 146.375 ;
        RECT 2027.990 145.345 2028.290 147.055 ;
        RECT 2407.950 146.025 2408.250 147.055 ;
        RECT 2407.935 145.695 2408.265 146.025 ;
        RECT 1635.135 145.015 1635.465 145.345 ;
        RECT 2027.975 145.015 2028.305 145.345 ;
        RECT 1436.415 144.335 1436.745 144.665 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1490.930 2918.120 1491.250 2918.180 ;
        RECT 2348.830 2918.120 2349.150 2918.180 ;
        RECT 1490.930 2917.980 2349.150 2918.120 ;
        RECT 1490.930 2917.920 1491.250 2917.980 ;
        RECT 2348.830 2917.920 2349.150 2917.980 ;
        RECT 2348.830 2497.540 2349.150 2497.600 ;
        RECT 2898.990 2497.540 2899.310 2497.600 ;
        RECT 2348.830 2497.400 2899.310 2497.540 ;
        RECT 2348.830 2497.340 2349.150 2497.400 ;
        RECT 2898.990 2497.340 2899.310 2497.400 ;
      LAYER via ;
        RECT 1490.960 2917.920 1491.220 2918.180 ;
        RECT 2348.860 2917.920 2349.120 2918.180 ;
        RECT 2348.860 2497.340 2349.120 2497.600 ;
        RECT 2899.020 2497.340 2899.280 2497.600 ;
      LAYER met2 ;
        RECT 1490.960 2917.890 1491.220 2918.210 ;
        RECT 2348.860 2917.890 2349.120 2918.210 ;
        RECT 1491.020 2900.000 1491.160 2917.890 ;
        RECT 1490.885 2896.000 1491.165 2900.000 ;
        RECT 2348.920 2497.630 2349.060 2917.890 ;
        RECT 2348.860 2497.310 2349.120 2497.630 ;
        RECT 2899.020 2497.310 2899.280 2497.630 ;
        RECT 2899.080 2493.405 2899.220 2497.310 ;
        RECT 2899.010 2493.035 2899.290 2493.405 ;
      LAYER via2 ;
        RECT 2899.010 2493.080 2899.290 2493.360 ;
      LAYER met3 ;
        RECT 2898.985 2493.370 2899.315 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2898.985 2493.070 2924.800 2493.370 ;
        RECT 2898.985 2493.055 2899.315 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1522.670 2918.460 1522.990 2918.520 ;
        RECT 2356.190 2918.460 2356.510 2918.520 ;
        RECT 1522.670 2918.320 2356.510 2918.460 ;
        RECT 1522.670 2918.260 1522.990 2918.320 ;
        RECT 2356.190 2918.260 2356.510 2918.320 ;
        RECT 2356.190 2732.140 2356.510 2732.200 ;
        RECT 2898.990 2732.140 2899.310 2732.200 ;
        RECT 2356.190 2732.000 2899.310 2732.140 ;
        RECT 2356.190 2731.940 2356.510 2732.000 ;
        RECT 2898.990 2731.940 2899.310 2732.000 ;
      LAYER via ;
        RECT 1522.700 2918.260 1522.960 2918.520 ;
        RECT 2356.220 2918.260 2356.480 2918.520 ;
        RECT 2356.220 2731.940 2356.480 2732.200 ;
        RECT 2899.020 2731.940 2899.280 2732.200 ;
      LAYER met2 ;
        RECT 1522.700 2918.230 1522.960 2918.550 ;
        RECT 2356.220 2918.230 2356.480 2918.550 ;
        RECT 1522.760 2900.000 1522.900 2918.230 ;
        RECT 1522.625 2896.000 1522.905 2900.000 ;
        RECT 2356.280 2732.230 2356.420 2918.230 ;
        RECT 2356.220 2731.910 2356.480 2732.230 ;
        RECT 2899.020 2731.910 2899.280 2732.230 ;
        RECT 2899.080 2728.005 2899.220 2731.910 ;
        RECT 2899.010 2727.635 2899.290 2728.005 ;
      LAYER via2 ;
        RECT 2899.010 2727.680 2899.290 2727.960 ;
      LAYER met3 ;
        RECT 2898.985 2727.970 2899.315 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2898.985 2727.670 2924.800 2727.970 ;
        RECT 2898.985 2727.655 2899.315 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1559.010 2960.280 1559.330 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 1559.010 2960.140 2901.150 2960.280 ;
        RECT 1559.010 2960.080 1559.330 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
      LAYER via ;
        RECT 1559.040 2960.080 1559.300 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 1559.040 2960.050 1559.300 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 1559.100 2900.610 1559.240 2960.050 ;
        RECT 1556.340 2900.470 1559.240 2900.610 ;
        RECT 1553.905 2899.250 1554.185 2900.000 ;
        RECT 1556.340 2899.250 1556.480 2900.470 ;
        RECT 1553.905 2899.110 1556.480 2899.250 ;
        RECT 1553.905 2896.000 1554.185 2899.110 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1586.610 3194.880 1586.930 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 1586.610 3194.740 2901.150 3194.880 ;
        RECT 1586.610 3194.680 1586.930 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 1586.640 3194.680 1586.900 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 1586.640 3194.650 1586.900 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 1585.645 2899.930 1585.925 2900.000 ;
        RECT 1586.700 2899.930 1586.840 3194.650 ;
        RECT 1585.645 2899.790 1586.840 2899.930 ;
        RECT 1585.645 2896.000 1585.925 2899.790 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2146.060 3429.680 2149.880 3429.820 ;
        RECT 1621.110 3429.480 1621.430 3429.540 ;
        RECT 2146.060 3429.480 2146.200 3429.680 ;
        RECT 1621.110 3429.340 2146.200 3429.480 ;
        RECT 2149.740 3429.480 2149.880 3429.680 ;
        RECT 2762.920 3429.680 2798.940 3429.820 ;
        RECT 2762.920 3429.480 2763.060 3429.680 ;
        RECT 2149.740 3429.340 2763.060 3429.480 ;
        RECT 2798.800 3429.480 2798.940 3429.680 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 2798.800 3429.340 2901.150 3429.480 ;
        RECT 1621.110 3429.280 1621.430 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 1621.140 3429.280 1621.400 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1621.140 3429.250 1621.400 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1616.925 2899.250 1617.205 2900.000 ;
        RECT 1621.200 2899.250 1621.340 3429.250 ;
        RECT 1616.925 2899.110 1621.340 2899.250 ;
        RECT 1616.925 2896.000 1617.205 2899.110 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1648.710 3503.940 1649.030 3504.000 ;
        RECT 2717.290 3503.940 2717.610 3504.000 ;
        RECT 1648.710 3503.800 2717.610 3503.940 ;
        RECT 1648.710 3503.740 1649.030 3503.800 ;
        RECT 2717.290 3503.740 2717.610 3503.800 ;
      LAYER via ;
        RECT 1648.740 3503.740 1649.000 3504.000 ;
        RECT 2717.320 3503.740 2717.580 3504.000 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3504.030 2717.520 3517.600 ;
        RECT 1648.740 3503.710 1649.000 3504.030 ;
        RECT 2717.320 3503.710 2717.580 3504.030 ;
        RECT 1648.800 2900.000 1648.940 3503.710 ;
        RECT 1648.665 2896.000 1648.945 2900.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1683.210 3500.880 1683.530 3500.940 ;
        RECT 2392.530 3500.880 2392.850 3500.940 ;
        RECT 1683.210 3500.740 2392.850 3500.880 ;
        RECT 1683.210 3500.680 1683.530 3500.740 ;
        RECT 2392.530 3500.680 2392.850 3500.740 ;
      LAYER via ;
        RECT 1683.240 3500.680 1683.500 3500.940 ;
        RECT 2392.560 3500.680 2392.820 3500.940 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3500.970 2392.760 3517.600 ;
        RECT 1683.240 3500.650 1683.500 3500.970 ;
        RECT 2392.560 3500.650 2392.820 3500.970 ;
        RECT 1680.405 2899.250 1680.685 2900.000 ;
        RECT 1683.300 2899.250 1683.440 3500.650 ;
        RECT 1680.405 2899.110 1683.440 2899.250 ;
        RECT 1680.405 2896.000 1680.685 2899.110 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1717.710 3499.180 1718.030 3499.240 ;
        RECT 2068.230 3499.180 2068.550 3499.240 ;
        RECT 1717.710 3499.040 2068.550 3499.180 ;
        RECT 1717.710 3498.980 1718.030 3499.040 ;
        RECT 2068.230 3498.980 2068.550 3499.040 ;
      LAYER via ;
        RECT 1717.740 3498.980 1718.000 3499.240 ;
        RECT 2068.260 3498.980 2068.520 3499.240 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3499.270 2068.460 3517.600 ;
        RECT 1717.740 3498.950 1718.000 3499.270 ;
        RECT 2068.260 3498.950 2068.520 3499.270 ;
        RECT 1711.685 2899.250 1711.965 2900.000 ;
        RECT 1717.800 2899.250 1717.940 3498.950 ;
        RECT 1711.685 2899.110 1717.940 2899.250 ;
        RECT 1711.685 2896.000 1711.965 2899.110 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1738.870 3498.500 1739.190 3498.560 ;
        RECT 1743.930 3498.500 1744.250 3498.560 ;
        RECT 1738.870 3498.360 1744.250 3498.500 ;
        RECT 1738.870 3498.300 1739.190 3498.360 ;
        RECT 1743.930 3498.300 1744.250 3498.360 ;
      LAYER via ;
        RECT 1738.900 3498.300 1739.160 3498.560 ;
        RECT 1743.960 3498.300 1744.220 3498.560 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3498.590 1744.160 3517.600 ;
        RECT 1738.900 3498.270 1739.160 3498.590 ;
        RECT 1743.960 3498.270 1744.220 3498.590 ;
        RECT 1738.960 2899.250 1739.100 3498.270 ;
        RECT 1743.425 2899.250 1743.705 2900.000 ;
        RECT 1738.960 2899.110 1743.705 2899.250 ;
        RECT 1743.425 2896.000 1743.705 2899.110 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.170 3499.520 1419.490 3499.580 ;
        RECT 1773.370 3499.520 1773.690 3499.580 ;
        RECT 1419.170 3499.380 1773.690 3499.520 ;
        RECT 1419.170 3499.320 1419.490 3499.380 ;
        RECT 1773.370 3499.320 1773.690 3499.380 ;
      LAYER via ;
        RECT 1419.200 3499.320 1419.460 3499.580 ;
        RECT 1773.400 3499.320 1773.660 3499.580 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3499.610 1419.400 3517.600 ;
        RECT 1419.200 3499.290 1419.460 3499.610 ;
        RECT 1773.400 3499.290 1773.660 3499.610 ;
        RECT 1773.460 2899.930 1773.600 3499.290 ;
        RECT 1775.165 2899.930 1775.445 2900.000 ;
        RECT 1773.460 2899.790 1775.445 2899.930 ;
        RECT 1775.165 2896.000 1775.445 2899.790 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1891.130 381.380 1891.450 381.440 ;
        RECT 1931.610 381.380 1931.930 381.440 ;
        RECT 1891.130 381.240 1931.930 381.380 ;
        RECT 1891.130 381.180 1891.450 381.240 ;
        RECT 1931.610 381.180 1931.930 381.240 ;
        RECT 2173.570 380.700 2173.890 380.760 ;
        RECT 2187.370 380.700 2187.690 380.760 ;
        RECT 2173.570 380.560 2187.690 380.700 ;
        RECT 2173.570 380.500 2173.890 380.560 ;
        RECT 2187.370 380.500 2187.690 380.560 ;
        RECT 2318.470 380.700 2318.790 380.760 ;
        RECT 2339.630 380.700 2339.950 380.760 ;
        RECT 2318.470 380.560 2339.950 380.700 ;
        RECT 2318.470 380.500 2318.790 380.560 ;
        RECT 2339.630 380.500 2339.950 380.560 ;
        RECT 2089.390 380.360 2089.710 380.420 ;
        RECT 2096.750 380.360 2097.070 380.420 ;
        RECT 2089.390 380.220 2097.070 380.360 ;
        RECT 2089.390 380.160 2089.710 380.220 ;
        RECT 2096.750 380.160 2097.070 380.220 ;
        RECT 1352.470 380.020 1352.790 380.080 ;
        RECT 1376.850 380.020 1377.170 380.080 ;
        RECT 1352.470 379.880 1377.170 380.020 ;
        RECT 1352.470 379.820 1352.790 379.880 ;
        RECT 1376.850 379.820 1377.170 379.880 ;
      LAYER via ;
        RECT 1891.160 381.180 1891.420 381.440 ;
        RECT 1931.640 381.180 1931.900 381.440 ;
        RECT 2173.600 380.500 2173.860 380.760 ;
        RECT 2187.400 380.500 2187.660 380.760 ;
        RECT 2318.500 380.500 2318.760 380.760 ;
        RECT 2339.660 380.500 2339.920 380.760 ;
        RECT 2089.420 380.160 2089.680 380.420 ;
        RECT 2096.780 380.160 2097.040 380.420 ;
        RECT 1352.500 379.820 1352.760 380.080 ;
        RECT 1376.880 379.820 1377.140 380.080 ;
      LAYER met2 ;
        RECT 1206.605 2896.530 1206.885 2900.000 ;
        RECT 1207.130 2896.530 1207.410 2896.645 ;
        RECT 1206.605 2896.390 1207.410 2896.530 ;
        RECT 1206.605 2896.000 1206.885 2896.390 ;
        RECT 1207.130 2896.275 1207.410 2896.390 ;
        RECT 2414.630 382.315 2414.910 382.685 ;
        RECT 1891.160 381.325 1891.420 381.470 ;
        RECT 1931.640 381.325 1931.900 381.470 ;
        RECT 1891.150 380.955 1891.430 381.325 ;
        RECT 1931.630 380.955 1931.910 381.325 ;
        RECT 2339.650 380.955 2339.930 381.325 ;
        RECT 2339.720 380.790 2339.860 380.955 ;
        RECT 2173.600 380.645 2173.860 380.790 ;
        RECT 2187.400 380.645 2187.660 380.790 ;
        RECT 2318.500 380.645 2318.760 380.790 ;
        RECT 1255.890 380.275 1256.170 380.645 ;
        RECT 1376.870 380.275 1377.150 380.645 ;
        RECT 1423.330 380.530 1423.610 380.645 ;
        RECT 1800.530 380.530 1800.810 380.645 ;
        RECT 1801.450 380.530 1801.730 380.645 ;
        RECT 1423.330 380.390 1424.000 380.530 ;
        RECT 1423.330 380.275 1423.610 380.390 ;
        RECT 1255.960 378.605 1256.100 380.275 ;
        RECT 1376.940 380.110 1377.080 380.275 ;
        RECT 1352.500 379.965 1352.760 380.110 ;
        RECT 1352.490 379.595 1352.770 379.965 ;
        RECT 1376.880 379.790 1377.140 380.110 ;
        RECT 1423.860 379.965 1424.000 380.390 ;
        RECT 1800.530 380.390 1801.730 380.530 ;
        RECT 1800.530 380.275 1800.810 380.390 ;
        RECT 1801.450 380.275 1801.730 380.390 ;
        RECT 2089.410 380.275 2089.690 380.645 ;
        RECT 2096.770 380.275 2097.050 380.645 ;
        RECT 2173.590 380.275 2173.870 380.645 ;
        RECT 2187.390 380.275 2187.670 380.645 ;
        RECT 2318.490 380.275 2318.770 380.645 ;
        RECT 2339.660 380.470 2339.920 380.790 ;
        RECT 2414.700 380.645 2414.840 382.315 ;
        RECT 2439.010 381.635 2439.290 382.005 ;
        RECT 2414.630 380.275 2414.910 380.645 ;
        RECT 2089.420 380.130 2089.680 380.275 ;
        RECT 2096.780 380.130 2097.040 380.275 ;
        RECT 2439.080 379.965 2439.220 381.635 ;
        RECT 1423.790 379.595 1424.070 379.965 ;
        RECT 2439.010 379.595 2439.290 379.965 ;
        RECT 1255.890 378.235 1256.170 378.605 ;
      LAYER via2 ;
        RECT 1207.130 2896.320 1207.410 2896.600 ;
        RECT 2414.630 382.360 2414.910 382.640 ;
        RECT 1891.150 381.000 1891.430 381.280 ;
        RECT 1931.630 381.000 1931.910 381.280 ;
        RECT 2339.650 381.000 2339.930 381.280 ;
        RECT 1255.890 380.320 1256.170 380.600 ;
        RECT 1376.870 380.320 1377.150 380.600 ;
        RECT 1423.330 380.320 1423.610 380.600 ;
        RECT 1352.490 379.640 1352.770 379.920 ;
        RECT 1800.530 380.320 1800.810 380.600 ;
        RECT 1801.450 380.320 1801.730 380.600 ;
        RECT 2089.410 380.320 2089.690 380.600 ;
        RECT 2096.770 380.320 2097.050 380.600 ;
        RECT 2173.590 380.320 2173.870 380.600 ;
        RECT 2187.390 380.320 2187.670 380.600 ;
        RECT 2318.490 380.320 2318.770 380.600 ;
        RECT 2439.010 381.680 2439.290 381.960 ;
        RECT 2414.630 380.320 2414.910 380.600 ;
        RECT 1423.790 379.640 1424.070 379.920 ;
        RECT 2439.010 379.640 2439.290 379.920 ;
        RECT 1255.890 378.280 1256.170 378.560 ;
      LAYER met3 ;
        RECT 1206.390 2896.610 1206.770 2896.620 ;
        RECT 1207.105 2896.610 1207.435 2896.625 ;
        RECT 1206.390 2896.310 1207.435 2896.610 ;
        RECT 1206.390 2896.300 1206.770 2896.310 ;
        RECT 1207.105 2896.295 1207.435 2896.310 ;
        RECT 2366.510 382.650 2366.890 382.660 ;
        RECT 2414.605 382.650 2414.935 382.665 ;
        RECT 2366.510 382.350 2414.935 382.650 ;
        RECT 2366.510 382.340 2366.890 382.350 ;
        RECT 2414.605 382.335 2414.935 382.350 ;
        RECT 2438.985 381.970 2439.315 381.985 ;
        RECT 1993.030 381.670 2028.290 381.970 ;
        RECT 1497.110 381.290 1497.490 381.300 ;
        RECT 1538.510 381.290 1538.890 381.300 ;
        RECT 1891.125 381.290 1891.455 381.305 ;
        RECT 1497.110 380.990 1538.890 381.290 ;
        RECT 1497.110 380.980 1497.490 380.990 ;
        RECT 1538.510 380.980 1538.890 380.990 ;
        RECT 1655.390 380.990 1704.450 381.290 ;
        RECT 1206.390 380.610 1206.770 380.620 ;
        RECT 1255.865 380.610 1256.195 380.625 ;
        RECT 1206.390 380.310 1256.195 380.610 ;
        RECT 1206.390 380.300 1206.770 380.310 ;
        RECT 1255.865 380.295 1256.195 380.310 ;
        RECT 1376.845 380.610 1377.175 380.625 ;
        RECT 1423.305 380.610 1423.635 380.625 ;
        RECT 1376.845 380.310 1423.635 380.610 ;
        RECT 1376.845 380.295 1377.175 380.310 ;
        RECT 1423.305 380.295 1423.635 380.310 ;
        RECT 1303.910 379.930 1304.290 379.940 ;
        RECT 1352.465 379.930 1352.795 379.945 ;
        RECT 1303.910 379.630 1352.795 379.930 ;
        RECT 1303.910 379.620 1304.290 379.630 ;
        RECT 1352.465 379.615 1352.795 379.630 ;
        RECT 1423.765 379.930 1424.095 379.945 ;
        RECT 1497.110 379.930 1497.490 379.940 ;
        RECT 1423.765 379.630 1424.770 379.930 ;
        RECT 1423.765 379.615 1424.095 379.630 ;
        RECT 1255.865 378.570 1256.195 378.585 ;
        RECT 1303.910 378.570 1304.290 378.580 ;
        RECT 1255.865 378.270 1304.290 378.570 ;
        RECT 1424.470 378.570 1424.770 379.630 ;
        RECT 1441.030 379.630 1497.490 379.930 ;
        RECT 1441.030 378.570 1441.330 379.630 ;
        RECT 1497.110 379.620 1497.490 379.630 ;
        RECT 1538.510 379.930 1538.890 379.940 ;
        RECT 1655.390 379.930 1655.690 380.990 ;
        RECT 1538.510 379.630 1655.690 379.930 ;
        RECT 1704.150 379.930 1704.450 380.990 ;
        RECT 1849.510 380.990 1891.455 381.290 ;
        RECT 1800.505 380.610 1800.835 380.625 ;
        RECT 1752.910 380.310 1800.835 380.610 ;
        RECT 1752.910 379.930 1753.210 380.310 ;
        RECT 1800.505 380.295 1800.835 380.310 ;
        RECT 1801.425 380.610 1801.755 380.625 ;
        RECT 1801.425 380.310 1848.890 380.610 ;
        RECT 1801.425 380.295 1801.755 380.310 ;
        RECT 1704.150 379.630 1753.210 379.930 ;
        RECT 1848.590 379.930 1848.890 380.310 ;
        RECT 1849.510 379.930 1849.810 380.990 ;
        RECT 1891.125 380.975 1891.455 380.990 ;
        RECT 1931.605 381.290 1931.935 381.305 ;
        RECT 1931.605 380.990 1945.490 381.290 ;
        RECT 1931.605 380.975 1931.935 380.990 ;
        RECT 1848.590 379.630 1849.810 379.930 ;
        RECT 1945.190 379.930 1945.490 380.990 ;
        RECT 1993.030 380.610 1993.330 381.670 ;
        RECT 1946.110 380.310 1993.330 380.610 ;
        RECT 1946.110 379.930 1946.410 380.310 ;
        RECT 1945.190 379.630 1946.410 379.930 ;
        RECT 2027.990 379.930 2028.290 381.670 ;
        RECT 2415.310 381.670 2439.315 381.970 ;
        RECT 2339.625 381.290 2339.955 381.305 ;
        RECT 2366.510 381.290 2366.890 381.300 ;
        RECT 2235.910 380.990 2283.130 381.290 ;
        RECT 2089.385 380.610 2089.715 380.625 ;
        RECT 2042.710 380.310 2089.715 380.610 ;
        RECT 2042.710 379.930 2043.010 380.310 ;
        RECT 2089.385 380.295 2089.715 380.310 ;
        RECT 2096.745 380.610 2097.075 380.625 ;
        RECT 2173.565 380.610 2173.895 380.625 ;
        RECT 2096.745 380.310 2124.890 380.610 ;
        RECT 2096.745 380.295 2097.075 380.310 ;
        RECT 2027.990 379.630 2043.010 379.930 ;
        RECT 2124.590 379.930 2124.890 380.310 ;
        RECT 2139.310 380.310 2173.895 380.610 ;
        RECT 2139.310 379.930 2139.610 380.310 ;
        RECT 2173.565 380.295 2173.895 380.310 ;
        RECT 2187.365 380.610 2187.695 380.625 ;
        RECT 2187.365 380.310 2221.490 380.610 ;
        RECT 2187.365 380.295 2187.695 380.310 ;
        RECT 2124.590 379.630 2139.610 379.930 ;
        RECT 2221.190 379.930 2221.490 380.310 ;
        RECT 2235.910 379.930 2236.210 380.990 ;
        RECT 2282.830 380.610 2283.130 380.990 ;
        RECT 2339.625 380.990 2366.890 381.290 ;
        RECT 2339.625 380.975 2339.955 380.990 ;
        RECT 2366.510 380.980 2366.890 380.990 ;
        RECT 2318.465 380.610 2318.795 380.625 ;
        RECT 2282.830 380.310 2318.795 380.610 ;
        RECT 2318.465 380.295 2318.795 380.310 ;
        RECT 2414.605 380.610 2414.935 380.625 ;
        RECT 2415.310 380.610 2415.610 381.670 ;
        RECT 2438.985 381.655 2439.315 381.670 ;
        RECT 2463.110 381.290 2463.490 381.300 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 2463.110 380.990 2546.250 381.290 ;
        RECT 2463.110 380.980 2463.490 380.990 ;
        RECT 2414.605 380.310 2415.610 380.610 ;
        RECT 2545.950 380.610 2546.250 380.990 ;
        RECT 2594.710 380.990 2642.850 381.290 ;
        RECT 2545.950 380.310 2594.090 380.610 ;
        RECT 2414.605 380.295 2414.935 380.310 ;
        RECT 2221.190 379.630 2236.210 379.930 ;
        RECT 2438.985 379.930 2439.315 379.945 ;
        RECT 2463.110 379.930 2463.490 379.940 ;
        RECT 2438.985 379.630 2463.490 379.930 ;
        RECT 2593.790 379.930 2594.090 380.310 ;
        RECT 2594.710 379.930 2595.010 380.990 ;
        RECT 2642.550 380.610 2642.850 380.990 ;
        RECT 2691.310 380.990 2739.450 381.290 ;
        RECT 2642.550 380.310 2690.690 380.610 ;
        RECT 2593.790 379.630 2595.010 379.930 ;
        RECT 2690.390 379.930 2690.690 380.310 ;
        RECT 2691.310 379.930 2691.610 380.990 ;
        RECT 2739.150 380.610 2739.450 380.990 ;
        RECT 2787.910 380.990 2836.050 381.290 ;
        RECT 2739.150 380.310 2787.290 380.610 ;
        RECT 2690.390 379.630 2691.610 379.930 ;
        RECT 2786.990 379.930 2787.290 380.310 ;
        RECT 2787.910 379.930 2788.210 380.990 ;
        RECT 2835.750 380.610 2836.050 380.990 ;
        RECT 2916.710 380.990 2924.800 381.290 ;
        RECT 2916.710 380.610 2917.010 380.990 ;
        RECT 2835.750 380.310 2883.890 380.610 ;
        RECT 2786.990 379.630 2788.210 379.930 ;
        RECT 2883.590 379.930 2883.890 380.310 ;
        RECT 2884.510 380.310 2917.010 380.610 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
        RECT 2884.510 379.930 2884.810 380.310 ;
        RECT 2883.590 379.630 2884.810 379.930 ;
        RECT 1538.510 379.620 1538.890 379.630 ;
        RECT 2438.985 379.615 2439.315 379.630 ;
        RECT 2463.110 379.620 2463.490 379.630 ;
        RECT 1424.470 378.270 1441.330 378.570 ;
        RECT 1255.865 378.255 1256.195 378.270 ;
        RECT 1303.910 378.260 1304.290 378.270 ;
      LAYER via3 ;
        RECT 1206.420 2896.300 1206.740 2896.620 ;
        RECT 2366.540 382.340 2366.860 382.660 ;
        RECT 1497.140 380.980 1497.460 381.300 ;
        RECT 1538.540 380.980 1538.860 381.300 ;
        RECT 1206.420 380.300 1206.740 380.620 ;
        RECT 1303.940 379.620 1304.260 379.940 ;
        RECT 1303.940 378.260 1304.260 378.580 ;
        RECT 1497.140 379.620 1497.460 379.940 ;
        RECT 1538.540 379.620 1538.860 379.940 ;
        RECT 2366.540 380.980 2366.860 381.300 ;
        RECT 2463.140 380.980 2463.460 381.300 ;
        RECT 2463.140 379.620 2463.460 379.940 ;
      LAYER met4 ;
        RECT 1206.415 2896.295 1206.745 2896.625 ;
        RECT 1206.430 380.625 1206.730 2896.295 ;
        RECT 2366.535 382.335 2366.865 382.665 ;
        RECT 2366.550 381.305 2366.850 382.335 ;
        RECT 1497.135 380.975 1497.465 381.305 ;
        RECT 1538.535 380.975 1538.865 381.305 ;
        RECT 2366.535 380.975 2366.865 381.305 ;
        RECT 2463.135 380.975 2463.465 381.305 ;
        RECT 1206.415 380.295 1206.745 380.625 ;
        RECT 1497.150 379.945 1497.450 380.975 ;
        RECT 1538.550 379.945 1538.850 380.975 ;
        RECT 2463.150 379.945 2463.450 380.975 ;
        RECT 1303.935 379.615 1304.265 379.945 ;
        RECT 1497.135 379.615 1497.465 379.945 ;
        RECT 1538.535 379.615 1538.865 379.945 ;
        RECT 2463.135 379.615 2463.465 379.945 ;
        RECT 1303.950 378.585 1304.250 379.615 ;
        RECT 1303.935 378.255 1304.265 378.585 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1094.870 3501.220 1095.190 3501.280 ;
        RECT 1800.970 3501.220 1801.290 3501.280 ;
        RECT 1094.870 3501.080 1801.290 3501.220 ;
        RECT 1094.870 3501.020 1095.190 3501.080 ;
        RECT 1800.970 3501.020 1801.290 3501.080 ;
      LAYER via ;
        RECT 1094.900 3501.020 1095.160 3501.280 ;
        RECT 1801.000 3501.020 1801.260 3501.280 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3501.310 1095.100 3517.600 ;
        RECT 1094.900 3500.990 1095.160 3501.310 ;
        RECT 1801.000 3500.990 1801.260 3501.310 ;
        RECT 1801.060 2900.610 1801.200 3500.990 ;
        RECT 1801.060 2900.470 1804.420 2900.610 ;
        RECT 1804.280 2899.250 1804.420 2900.470 ;
        RECT 1806.445 2899.250 1806.725 2900.000 ;
        RECT 1804.280 2899.110 1806.725 2899.250 ;
        RECT 1806.445 2896.000 1806.725 2899.110 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 770.570 3503.600 770.890 3503.660 ;
        RECT 1835.470 3503.600 1835.790 3503.660 ;
        RECT 770.570 3503.460 1835.790 3503.600 ;
        RECT 770.570 3503.400 770.890 3503.460 ;
        RECT 1835.470 3503.400 1835.790 3503.460 ;
      LAYER via ;
        RECT 770.600 3503.400 770.860 3503.660 ;
        RECT 1835.500 3503.400 1835.760 3503.660 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3503.690 770.800 3517.600 ;
        RECT 770.600 3503.370 770.860 3503.690 ;
        RECT 1835.500 3503.370 1835.760 3503.690 ;
        RECT 1835.560 2899.250 1835.700 3503.370 ;
        RECT 1838.185 2899.250 1838.465 2900.000 ;
        RECT 1835.560 2899.110 1838.465 2899.250 ;
        RECT 1838.185 2896.000 1838.465 2899.110 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3502.580 446.130 3502.640 ;
        RECT 1869.970 3502.580 1870.290 3502.640 ;
        RECT 445.810 3502.440 1870.290 3502.580 ;
        RECT 445.810 3502.380 446.130 3502.440 ;
        RECT 1869.970 3502.380 1870.290 3502.440 ;
      LAYER via ;
        RECT 445.840 3502.380 446.100 3502.640 ;
        RECT 1870.000 3502.380 1870.260 3502.640 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3502.670 446.040 3517.600 ;
        RECT 445.840 3502.350 446.100 3502.670 ;
        RECT 1870.000 3502.350 1870.260 3502.670 ;
        RECT 1870.060 2900.000 1870.200 3502.350 ;
        RECT 1869.925 2896.000 1870.205 2900.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 121.510 3501.560 121.830 3501.620 ;
        RECT 1897.570 3501.560 1897.890 3501.620 ;
        RECT 121.510 3501.420 1897.890 3501.560 ;
        RECT 121.510 3501.360 121.830 3501.420 ;
        RECT 1897.570 3501.360 1897.890 3501.420 ;
      LAYER via ;
        RECT 121.540 3501.360 121.800 3501.620 ;
        RECT 1897.600 3501.360 1897.860 3501.620 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3501.650 121.740 3517.600 ;
        RECT 121.540 3501.330 121.800 3501.650 ;
        RECT 1897.600 3501.330 1897.860 3501.650 ;
        RECT 1897.660 2899.250 1897.800 3501.330 ;
        RECT 1901.205 2899.250 1901.485 2900.000 ;
        RECT 1897.660 2899.110 1901.485 2899.250 ;
        RECT 1901.205 2896.000 1901.485 2899.110 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3339.720 17.410 3339.780 ;
        RECT 1932.070 3339.720 1932.390 3339.780 ;
        RECT 17.090 3339.580 1932.390 3339.720 ;
        RECT 17.090 3339.520 17.410 3339.580 ;
        RECT 1932.070 3339.520 1932.390 3339.580 ;
      LAYER via ;
        RECT 17.120 3339.520 17.380 3339.780 ;
        RECT 1932.100 3339.520 1932.360 3339.780 ;
      LAYER met2 ;
        RECT 17.110 3339.635 17.390 3340.005 ;
        RECT 17.120 3339.490 17.380 3339.635 ;
        RECT 1932.100 3339.490 1932.360 3339.810 ;
        RECT 1932.160 2899.930 1932.300 3339.490 ;
        RECT 1932.945 2899.930 1933.225 2900.000 ;
        RECT 1932.160 2899.790 1933.225 2899.930 ;
        RECT 1932.945 2896.000 1933.225 2899.790 ;
      LAYER via2 ;
        RECT 17.110 3339.680 17.390 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.085 3339.970 17.415 3339.985 ;
        RECT -4.800 3339.670 17.415 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.085 3339.655 17.415 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.090 3050.040 17.410 3050.100 ;
        RECT 1959.670 3050.040 1959.990 3050.100 ;
        RECT 17.090 3049.900 1959.990 3050.040 ;
        RECT 17.090 3049.840 17.410 3049.900 ;
        RECT 1959.670 3049.840 1959.990 3049.900 ;
      LAYER via ;
        RECT 17.120 3049.840 17.380 3050.100 ;
        RECT 1959.700 3049.840 1959.960 3050.100 ;
      LAYER met2 ;
        RECT 17.110 3051.995 17.390 3052.365 ;
        RECT 17.180 3050.130 17.320 3051.995 ;
        RECT 17.120 3049.810 17.380 3050.130 ;
        RECT 1959.700 3049.810 1959.960 3050.130 ;
        RECT 1959.760 2900.610 1959.900 3049.810 ;
        RECT 1959.760 2900.470 1962.660 2900.610 ;
        RECT 1962.520 2899.250 1962.660 2900.470 ;
        RECT 1964.685 2899.250 1964.965 2900.000 ;
        RECT 1962.520 2899.110 1964.965 2899.250 ;
        RECT 1964.685 2896.000 1964.965 2899.110 ;
      LAYER via2 ;
        RECT 17.110 3052.040 17.390 3052.320 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 17.085 3052.330 17.415 3052.345 ;
        RECT -4.800 3052.030 17.415 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 17.085 3052.015 17.415 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 33.190 2916.760 33.510 2916.820 ;
        RECT 1996.010 2916.760 1996.330 2916.820 ;
        RECT 33.190 2916.620 1996.330 2916.760 ;
        RECT 33.190 2916.560 33.510 2916.620 ;
        RECT 1996.010 2916.560 1996.330 2916.620 ;
        RECT 15.710 2766.820 16.030 2766.880 ;
        RECT 33.190 2766.820 33.510 2766.880 ;
        RECT 15.710 2766.680 33.510 2766.820 ;
        RECT 15.710 2766.620 16.030 2766.680 ;
        RECT 33.190 2766.620 33.510 2766.680 ;
      LAYER via ;
        RECT 33.220 2916.560 33.480 2916.820 ;
        RECT 1996.040 2916.560 1996.300 2916.820 ;
        RECT 15.740 2766.620 16.000 2766.880 ;
        RECT 33.220 2766.620 33.480 2766.880 ;
      LAYER met2 ;
        RECT 33.220 2916.530 33.480 2916.850 ;
        RECT 1996.040 2916.530 1996.300 2916.850 ;
        RECT 33.280 2766.910 33.420 2916.530 ;
        RECT 1996.100 2900.000 1996.240 2916.530 ;
        RECT 1995.965 2896.000 1996.245 2900.000 ;
        RECT 15.740 2766.590 16.000 2766.910 ;
        RECT 33.220 2766.590 33.480 2766.910 ;
        RECT 15.800 2765.405 15.940 2766.590 ;
        RECT 15.730 2765.035 16.010 2765.405 ;
      LAYER via2 ;
        RECT 15.730 2765.080 16.010 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 15.705 2765.370 16.035 2765.385 ;
        RECT -4.800 2765.070 16.035 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 15.705 2765.055 16.035 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 23.530 2916.080 23.850 2916.140 ;
        RECT 2027.750 2916.080 2028.070 2916.140 ;
        RECT 23.530 2915.940 2028.070 2916.080 ;
        RECT 23.530 2915.880 23.850 2915.940 ;
        RECT 2027.750 2915.880 2028.070 2915.940 ;
        RECT 13.870 2478.840 14.190 2478.900 ;
        RECT 23.530 2478.840 23.850 2478.900 ;
        RECT 13.870 2478.700 23.850 2478.840 ;
        RECT 13.870 2478.640 14.190 2478.700 ;
        RECT 23.530 2478.640 23.850 2478.700 ;
      LAYER via ;
        RECT 23.560 2915.880 23.820 2916.140 ;
        RECT 2027.780 2915.880 2028.040 2916.140 ;
        RECT 13.900 2478.640 14.160 2478.900 ;
        RECT 23.560 2478.640 23.820 2478.900 ;
      LAYER met2 ;
        RECT 23.560 2915.850 23.820 2916.170 ;
        RECT 2027.780 2915.850 2028.040 2916.170 ;
        RECT 23.620 2478.930 23.760 2915.850 ;
        RECT 2027.840 2900.000 2027.980 2915.850 ;
        RECT 2027.705 2896.000 2027.985 2900.000 ;
        RECT 13.900 2478.610 14.160 2478.930 ;
        RECT 23.560 2478.610 23.820 2478.930 ;
        RECT 13.960 2477.765 14.100 2478.610 ;
        RECT 13.890 2477.395 14.170 2477.765 ;
      LAYER via2 ;
        RECT 13.890 2477.440 14.170 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 13.865 2477.730 14.195 2477.745 ;
        RECT -4.800 2477.430 14.195 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 13.865 2477.415 14.195 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 27.210 2915.060 27.530 2915.120 ;
        RECT 2059.490 2915.060 2059.810 2915.120 ;
        RECT 27.210 2914.920 2059.810 2915.060 ;
        RECT 27.210 2914.860 27.530 2914.920 ;
        RECT 2059.490 2914.860 2059.810 2914.920 ;
        RECT 13.870 2192.900 14.190 2192.960 ;
        RECT 27.210 2192.900 27.530 2192.960 ;
        RECT 13.870 2192.760 27.530 2192.900 ;
        RECT 13.870 2192.700 14.190 2192.760 ;
        RECT 27.210 2192.700 27.530 2192.760 ;
      LAYER via ;
        RECT 27.240 2914.860 27.500 2915.120 ;
        RECT 2059.520 2914.860 2059.780 2915.120 ;
        RECT 13.900 2192.700 14.160 2192.960 ;
        RECT 27.240 2192.700 27.500 2192.960 ;
      LAYER met2 ;
        RECT 27.240 2914.830 27.500 2915.150 ;
        RECT 2059.520 2914.830 2059.780 2915.150 ;
        RECT 27.300 2192.990 27.440 2914.830 ;
        RECT 2059.580 2900.000 2059.720 2914.830 ;
        RECT 2059.445 2896.000 2059.725 2900.000 ;
        RECT 13.900 2192.670 14.160 2192.990 ;
        RECT 27.240 2192.670 27.500 2192.990 ;
        RECT 13.960 2190.125 14.100 2192.670 ;
        RECT 13.890 2189.755 14.170 2190.125 ;
      LAYER via2 ;
        RECT 13.890 2189.800 14.170 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 13.865 2190.090 14.195 2190.105 ;
        RECT -4.800 2189.790 14.195 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 13.865 2189.775 14.195 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 26.290 2914.380 26.610 2914.440 ;
        RECT 2090.770 2914.380 2091.090 2914.440 ;
        RECT 26.290 2914.240 2091.090 2914.380 ;
        RECT 26.290 2914.180 26.610 2914.240 ;
        RECT 2090.770 2914.180 2091.090 2914.240 ;
        RECT 13.870 1903.900 14.190 1903.960 ;
        RECT 26.290 1903.900 26.610 1903.960 ;
        RECT 13.870 1903.760 26.610 1903.900 ;
        RECT 13.870 1903.700 14.190 1903.760 ;
        RECT 26.290 1903.700 26.610 1903.760 ;
      LAYER via ;
        RECT 26.320 2914.180 26.580 2914.440 ;
        RECT 2090.800 2914.180 2091.060 2914.440 ;
        RECT 13.900 1903.700 14.160 1903.960 ;
        RECT 26.320 1903.700 26.580 1903.960 ;
      LAYER met2 ;
        RECT 26.320 2914.150 26.580 2914.470 ;
        RECT 2090.800 2914.150 2091.060 2914.470 ;
        RECT 26.380 1903.990 26.520 2914.150 ;
        RECT 2090.860 2900.000 2091.000 2914.150 ;
        RECT 2090.725 2896.000 2091.005 2900.000 ;
        RECT 13.900 1903.670 14.160 1903.990 ;
        RECT 26.320 1903.670 26.580 1903.990 ;
        RECT 13.960 1903.165 14.100 1903.670 ;
        RECT 13.890 1902.795 14.170 1903.165 ;
      LAYER via2 ;
        RECT 13.890 1902.840 14.170 1903.120 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 13.865 1903.130 14.195 1903.145 ;
        RECT -4.800 1902.830 14.195 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 13.865 1902.815 14.195 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2282.590 615.640 2282.910 615.700 ;
        RECT 2287.190 615.640 2287.510 615.700 ;
        RECT 2282.590 615.500 2287.510 615.640 ;
        RECT 2282.590 615.440 2282.910 615.500 ;
        RECT 2287.190 615.440 2287.510 615.500 ;
        RECT 1530.030 615.300 1530.350 615.360 ;
        RECT 1572.810 615.300 1573.130 615.360 ;
        RECT 1530.030 615.160 1573.130 615.300 ;
        RECT 1530.030 615.100 1530.350 615.160 ;
        RECT 1572.810 615.100 1573.130 615.160 ;
        RECT 1848.350 615.300 1848.670 615.360 ;
        RECT 1883.310 615.300 1883.630 615.360 ;
        RECT 1848.350 615.160 1883.630 615.300 ;
        RECT 1848.350 615.100 1848.670 615.160 ;
        RECT 1883.310 615.100 1883.630 615.160 ;
        RECT 2089.390 614.960 2089.710 615.020 ;
        RECT 2096.750 614.960 2097.070 615.020 ;
        RECT 2089.390 614.820 2097.070 614.960 ;
        RECT 2089.390 614.760 2089.710 614.820 ;
        RECT 2096.750 614.760 2097.070 614.820 ;
        RECT 2185.990 614.960 2186.310 615.020 ;
        RECT 2187.370 614.960 2187.690 615.020 ;
        RECT 2185.990 614.820 2187.690 614.960 ;
        RECT 2185.990 614.760 2186.310 614.820 ;
        RECT 2187.370 614.760 2187.690 614.820 ;
      LAYER via ;
        RECT 2282.620 615.440 2282.880 615.700 ;
        RECT 2287.220 615.440 2287.480 615.700 ;
        RECT 1530.060 615.100 1530.320 615.360 ;
        RECT 1572.840 615.100 1573.100 615.360 ;
        RECT 1848.380 615.100 1848.640 615.360 ;
        RECT 1883.340 615.100 1883.600 615.360 ;
        RECT 2089.420 614.760 2089.680 615.020 ;
        RECT 2096.780 614.760 2097.040 615.020 ;
        RECT 2186.020 614.760 2186.280 615.020 ;
        RECT 2187.400 614.760 2187.660 615.020 ;
      LAYER met2 ;
        RECT 1238.345 2896.530 1238.625 2900.000 ;
        RECT 1239.330 2896.530 1239.610 2896.645 ;
        RECT 1238.345 2896.390 1239.610 2896.530 ;
        RECT 1238.345 2896.000 1238.625 2896.390 ;
        RECT 1239.330 2896.275 1239.610 2896.390 ;
        RECT 1628.030 617.595 1628.310 617.965 ;
        RECT 1368.590 616.490 1368.870 616.605 ;
        RECT 1369.510 616.490 1369.790 616.605 ;
        RECT 1368.590 616.350 1369.790 616.490 ;
        RECT 1368.590 616.235 1368.870 616.350 ;
        RECT 1369.510 616.235 1369.790 616.350 ;
        RECT 1482.670 616.235 1482.950 616.605 ;
        RECT 1572.830 616.235 1573.110 616.605 ;
        RECT 1482.740 615.245 1482.880 616.235 ;
        RECT 1572.900 615.390 1573.040 616.235 ;
        RECT 1530.060 615.245 1530.320 615.390 ;
        RECT 1482.670 614.875 1482.950 615.245 ;
        RECT 1530.050 614.875 1530.330 615.245 ;
        RECT 1572.840 615.070 1573.100 615.390 ;
        RECT 1628.100 615.245 1628.240 617.595 ;
        RECT 2439.010 616.235 2439.290 616.605 ;
        RECT 1642.290 615.555 1642.570 615.925 ;
        RECT 1883.330 615.555 1883.610 615.925 ;
        RECT 2282.610 615.555 2282.890 615.925 ;
        RECT 1642.360 615.245 1642.500 615.555 ;
        RECT 1883.400 615.390 1883.540 615.555 ;
        RECT 2282.620 615.410 2282.880 615.555 ;
        RECT 2287.220 615.410 2287.480 615.730 ;
        RECT 2359.430 615.555 2359.710 615.925 ;
        RECT 2380.130 615.555 2380.410 615.925 ;
        RECT 1628.030 614.875 1628.310 615.245 ;
        RECT 1642.290 614.875 1642.570 615.245 ;
        RECT 1828.130 614.875 1828.410 615.245 ;
        RECT 1848.380 615.070 1848.640 615.390 ;
        RECT 1883.340 615.070 1883.600 615.390 ;
        RECT 2287.280 615.245 2287.420 615.410 ;
        RECT 1828.200 614.565 1828.340 614.875 ;
        RECT 1848.440 614.565 1848.580 615.070 ;
        RECT 2089.410 614.875 2089.690 615.245 ;
        RECT 2096.770 614.875 2097.050 615.245 ;
        RECT 2186.010 614.875 2186.290 615.245 ;
        RECT 2187.390 614.875 2187.670 615.245 ;
        RECT 2287.210 614.875 2287.490 615.245 ;
        RECT 2089.420 614.730 2089.680 614.875 ;
        RECT 2096.780 614.730 2097.040 614.875 ;
        RECT 2186.020 614.730 2186.280 614.875 ;
        RECT 2187.400 614.730 2187.660 614.875 ;
        RECT 1828.130 614.195 1828.410 614.565 ;
        RECT 1848.370 614.195 1848.650 614.565 ;
        RECT 2359.500 613.885 2359.640 615.555 ;
        RECT 2380.200 615.130 2380.340 615.555 ;
        RECT 2381.050 615.130 2381.330 615.245 ;
        RECT 2380.200 614.990 2381.330 615.130 ;
        RECT 2381.050 614.875 2381.330 614.990 ;
        RECT 2439.080 614.565 2439.220 616.235 ;
        RECT 2439.010 614.195 2439.290 614.565 ;
        RECT 2359.430 613.515 2359.710 613.885 ;
      LAYER via2 ;
        RECT 1239.330 2896.320 1239.610 2896.600 ;
        RECT 1628.030 617.640 1628.310 617.920 ;
        RECT 1368.590 616.280 1368.870 616.560 ;
        RECT 1369.510 616.280 1369.790 616.560 ;
        RECT 1482.670 616.280 1482.950 616.560 ;
        RECT 1572.830 616.280 1573.110 616.560 ;
        RECT 1482.670 614.920 1482.950 615.200 ;
        RECT 1530.050 614.920 1530.330 615.200 ;
        RECT 2439.010 616.280 2439.290 616.560 ;
        RECT 1642.290 615.600 1642.570 615.880 ;
        RECT 1883.330 615.600 1883.610 615.880 ;
        RECT 2282.610 615.600 2282.890 615.880 ;
        RECT 2359.430 615.600 2359.710 615.880 ;
        RECT 2380.130 615.600 2380.410 615.880 ;
        RECT 1628.030 614.920 1628.310 615.200 ;
        RECT 1642.290 614.920 1642.570 615.200 ;
        RECT 1828.130 614.920 1828.410 615.200 ;
        RECT 2089.410 614.920 2089.690 615.200 ;
        RECT 2096.770 614.920 2097.050 615.200 ;
        RECT 2186.010 614.920 2186.290 615.200 ;
        RECT 2187.390 614.920 2187.670 615.200 ;
        RECT 2287.210 614.920 2287.490 615.200 ;
        RECT 1828.130 614.240 1828.410 614.520 ;
        RECT 1848.370 614.240 1848.650 614.520 ;
        RECT 2381.050 614.920 2381.330 615.200 ;
        RECT 2439.010 614.240 2439.290 614.520 ;
        RECT 2359.430 613.560 2359.710 613.840 ;
      LAYER met3 ;
        RECT 1239.305 2896.610 1239.635 2896.625 ;
        RECT 1241.350 2896.610 1241.730 2896.620 ;
        RECT 1239.305 2896.310 1241.730 2896.610 ;
        RECT 1239.305 2896.295 1239.635 2896.310 ;
        RECT 1241.350 2896.300 1241.730 2896.310 ;
        RECT 1579.910 617.930 1580.290 617.940 ;
        RECT 1628.005 617.930 1628.335 617.945 ;
        RECT 1579.910 617.630 1628.335 617.930 ;
        RECT 1579.910 617.620 1580.290 617.630 ;
        RECT 1628.005 617.615 1628.335 617.630 ;
        RECT 1338.870 616.570 1339.250 616.580 ;
        RECT 1368.565 616.570 1368.895 616.585 ;
        RECT 1338.870 616.270 1368.895 616.570 ;
        RECT 1338.870 616.260 1339.250 616.270 ;
        RECT 1368.565 616.255 1368.895 616.270 ;
        RECT 1369.485 616.570 1369.815 616.585 ;
        RECT 1482.645 616.570 1482.975 616.585 ;
        RECT 1369.485 616.270 1482.975 616.570 ;
        RECT 1369.485 616.255 1369.815 616.270 ;
        RECT 1482.645 616.255 1482.975 616.270 ;
        RECT 1572.805 616.570 1573.135 616.585 ;
        RECT 1579.910 616.570 1580.290 616.580 ;
        RECT 2438.985 616.570 2439.315 616.585 ;
        RECT 1572.805 616.270 1580.290 616.570 ;
        RECT 1572.805 616.255 1573.135 616.270 ;
        RECT 1579.910 616.260 1580.290 616.270 ;
        RECT 1993.030 616.270 2028.290 616.570 ;
        RECT 1241.350 615.890 1241.730 615.900 ;
        RECT 1642.265 615.890 1642.595 615.905 ;
        RECT 1883.305 615.890 1883.635 615.905 ;
        RECT 1241.350 615.590 1270.210 615.890 ;
        RECT 1241.350 615.580 1241.730 615.590 ;
        RECT 1269.910 615.210 1270.210 615.590 ;
        RECT 1642.265 615.590 1704.450 615.890 ;
        RECT 1642.265 615.575 1642.595 615.590 ;
        RECT 1338.870 615.210 1339.250 615.220 ;
        RECT 1269.910 614.910 1339.250 615.210 ;
        RECT 1338.870 614.900 1339.250 614.910 ;
        RECT 1482.645 615.210 1482.975 615.225 ;
        RECT 1530.025 615.210 1530.355 615.225 ;
        RECT 1482.645 614.910 1530.355 615.210 ;
        RECT 1482.645 614.895 1482.975 614.910 ;
        RECT 1530.025 614.895 1530.355 614.910 ;
        RECT 1628.005 615.210 1628.335 615.225 ;
        RECT 1642.265 615.210 1642.595 615.225 ;
        RECT 1628.005 614.910 1642.595 615.210 ;
        RECT 1628.005 614.895 1628.335 614.910 ;
        RECT 1642.265 614.895 1642.595 614.910 ;
        RECT 1704.150 614.530 1704.450 615.590 ;
        RECT 1883.305 615.590 1897.650 615.890 ;
        RECT 1883.305 615.575 1883.635 615.590 ;
        RECT 1828.105 615.210 1828.435 615.225 ;
        RECT 1752.910 614.910 1828.435 615.210 ;
        RECT 1752.910 614.530 1753.210 614.910 ;
        RECT 1828.105 614.895 1828.435 614.910 ;
        RECT 1704.150 614.230 1753.210 614.530 ;
        RECT 1828.105 614.530 1828.435 614.545 ;
        RECT 1848.345 614.530 1848.675 614.545 ;
        RECT 1828.105 614.230 1848.675 614.530 ;
        RECT 1897.350 614.530 1897.650 615.590 ;
        RECT 1993.030 615.210 1993.330 616.270 ;
        RECT 1942.430 614.910 1993.330 615.210 ;
        RECT 1942.430 614.530 1942.730 614.910 ;
        RECT 1897.350 614.230 1942.730 614.530 ;
        RECT 2027.990 614.530 2028.290 616.270 ;
        RECT 2415.310 616.270 2439.315 616.570 ;
        RECT 2282.585 615.890 2282.915 615.905 ;
        RECT 2235.910 615.590 2282.915 615.890 ;
        RECT 2089.385 615.210 2089.715 615.225 ;
        RECT 2042.710 614.910 2089.715 615.210 ;
        RECT 2042.710 614.530 2043.010 614.910 ;
        RECT 2089.385 614.895 2089.715 614.910 ;
        RECT 2096.745 615.210 2097.075 615.225 ;
        RECT 2185.985 615.210 2186.315 615.225 ;
        RECT 2096.745 614.910 2124.890 615.210 ;
        RECT 2096.745 614.895 2097.075 614.910 ;
        RECT 2027.990 614.230 2043.010 614.530 ;
        RECT 2124.590 614.530 2124.890 614.910 ;
        RECT 2139.310 614.910 2186.315 615.210 ;
        RECT 2139.310 614.530 2139.610 614.910 ;
        RECT 2185.985 614.895 2186.315 614.910 ;
        RECT 2187.365 615.210 2187.695 615.225 ;
        RECT 2187.365 614.910 2221.490 615.210 ;
        RECT 2187.365 614.895 2187.695 614.910 ;
        RECT 2124.590 614.230 2139.610 614.530 ;
        RECT 2221.190 614.530 2221.490 614.910 ;
        RECT 2235.910 614.530 2236.210 615.590 ;
        RECT 2282.585 615.575 2282.915 615.590 ;
        RECT 2359.405 615.890 2359.735 615.905 ;
        RECT 2380.105 615.890 2380.435 615.905 ;
        RECT 2359.405 615.590 2380.435 615.890 ;
        RECT 2359.405 615.575 2359.735 615.590 ;
        RECT 2380.105 615.575 2380.435 615.590 ;
        RECT 2287.185 615.210 2287.515 615.225 ;
        RECT 2311.310 615.210 2311.690 615.220 ;
        RECT 2287.185 614.910 2311.690 615.210 ;
        RECT 2287.185 614.895 2287.515 614.910 ;
        RECT 2311.310 614.900 2311.690 614.910 ;
        RECT 2381.025 615.210 2381.355 615.225 ;
        RECT 2415.310 615.210 2415.610 616.270 ;
        RECT 2438.985 616.255 2439.315 616.270 ;
        RECT 2463.110 615.890 2463.490 615.900 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2463.110 615.590 2546.250 615.890 ;
        RECT 2463.110 615.580 2463.490 615.590 ;
        RECT 2381.025 614.910 2415.610 615.210 ;
        RECT 2545.950 615.210 2546.250 615.590 ;
        RECT 2594.710 615.590 2642.850 615.890 ;
        RECT 2545.950 614.910 2594.090 615.210 ;
        RECT 2381.025 614.895 2381.355 614.910 ;
        RECT 2221.190 614.230 2236.210 614.530 ;
        RECT 2438.985 614.530 2439.315 614.545 ;
        RECT 2463.110 614.530 2463.490 614.540 ;
        RECT 2438.985 614.230 2463.490 614.530 ;
        RECT 2593.790 614.530 2594.090 614.910 ;
        RECT 2594.710 614.530 2595.010 615.590 ;
        RECT 2642.550 615.210 2642.850 615.590 ;
        RECT 2691.310 615.590 2739.450 615.890 ;
        RECT 2642.550 614.910 2690.690 615.210 ;
        RECT 2593.790 614.230 2595.010 614.530 ;
        RECT 2690.390 614.530 2690.690 614.910 ;
        RECT 2691.310 614.530 2691.610 615.590 ;
        RECT 2739.150 615.210 2739.450 615.590 ;
        RECT 2787.910 615.590 2836.050 615.890 ;
        RECT 2739.150 614.910 2787.290 615.210 ;
        RECT 2690.390 614.230 2691.610 614.530 ;
        RECT 2786.990 614.530 2787.290 614.910 ;
        RECT 2787.910 614.530 2788.210 615.590 ;
        RECT 2835.750 615.210 2836.050 615.590 ;
        RECT 2916.710 615.590 2924.800 615.890 ;
        RECT 2916.710 615.210 2917.010 615.590 ;
        RECT 2835.750 614.910 2883.890 615.210 ;
        RECT 2786.990 614.230 2788.210 614.530 ;
        RECT 2883.590 614.530 2883.890 614.910 ;
        RECT 2884.510 614.910 2917.010 615.210 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
        RECT 2884.510 614.530 2884.810 614.910 ;
        RECT 2883.590 614.230 2884.810 614.530 ;
        RECT 1828.105 614.215 1828.435 614.230 ;
        RECT 1848.345 614.215 1848.675 614.230 ;
        RECT 2438.985 614.215 2439.315 614.230 ;
        RECT 2463.110 614.220 2463.490 614.230 ;
        RECT 2311.310 613.850 2311.690 613.860 ;
        RECT 2359.405 613.850 2359.735 613.865 ;
        RECT 2311.310 613.550 2359.735 613.850 ;
        RECT 2311.310 613.540 2311.690 613.550 ;
        RECT 2359.405 613.535 2359.735 613.550 ;
      LAYER via3 ;
        RECT 1241.380 2896.300 1241.700 2896.620 ;
        RECT 1579.940 617.620 1580.260 617.940 ;
        RECT 1338.900 616.260 1339.220 616.580 ;
        RECT 1579.940 616.260 1580.260 616.580 ;
        RECT 1241.380 615.580 1241.700 615.900 ;
        RECT 1338.900 614.900 1339.220 615.220 ;
        RECT 2311.340 614.900 2311.660 615.220 ;
        RECT 2463.140 615.580 2463.460 615.900 ;
        RECT 2463.140 614.220 2463.460 614.540 ;
        RECT 2311.340 613.540 2311.660 613.860 ;
      LAYER met4 ;
        RECT 1241.375 2896.295 1241.705 2896.625 ;
        RECT 1241.390 615.905 1241.690 2896.295 ;
        RECT 1579.935 617.615 1580.265 617.945 ;
        RECT 1579.950 616.585 1580.250 617.615 ;
        RECT 1338.895 616.255 1339.225 616.585 ;
        RECT 1579.935 616.255 1580.265 616.585 ;
        RECT 1241.375 615.575 1241.705 615.905 ;
        RECT 1338.910 615.225 1339.210 616.255 ;
        RECT 2463.135 615.575 2463.465 615.905 ;
        RECT 1338.895 614.895 1339.225 615.225 ;
        RECT 2311.335 614.895 2311.665 615.225 ;
        RECT 2311.350 613.865 2311.650 614.895 ;
        RECT 2463.150 614.545 2463.450 615.575 ;
        RECT 2463.135 614.215 2463.465 614.545 ;
        RECT 2311.335 613.535 2311.665 613.865 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 72.290 2914.720 72.610 2914.780 ;
        RECT 2122.510 2914.720 2122.830 2914.780 ;
        RECT 72.290 2914.580 2122.830 2914.720 ;
        RECT 72.290 2914.520 72.610 2914.580 ;
        RECT 2122.510 2914.520 2122.830 2914.580 ;
        RECT 16.630 1621.360 16.950 1621.420 ;
        RECT 72.290 1621.360 72.610 1621.420 ;
        RECT 16.630 1621.220 72.610 1621.360 ;
        RECT 16.630 1621.160 16.950 1621.220 ;
        RECT 72.290 1621.160 72.610 1621.220 ;
      LAYER via ;
        RECT 72.320 2914.520 72.580 2914.780 ;
        RECT 2122.540 2914.520 2122.800 2914.780 ;
        RECT 16.660 1621.160 16.920 1621.420 ;
        RECT 72.320 1621.160 72.580 1621.420 ;
      LAYER met2 ;
        RECT 72.320 2914.490 72.580 2914.810 ;
        RECT 2122.540 2914.490 2122.800 2914.810 ;
        RECT 72.380 1621.450 72.520 2914.490 ;
        RECT 2122.600 2900.000 2122.740 2914.490 ;
        RECT 2122.465 2896.000 2122.745 2900.000 ;
        RECT 16.660 1621.130 16.920 1621.450 ;
        RECT 72.320 1621.130 72.580 1621.450 ;
        RECT 16.720 1615.525 16.860 1621.130 ;
        RECT 16.650 1615.155 16.930 1615.525 ;
      LAYER via2 ;
        RECT 16.650 1615.200 16.930 1615.480 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 16.625 1615.490 16.955 1615.505 ;
        RECT -4.800 1615.190 16.955 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 16.625 1615.175 16.955 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 79.190 2914.040 79.510 2914.100 ;
        RECT 2154.250 2914.040 2154.570 2914.100 ;
        RECT 79.190 2913.900 2154.570 2914.040 ;
        RECT 79.190 2913.840 79.510 2913.900 ;
        RECT 2154.250 2913.840 2154.570 2913.900 ;
        RECT 16.630 1400.700 16.950 1400.760 ;
        RECT 79.190 1400.700 79.510 1400.760 ;
        RECT 16.630 1400.560 79.510 1400.700 ;
        RECT 16.630 1400.500 16.950 1400.560 ;
        RECT 79.190 1400.500 79.510 1400.560 ;
      LAYER via ;
        RECT 79.220 2913.840 79.480 2914.100 ;
        RECT 2154.280 2913.840 2154.540 2914.100 ;
        RECT 16.660 1400.500 16.920 1400.760 ;
        RECT 79.220 1400.500 79.480 1400.760 ;
      LAYER met2 ;
        RECT 79.220 2913.810 79.480 2914.130 ;
        RECT 2154.280 2913.810 2154.540 2914.130 ;
        RECT 79.280 1400.790 79.420 2913.810 ;
        RECT 2154.340 2900.000 2154.480 2913.810 ;
        RECT 2154.205 2896.000 2154.485 2900.000 ;
        RECT 16.660 1400.645 16.920 1400.790 ;
        RECT 16.650 1400.275 16.930 1400.645 ;
        RECT 79.220 1400.470 79.480 1400.790 ;
      LAYER via2 ;
        RECT 16.650 1400.320 16.930 1400.600 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 16.625 1400.610 16.955 1400.625 ;
        RECT -4.800 1400.310 16.955 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 16.625 1400.295 16.955 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 86.090 2913.360 86.410 2913.420 ;
        RECT 2185.530 2913.360 2185.850 2913.420 ;
        RECT 86.090 2913.220 2185.850 2913.360 ;
        RECT 86.090 2913.160 86.410 2913.220 ;
        RECT 2185.530 2913.160 2185.850 2913.220 ;
        RECT 16.630 1186.840 16.950 1186.900 ;
        RECT 86.090 1186.840 86.410 1186.900 ;
        RECT 16.630 1186.700 86.410 1186.840 ;
        RECT 16.630 1186.640 16.950 1186.700 ;
        RECT 86.090 1186.640 86.410 1186.700 ;
      LAYER via ;
        RECT 86.120 2913.160 86.380 2913.420 ;
        RECT 2185.560 2913.160 2185.820 2913.420 ;
        RECT 16.660 1186.640 16.920 1186.900 ;
        RECT 86.120 1186.640 86.380 1186.900 ;
      LAYER met2 ;
        RECT 86.120 2913.130 86.380 2913.450 ;
        RECT 2185.560 2913.130 2185.820 2913.450 ;
        RECT 86.180 1186.930 86.320 2913.130 ;
        RECT 2185.620 2900.000 2185.760 2913.130 ;
        RECT 2185.485 2896.000 2185.765 2900.000 ;
        RECT 16.660 1186.610 16.920 1186.930 ;
        RECT 86.120 1186.610 86.380 1186.930 ;
        RECT 16.720 1185.085 16.860 1186.610 ;
        RECT 16.650 1184.715 16.930 1185.085 ;
      LAYER via2 ;
        RECT 16.650 1184.760 16.930 1185.040 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 16.625 1185.050 16.955 1185.065 ;
        RECT -4.800 1184.750 16.955 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 16.625 1184.735 16.955 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 2912.340 18.790 2912.400 ;
        RECT 2217.270 2912.340 2217.590 2912.400 ;
        RECT 18.470 2912.200 2217.590 2912.340 ;
        RECT 18.470 2912.140 18.790 2912.200 ;
        RECT 2217.270 2912.140 2217.590 2912.200 ;
      LAYER via ;
        RECT 18.500 2912.140 18.760 2912.400 ;
        RECT 2217.300 2912.140 2217.560 2912.400 ;
      LAYER met2 ;
        RECT 18.500 2912.110 18.760 2912.430 ;
        RECT 2217.300 2912.110 2217.560 2912.430 ;
        RECT 18.560 969.525 18.700 2912.110 ;
        RECT 2217.360 2900.000 2217.500 2912.110 ;
        RECT 2217.225 2896.000 2217.505 2900.000 ;
        RECT 18.490 969.155 18.770 969.525 ;
      LAYER via2 ;
        RECT 18.490 969.200 18.770 969.480 ;
      LAYER met3 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 18.465 969.490 18.795 969.505 ;
        RECT -4.800 969.190 18.795 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 18.465 969.175 18.795 969.190 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 120.590 2913.020 120.910 2913.080 ;
        RECT 2249.010 2913.020 2249.330 2913.080 ;
        RECT 120.590 2912.880 2249.330 2913.020 ;
        RECT 120.590 2912.820 120.910 2912.880 ;
        RECT 2249.010 2912.820 2249.330 2912.880 ;
        RECT 16.630 758.780 16.950 758.840 ;
        RECT 120.590 758.780 120.910 758.840 ;
        RECT 16.630 758.640 120.910 758.780 ;
        RECT 16.630 758.580 16.950 758.640 ;
        RECT 120.590 758.580 120.910 758.640 ;
      LAYER via ;
        RECT 120.620 2912.820 120.880 2913.080 ;
        RECT 2249.040 2912.820 2249.300 2913.080 ;
        RECT 16.660 758.580 16.920 758.840 ;
        RECT 120.620 758.580 120.880 758.840 ;
      LAYER met2 ;
        RECT 120.620 2912.790 120.880 2913.110 ;
        RECT 2249.040 2912.790 2249.300 2913.110 ;
        RECT 120.680 758.870 120.820 2912.790 ;
        RECT 2249.100 2900.000 2249.240 2912.790 ;
        RECT 2248.965 2896.000 2249.245 2900.000 ;
        RECT 16.660 758.550 16.920 758.870 ;
        RECT 120.620 758.550 120.880 758.870 ;
        RECT 16.720 753.965 16.860 758.550 ;
        RECT 16.650 753.595 16.930 753.965 ;
      LAYER via2 ;
        RECT 16.650 753.640 16.930 753.920 ;
      LAYER met3 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 16.625 753.930 16.955 753.945 ;
        RECT -4.800 753.630 16.955 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 16.625 753.615 16.955 753.630 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2278.985 2891.105 2279.155 2896.715 ;
      LAYER mcon ;
        RECT 2278.985 2896.545 2279.155 2896.715 ;
      LAYER met1 ;
        RECT 2278.910 2896.700 2279.230 2896.760 ;
        RECT 2278.715 2896.560 2279.230 2896.700 ;
        RECT 2278.910 2896.500 2279.230 2896.560 ;
        RECT 17.550 2891.260 17.870 2891.320 ;
        RECT 2278.925 2891.260 2279.215 2891.305 ;
        RECT 17.550 2891.120 2279.215 2891.260 ;
        RECT 17.550 2891.060 17.870 2891.120 ;
        RECT 2278.925 2891.075 2279.215 2891.120 ;
      LAYER via ;
        RECT 2278.940 2896.500 2279.200 2896.760 ;
        RECT 17.580 2891.060 17.840 2891.320 ;
      LAYER met2 ;
        RECT 2278.940 2896.530 2279.200 2896.790 ;
        RECT 2280.245 2896.530 2280.525 2900.000 ;
        RECT 2278.940 2896.470 2280.525 2896.530 ;
        RECT 2279.000 2896.390 2280.525 2896.470 ;
        RECT 2280.245 2896.000 2280.525 2896.390 ;
        RECT 17.580 2891.030 17.840 2891.350 ;
        RECT 17.640 538.405 17.780 2891.030 ;
        RECT 17.570 538.035 17.850 538.405 ;
      LAYER via2 ;
        RECT 17.570 538.080 17.850 538.360 ;
      LAYER met3 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 17.545 538.370 17.875 538.385 ;
        RECT -4.800 538.070 17.875 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 17.545 538.055 17.875 538.070 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 324.260 16.950 324.320 ;
        RECT 155.090 324.260 155.410 324.320 ;
        RECT 16.630 324.120 155.410 324.260 ;
        RECT 16.630 324.060 16.950 324.120 ;
        RECT 155.090 324.060 155.410 324.120 ;
      LAYER via ;
        RECT 16.660 324.060 16.920 324.320 ;
        RECT 155.120 324.060 155.380 324.320 ;
      LAYER met2 ;
        RECT 155.110 2912.595 155.390 2912.965 ;
        RECT 2312.050 2912.595 2312.330 2912.965 ;
        RECT 155.180 324.350 155.320 2912.595 ;
        RECT 2312.120 2900.000 2312.260 2912.595 ;
        RECT 2311.985 2896.000 2312.265 2900.000 ;
        RECT 16.660 324.030 16.920 324.350 ;
        RECT 155.120 324.030 155.380 324.350 ;
        RECT 16.720 322.845 16.860 324.030 ;
        RECT 16.650 322.475 16.930 322.845 ;
      LAYER via2 ;
        RECT 155.110 2912.640 155.390 2912.920 ;
        RECT 2312.050 2912.640 2312.330 2912.920 ;
        RECT 16.650 322.520 16.930 322.800 ;
      LAYER met3 ;
        RECT 155.085 2912.930 155.415 2912.945 ;
        RECT 2312.025 2912.930 2312.355 2912.945 ;
        RECT 155.085 2912.630 2312.355 2912.930 ;
        RECT 155.085 2912.615 155.415 2912.630 ;
        RECT 2312.025 2912.615 2312.355 2912.630 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 16.625 322.810 16.955 322.825 ;
        RECT -4.800 322.510 16.955 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
        RECT 16.625 322.495 16.955 322.510 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2342.870 2896.530 2343.150 2896.645 ;
        RECT 2343.725 2896.530 2344.005 2900.000 ;
        RECT 2342.870 2896.390 2344.005 2896.530 ;
        RECT 2342.870 2896.275 2343.150 2896.390 ;
        RECT 2343.725 2896.000 2344.005 2896.390 ;
      LAYER via2 ;
        RECT 2342.870 2896.320 2343.150 2896.600 ;
      LAYER met3 ;
        RECT 2338.910 2896.610 2339.290 2896.620 ;
        RECT 2342.845 2896.610 2343.175 2896.625 ;
        RECT 2338.910 2896.310 2343.175 2896.610 ;
        RECT 2338.910 2896.300 2339.290 2896.310 ;
        RECT 2342.845 2896.295 2343.175 2896.310 ;
        RECT 2338.910 109.970 2339.290 109.980 ;
        RECT 3.070 109.670 2339.290 109.970 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 3.070 107.250 3.370 109.670 ;
        RECT 2338.910 109.660 2339.290 109.670 ;
        RECT -4.800 106.950 3.370 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
      LAYER via3 ;
        RECT 2338.940 2896.300 2339.260 2896.620 ;
        RECT 2338.940 109.660 2339.260 109.980 ;
      LAYER met4 ;
        RECT 2338.935 2896.295 2339.265 2896.625 ;
        RECT 2338.950 109.985 2339.250 2896.295 ;
        RECT 2338.935 109.655 2339.265 109.985 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1270.590 2896.500 1270.910 2896.760 ;
        RECT 1270.680 2893.300 1270.820 2896.500 ;
        RECT 2901.290 2893.300 2901.610 2893.360 ;
        RECT 1270.680 2893.160 2901.610 2893.300 ;
        RECT 2901.290 2893.100 2901.610 2893.160 ;
      LAYER via ;
        RECT 1270.620 2896.500 1270.880 2896.760 ;
        RECT 2901.320 2893.100 2901.580 2893.360 ;
      LAYER met2 ;
        RECT 1269.625 2896.530 1269.905 2900.000 ;
        RECT 1270.620 2896.530 1270.880 2896.790 ;
        RECT 1269.625 2896.470 1270.880 2896.530 ;
        RECT 1269.625 2896.390 1270.820 2896.470 ;
        RECT 1269.625 2896.000 1269.905 2896.390 ;
        RECT 2901.320 2893.070 2901.580 2893.390 ;
        RECT 2901.380 850.525 2901.520 2893.070 ;
        RECT 2901.310 850.155 2901.590 850.525 ;
      LAYER via2 ;
        RECT 2901.310 850.200 2901.590 850.480 ;
      LAYER met3 ;
        RECT 2901.285 850.490 2901.615 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2901.285 850.190 2924.800 850.490 ;
        RECT 2901.285 850.175 2901.615 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.250 2896.500 1303.570 2896.760 ;
        RECT 1303.340 2893.640 1303.480 2896.500 ;
        RECT 2902.670 2893.640 2902.990 2893.700 ;
        RECT 1303.340 2893.500 2902.990 2893.640 ;
        RECT 2902.670 2893.440 2902.990 2893.500 ;
      LAYER via ;
        RECT 1303.280 2896.500 1303.540 2896.760 ;
        RECT 2902.700 2893.440 2902.960 2893.700 ;
      LAYER met2 ;
        RECT 1301.365 2896.530 1301.645 2900.000 ;
        RECT 1303.280 2896.530 1303.540 2896.790 ;
        RECT 1301.365 2896.470 1303.540 2896.530 ;
        RECT 1301.365 2896.390 1303.480 2896.470 ;
        RECT 1301.365 2896.000 1301.645 2896.390 ;
        RECT 2902.700 2893.410 2902.960 2893.730 ;
        RECT 2902.760 1085.125 2902.900 2893.410 ;
        RECT 2902.690 1084.755 2902.970 1085.125 ;
      LAYER via2 ;
        RECT 2902.690 1084.800 2902.970 1085.080 ;
      LAYER met3 ;
        RECT 2902.665 1085.090 2902.995 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2902.665 1084.790 2924.800 1085.090 ;
        RECT 2902.665 1084.775 2902.995 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1334.070 2896.500 1334.390 2896.760 ;
        RECT 1334.160 2893.980 1334.300 2896.500 ;
        RECT 2904.050 2893.980 2904.370 2894.040 ;
        RECT 1334.160 2893.840 2904.370 2893.980 ;
        RECT 2904.050 2893.780 2904.370 2893.840 ;
      LAYER via ;
        RECT 1334.100 2896.500 1334.360 2896.760 ;
        RECT 2904.080 2893.780 2904.340 2894.040 ;
      LAYER met2 ;
        RECT 1333.105 2896.530 1333.385 2900.000 ;
        RECT 1334.100 2896.530 1334.360 2896.790 ;
        RECT 1333.105 2896.470 1334.360 2896.530 ;
        RECT 1333.105 2896.390 1334.300 2896.470 ;
        RECT 1333.105 2896.000 1333.385 2896.390 ;
        RECT 2904.080 2893.750 2904.340 2894.070 ;
        RECT 2904.140 1319.725 2904.280 2893.750 ;
        RECT 2904.070 1319.355 2904.350 1319.725 ;
      LAYER via2 ;
        RECT 2904.070 1319.400 2904.350 1319.680 ;
      LAYER met3 ;
        RECT 2904.045 1319.690 2904.375 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2904.045 1319.390 2924.800 1319.690 ;
        RECT 2904.045 1319.375 2904.375 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1365.810 2896.500 1366.130 2896.760 ;
        RECT 1365.900 2894.320 1366.040 2896.500 ;
        RECT 2900.830 2894.320 2901.150 2894.380 ;
        RECT 1365.900 2894.180 2901.150 2894.320 ;
        RECT 2900.830 2894.120 2901.150 2894.180 ;
      LAYER via ;
        RECT 1365.840 2896.500 1366.100 2896.760 ;
        RECT 2900.860 2894.120 2901.120 2894.380 ;
      LAYER met2 ;
        RECT 1364.385 2896.530 1364.665 2900.000 ;
        RECT 1365.840 2896.530 1366.100 2896.790 ;
        RECT 1364.385 2896.470 1366.100 2896.530 ;
        RECT 1364.385 2896.390 1366.040 2896.470 ;
        RECT 1364.385 2896.000 1364.665 2896.390 ;
        RECT 2900.860 2894.090 2901.120 2894.410 ;
        RECT 2900.920 1554.325 2901.060 2894.090 ;
        RECT 2900.850 1553.955 2901.130 1554.325 ;
      LAYER via2 ;
        RECT 2900.850 1554.000 2901.130 1554.280 ;
      LAYER met3 ;
        RECT 2900.825 1554.290 2901.155 1554.305 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2900.825 1553.990 2924.800 1554.290 ;
        RECT 2900.825 1553.975 2901.155 1553.990 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1398.010 2896.500 1398.330 2896.760 ;
        RECT 1398.100 2895.000 1398.240 2896.500 ;
        RECT 2900.370 2895.000 2900.690 2895.060 ;
        RECT 1398.100 2894.860 2900.690 2895.000 ;
        RECT 2900.370 2894.800 2900.690 2894.860 ;
      LAYER via ;
        RECT 1398.040 2896.500 1398.300 2896.760 ;
        RECT 2900.400 2894.800 2900.660 2895.060 ;
      LAYER met2 ;
        RECT 1396.125 2896.530 1396.405 2900.000 ;
        RECT 1398.040 2896.530 1398.300 2896.790 ;
        RECT 1396.125 2896.470 1398.300 2896.530 ;
        RECT 1396.125 2896.390 1398.240 2896.470 ;
        RECT 1396.125 2896.000 1396.405 2896.390 ;
        RECT 2900.400 2894.770 2900.660 2895.090 ;
        RECT 2900.460 1789.605 2900.600 2894.770 ;
        RECT 2900.390 1789.235 2900.670 1789.605 ;
      LAYER via2 ;
        RECT 2900.390 1789.280 2900.670 1789.560 ;
      LAYER met3 ;
        RECT 2900.365 1789.570 2900.695 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2900.365 1789.270 2924.800 1789.570 ;
        RECT 2900.365 1789.255 2900.695 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1428.830 2896.500 1429.150 2896.760 ;
        RECT 1428.920 2896.020 1429.060 2896.500 ;
        RECT 2351.130 2896.020 2351.450 2896.080 ;
        RECT 1428.920 2895.880 2351.450 2896.020 ;
        RECT 2351.130 2895.820 2351.450 2895.880 ;
        RECT 2351.130 2028.340 2351.450 2028.400 ;
        RECT 2899.450 2028.340 2899.770 2028.400 ;
        RECT 2351.130 2028.200 2899.770 2028.340 ;
        RECT 2351.130 2028.140 2351.450 2028.200 ;
        RECT 2899.450 2028.140 2899.770 2028.200 ;
      LAYER via ;
        RECT 1428.860 2896.500 1429.120 2896.760 ;
        RECT 2351.160 2895.820 2351.420 2896.080 ;
        RECT 2351.160 2028.140 2351.420 2028.400 ;
        RECT 2899.480 2028.140 2899.740 2028.400 ;
      LAYER met2 ;
        RECT 1427.865 2896.530 1428.145 2900.000 ;
        RECT 1428.860 2896.530 1429.120 2896.790 ;
        RECT 1427.865 2896.470 1429.120 2896.530 ;
        RECT 1427.865 2896.390 1429.060 2896.470 ;
        RECT 1427.865 2896.000 1428.145 2896.390 ;
        RECT 2351.160 2895.790 2351.420 2896.110 ;
        RECT 2351.220 2028.430 2351.360 2895.790 ;
        RECT 2351.160 2028.110 2351.420 2028.430 ;
        RECT 2899.480 2028.110 2899.740 2028.430 ;
        RECT 2899.540 2024.205 2899.680 2028.110 ;
        RECT 2899.470 2023.835 2899.750 2024.205 ;
      LAYER via2 ;
        RECT 2899.470 2023.880 2899.750 2024.160 ;
      LAYER met3 ;
        RECT 2899.445 2024.170 2899.775 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2899.445 2023.870 2924.800 2024.170 ;
        RECT 2899.445 2023.855 2899.775 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1460.645 2895.185 1460.815 2896.715 ;
      LAYER mcon ;
        RECT 1460.645 2896.545 1460.815 2896.715 ;
      LAYER met1 ;
        RECT 1460.570 2896.700 1460.890 2896.760 ;
        RECT 1460.375 2896.560 1460.890 2896.700 ;
        RECT 1460.570 2896.500 1460.890 2896.560 ;
        RECT 1460.585 2895.340 1460.875 2895.385 ;
        RECT 2899.450 2895.340 2899.770 2895.400 ;
        RECT 1460.585 2895.200 2899.770 2895.340 ;
        RECT 1460.585 2895.155 1460.875 2895.200 ;
        RECT 2899.450 2895.140 2899.770 2895.200 ;
      LAYER via ;
        RECT 1460.600 2896.500 1460.860 2896.760 ;
        RECT 2899.480 2895.140 2899.740 2895.400 ;
      LAYER met2 ;
        RECT 1459.145 2896.530 1459.425 2900.000 ;
        RECT 1460.600 2896.530 1460.860 2896.790 ;
        RECT 1459.145 2896.470 1460.860 2896.530 ;
        RECT 1459.145 2896.390 1460.800 2896.470 ;
        RECT 1459.145 2896.000 1459.425 2896.390 ;
        RECT 2899.480 2895.110 2899.740 2895.430 ;
        RECT 2899.540 2258.805 2899.680 2895.110 ;
        RECT 2899.470 2258.435 2899.750 2258.805 ;
      LAYER via2 ;
        RECT 2899.470 2258.480 2899.750 2258.760 ;
      LAYER met3 ;
        RECT 2899.445 2258.770 2899.775 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2899.445 2258.470 2924.800 2258.770 ;
        RECT 2899.445 2258.455 2899.775 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 634.410 59.060 634.730 59.120 ;
        RECT 1407.670 59.060 1407.990 59.120 ;
        RECT 634.410 58.920 1407.990 59.060 ;
        RECT 634.410 58.860 634.730 58.920 ;
        RECT 1407.670 58.860 1407.990 58.920 ;
      LAYER via ;
        RECT 634.440 58.860 634.700 59.120 ;
        RECT 1407.700 58.860 1407.960 59.120 ;
      LAYER met2 ;
        RECT 1409.465 1700.410 1409.745 1704.000 ;
        RECT 1407.760 1700.270 1409.745 1700.410 ;
        RECT 1407.760 59.150 1407.900 1700.270 ;
        RECT 1409.465 1700.000 1409.745 1700.270 ;
        RECT 634.440 58.830 634.700 59.150 ;
        RECT 1407.700 58.830 1407.960 59.150 ;
        RECT 634.500 17.410 634.640 58.830 ;
        RECT 633.120 17.270 634.640 17.410 ;
        RECT 633.120 2.400 633.260 17.270 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2145.510 29.480 2145.830 29.540 ;
        RECT 2417.370 29.480 2417.690 29.540 ;
        RECT 2145.510 29.340 2417.690 29.480 ;
        RECT 2145.510 29.280 2145.830 29.340 ;
        RECT 2417.370 29.280 2417.690 29.340 ;
      LAYER via ;
        RECT 2145.540 29.280 2145.800 29.540 ;
        RECT 2417.400 29.280 2417.660 29.540 ;
      LAYER met2 ;
        RECT 2144.085 1700.410 2144.365 1704.000 ;
        RECT 2144.085 1700.270 2145.740 1700.410 ;
        RECT 2144.085 1700.000 2144.365 1700.270 ;
        RECT 2145.600 29.570 2145.740 1700.270 ;
        RECT 2145.540 29.250 2145.800 29.570 ;
        RECT 2417.400 29.250 2417.660 29.570 ;
        RECT 2417.460 2.400 2417.600 29.250 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2152.410 30.160 2152.730 30.220 ;
        RECT 2434.850 30.160 2435.170 30.220 ;
        RECT 2152.410 30.020 2435.170 30.160 ;
        RECT 2152.410 29.960 2152.730 30.020 ;
        RECT 2434.850 29.960 2435.170 30.020 ;
      LAYER via ;
        RECT 2152.440 29.960 2152.700 30.220 ;
        RECT 2434.880 29.960 2435.140 30.220 ;
      LAYER met2 ;
        RECT 2151.445 1700.410 2151.725 1704.000 ;
        RECT 2151.445 1700.270 2152.640 1700.410 ;
        RECT 2151.445 1700.000 2151.725 1700.270 ;
        RECT 2152.500 30.250 2152.640 1700.270 ;
        RECT 2152.440 29.930 2152.700 30.250 ;
        RECT 2434.880 29.930 2435.140 30.250 ;
        RECT 2434.940 2.400 2435.080 29.930 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2159.310 34.240 2159.630 34.300 ;
        RECT 2452.790 34.240 2453.110 34.300 ;
        RECT 2159.310 34.100 2453.110 34.240 ;
        RECT 2159.310 34.040 2159.630 34.100 ;
        RECT 2452.790 34.040 2453.110 34.100 ;
      LAYER via ;
        RECT 2159.340 34.040 2159.600 34.300 ;
        RECT 2452.820 34.040 2453.080 34.300 ;
      LAYER met2 ;
        RECT 2158.805 1700.410 2159.085 1704.000 ;
        RECT 2158.805 1700.270 2159.540 1700.410 ;
        RECT 2158.805 1700.000 2159.085 1700.270 ;
        RECT 2159.400 34.330 2159.540 1700.270 ;
        RECT 2159.340 34.010 2159.600 34.330 ;
        RECT 2452.820 34.010 2453.080 34.330 ;
        RECT 2452.880 2.400 2453.020 34.010 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2166.210 33.220 2166.530 33.280 ;
        RECT 2470.730 33.220 2471.050 33.280 ;
        RECT 2166.210 33.080 2471.050 33.220 ;
        RECT 2166.210 33.020 2166.530 33.080 ;
        RECT 2470.730 33.020 2471.050 33.080 ;
      LAYER via ;
        RECT 2166.240 33.020 2166.500 33.280 ;
        RECT 2470.760 33.020 2471.020 33.280 ;
      LAYER met2 ;
        RECT 2166.165 1700.000 2166.445 1704.000 ;
        RECT 2166.300 33.310 2166.440 1700.000 ;
        RECT 2166.240 32.990 2166.500 33.310 ;
        RECT 2470.760 32.990 2471.020 33.310 ;
        RECT 2470.820 2.400 2470.960 32.990 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2173.570 1684.260 2173.890 1684.320 ;
        RECT 2179.550 1684.260 2179.870 1684.320 ;
        RECT 2173.570 1684.120 2179.870 1684.260 ;
        RECT 2173.570 1684.060 2173.890 1684.120 ;
        RECT 2179.550 1684.060 2179.870 1684.120 ;
        RECT 2179.550 32.880 2179.870 32.940 ;
        RECT 2488.670 32.880 2488.990 32.940 ;
        RECT 2179.550 32.740 2488.990 32.880 ;
        RECT 2179.550 32.680 2179.870 32.740 ;
        RECT 2488.670 32.680 2488.990 32.740 ;
      LAYER via ;
        RECT 2173.600 1684.060 2173.860 1684.320 ;
        RECT 2179.580 1684.060 2179.840 1684.320 ;
        RECT 2179.580 32.680 2179.840 32.940 ;
        RECT 2488.700 32.680 2488.960 32.940 ;
      LAYER met2 ;
        RECT 2173.525 1700.000 2173.805 1704.000 ;
        RECT 2173.660 1684.350 2173.800 1700.000 ;
        RECT 2173.600 1684.030 2173.860 1684.350 ;
        RECT 2179.580 1684.030 2179.840 1684.350 ;
        RECT 2179.640 32.970 2179.780 1684.030 ;
        RECT 2179.580 32.650 2179.840 32.970 ;
        RECT 2488.700 32.650 2488.960 32.970 ;
        RECT 2488.760 2.400 2488.900 32.650 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2180.930 1683.920 2181.250 1683.980 ;
        RECT 2186.910 1683.920 2187.230 1683.980 ;
        RECT 2180.930 1683.780 2187.230 1683.920 ;
        RECT 2180.930 1683.720 2181.250 1683.780 ;
        RECT 2186.910 1683.720 2187.230 1683.780 ;
        RECT 2186.910 32.200 2187.230 32.260 ;
        RECT 2506.150 32.200 2506.470 32.260 ;
        RECT 2186.910 32.060 2506.470 32.200 ;
        RECT 2186.910 32.000 2187.230 32.060 ;
        RECT 2506.150 32.000 2506.470 32.060 ;
      LAYER via ;
        RECT 2180.960 1683.720 2181.220 1683.980 ;
        RECT 2186.940 1683.720 2187.200 1683.980 ;
        RECT 2186.940 32.000 2187.200 32.260 ;
        RECT 2506.180 32.000 2506.440 32.260 ;
      LAYER met2 ;
        RECT 2180.885 1700.000 2181.165 1704.000 ;
        RECT 2181.020 1684.010 2181.160 1700.000 ;
        RECT 2180.960 1683.690 2181.220 1684.010 ;
        RECT 2186.940 1683.690 2187.200 1684.010 ;
        RECT 2187.000 32.290 2187.140 1683.690 ;
        RECT 2186.940 31.970 2187.200 32.290 ;
        RECT 2506.180 31.970 2506.440 32.290 ;
        RECT 2506.240 2.400 2506.380 31.970 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2188.290 1688.000 2188.610 1688.060 ;
        RECT 2193.350 1688.000 2193.670 1688.060 ;
        RECT 2188.290 1687.860 2193.670 1688.000 ;
        RECT 2188.290 1687.800 2188.610 1687.860 ;
        RECT 2193.350 1687.800 2193.670 1687.860 ;
        RECT 2193.350 31.520 2193.670 31.580 ;
        RECT 2524.090 31.520 2524.410 31.580 ;
        RECT 2193.350 31.380 2524.410 31.520 ;
        RECT 2193.350 31.320 2193.670 31.380 ;
        RECT 2524.090 31.320 2524.410 31.380 ;
      LAYER via ;
        RECT 2188.320 1687.800 2188.580 1688.060 ;
        RECT 2193.380 1687.800 2193.640 1688.060 ;
        RECT 2193.380 31.320 2193.640 31.580 ;
        RECT 2524.120 31.320 2524.380 31.580 ;
      LAYER met2 ;
        RECT 2188.245 1700.000 2188.525 1704.000 ;
        RECT 2188.380 1688.090 2188.520 1700.000 ;
        RECT 2188.320 1687.770 2188.580 1688.090 ;
        RECT 2193.380 1687.770 2193.640 1688.090 ;
        RECT 2193.440 31.610 2193.580 1687.770 ;
        RECT 2193.380 31.290 2193.640 31.610 ;
        RECT 2524.120 31.290 2524.380 31.610 ;
        RECT 2524.180 2.400 2524.320 31.290 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2195.650 1688.680 2195.970 1688.740 ;
        RECT 2200.710 1688.680 2201.030 1688.740 ;
        RECT 2195.650 1688.540 2201.030 1688.680 ;
        RECT 2195.650 1688.480 2195.970 1688.540 ;
        RECT 2200.710 1688.480 2201.030 1688.540 ;
        RECT 2200.710 30.840 2201.030 30.900 ;
        RECT 2542.030 30.840 2542.350 30.900 ;
        RECT 2200.710 30.700 2542.350 30.840 ;
        RECT 2200.710 30.640 2201.030 30.700 ;
        RECT 2542.030 30.640 2542.350 30.700 ;
      LAYER via ;
        RECT 2195.680 1688.480 2195.940 1688.740 ;
        RECT 2200.740 1688.480 2201.000 1688.740 ;
        RECT 2200.740 30.640 2201.000 30.900 ;
        RECT 2542.060 30.640 2542.320 30.900 ;
      LAYER met2 ;
        RECT 2195.605 1700.000 2195.885 1704.000 ;
        RECT 2195.740 1688.770 2195.880 1700.000 ;
        RECT 2195.680 1688.450 2195.940 1688.770 ;
        RECT 2200.740 1688.450 2201.000 1688.770 ;
        RECT 2200.800 30.930 2200.940 1688.450 ;
        RECT 2200.740 30.610 2201.000 30.930 ;
        RECT 2542.060 30.610 2542.320 30.930 ;
        RECT 2542.120 2.400 2542.260 30.610 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2203.010 1688.000 2203.330 1688.060 ;
        RECT 2207.610 1688.000 2207.930 1688.060 ;
        RECT 2203.010 1687.860 2207.930 1688.000 ;
        RECT 2203.010 1687.800 2203.330 1687.860 ;
        RECT 2207.610 1687.800 2207.930 1687.860 ;
        RECT 2207.610 21.320 2207.930 21.380 ;
        RECT 2559.970 21.320 2560.290 21.380 ;
        RECT 2207.610 21.180 2560.290 21.320 ;
        RECT 2207.610 21.120 2207.930 21.180 ;
        RECT 2559.970 21.120 2560.290 21.180 ;
      LAYER via ;
        RECT 2203.040 1687.800 2203.300 1688.060 ;
        RECT 2207.640 1687.800 2207.900 1688.060 ;
        RECT 2207.640 21.120 2207.900 21.380 ;
        RECT 2560.000 21.120 2560.260 21.380 ;
      LAYER met2 ;
        RECT 2202.965 1700.000 2203.245 1704.000 ;
        RECT 2203.100 1688.090 2203.240 1700.000 ;
        RECT 2203.040 1687.770 2203.300 1688.090 ;
        RECT 2207.640 1687.770 2207.900 1688.090 ;
        RECT 2207.700 21.410 2207.840 1687.770 ;
        RECT 2207.640 21.090 2207.900 21.410 ;
        RECT 2560.000 21.090 2560.260 21.410 ;
        RECT 2560.060 2.400 2560.200 21.090 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2210.370 1688.340 2210.690 1688.400 ;
        RECT 2214.510 1688.340 2214.830 1688.400 ;
        RECT 2210.370 1688.200 2214.830 1688.340 ;
        RECT 2210.370 1688.140 2210.690 1688.200 ;
        RECT 2214.510 1688.140 2214.830 1688.200 ;
        RECT 2214.510 21.660 2214.830 21.720 ;
        RECT 2577.910 21.660 2578.230 21.720 ;
        RECT 2214.510 21.520 2578.230 21.660 ;
        RECT 2214.510 21.460 2214.830 21.520 ;
        RECT 2577.910 21.460 2578.230 21.520 ;
      LAYER via ;
        RECT 2210.400 1688.140 2210.660 1688.400 ;
        RECT 2214.540 1688.140 2214.800 1688.400 ;
        RECT 2214.540 21.460 2214.800 21.720 ;
        RECT 2577.940 21.460 2578.200 21.720 ;
      LAYER met2 ;
        RECT 2210.325 1700.000 2210.605 1704.000 ;
        RECT 2210.460 1688.430 2210.600 1700.000 ;
        RECT 2210.400 1688.110 2210.660 1688.430 ;
        RECT 2214.540 1688.110 2214.800 1688.430 ;
        RECT 2214.600 21.750 2214.740 1688.110 ;
        RECT 2214.540 21.430 2214.800 21.750 ;
        RECT 2577.940 21.430 2578.200 21.750 ;
        RECT 2578.000 2.400 2578.140 21.430 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1478.585 582.845 1478.755 613.955 ;
        RECT 1478.585 510.765 1478.755 558.875 ;
        RECT 1477.665 241.485 1477.835 307.275 ;
        RECT 1477.665 60.945 1477.835 96.475 ;
      LAYER mcon ;
        RECT 1478.585 613.785 1478.755 613.955 ;
        RECT 1478.585 558.705 1478.755 558.875 ;
        RECT 1477.665 307.105 1477.835 307.275 ;
        RECT 1477.665 96.305 1477.835 96.475 ;
      LAYER met1 ;
        RECT 1477.590 1642.100 1477.910 1642.160 ;
        RECT 1478.510 1642.100 1478.830 1642.160 ;
        RECT 1477.590 1641.960 1478.830 1642.100 ;
        RECT 1477.590 1641.900 1477.910 1641.960 ;
        RECT 1478.510 1641.900 1478.830 1641.960 ;
        RECT 1477.590 1521.400 1477.910 1521.460 ;
        RECT 1478.510 1521.400 1478.830 1521.460 ;
        RECT 1477.590 1521.260 1478.830 1521.400 ;
        RECT 1477.590 1521.200 1477.910 1521.260 ;
        RECT 1478.510 1521.200 1478.830 1521.260 ;
        RECT 1477.590 1462.720 1477.910 1462.980 ;
        RECT 1477.680 1462.580 1477.820 1462.720 ;
        RECT 1478.050 1462.580 1478.370 1462.640 ;
        RECT 1477.680 1462.440 1478.370 1462.580 ;
        RECT 1478.050 1462.380 1478.370 1462.440 ;
        RECT 1478.050 1414.980 1478.370 1415.040 ;
        RECT 1477.680 1414.840 1478.370 1414.980 ;
        RECT 1477.680 1414.360 1477.820 1414.840 ;
        RECT 1478.050 1414.780 1478.370 1414.840 ;
        RECT 1477.590 1414.100 1477.910 1414.360 ;
        RECT 1477.590 1345.620 1477.910 1345.680 ;
        RECT 1478.970 1345.620 1479.290 1345.680 ;
        RECT 1477.590 1345.480 1479.290 1345.620 ;
        RECT 1477.590 1345.420 1477.910 1345.480 ;
        RECT 1478.970 1345.420 1479.290 1345.480 ;
        RECT 1477.590 1290.200 1477.910 1290.260 ;
        RECT 1478.510 1290.200 1478.830 1290.260 ;
        RECT 1477.590 1290.060 1478.830 1290.200 ;
        RECT 1477.590 1290.000 1477.910 1290.060 ;
        RECT 1478.510 1290.000 1478.830 1290.060 ;
        RECT 1477.590 1111.020 1477.910 1111.080 ;
        RECT 1478.050 1111.020 1478.370 1111.080 ;
        RECT 1477.590 1110.880 1478.370 1111.020 ;
        RECT 1477.590 1110.820 1477.910 1110.880 ;
        RECT 1478.050 1110.820 1478.370 1110.880 ;
        RECT 1477.590 1014.460 1477.910 1014.520 ;
        RECT 1478.050 1014.460 1478.370 1014.520 ;
        RECT 1477.590 1014.320 1478.370 1014.460 ;
        RECT 1477.590 1014.260 1477.910 1014.320 ;
        RECT 1478.050 1014.260 1478.370 1014.320 ;
        RECT 1478.050 931.840 1478.370 931.900 ;
        RECT 1477.680 931.700 1478.370 931.840 ;
        RECT 1477.680 931.560 1477.820 931.700 ;
        RECT 1478.050 931.640 1478.370 931.700 ;
        RECT 1477.590 931.300 1477.910 931.560 ;
        RECT 1477.590 893.760 1477.910 893.820 ;
        RECT 1478.510 893.760 1478.830 893.820 ;
        RECT 1477.590 893.620 1478.830 893.760 ;
        RECT 1477.590 893.560 1477.910 893.620 ;
        RECT 1478.510 893.560 1478.830 893.620 ;
        RECT 1478.050 807.400 1478.370 807.460 ;
        RECT 1478.510 807.400 1478.830 807.460 ;
        RECT 1478.050 807.260 1478.830 807.400 ;
        RECT 1478.050 807.200 1478.370 807.260 ;
        RECT 1478.510 807.200 1478.830 807.260 ;
        RECT 1477.590 662.560 1477.910 662.620 ;
        RECT 1478.050 662.560 1478.370 662.620 ;
        RECT 1477.590 662.420 1478.370 662.560 ;
        RECT 1477.590 662.360 1477.910 662.420 ;
        RECT 1478.050 662.360 1478.370 662.420 ;
        RECT 1478.510 613.940 1478.830 614.000 ;
        RECT 1478.315 613.800 1478.830 613.940 ;
        RECT 1478.510 613.740 1478.830 613.800 ;
        RECT 1478.525 583.000 1478.815 583.045 ;
        RECT 1478.970 583.000 1479.290 583.060 ;
        RECT 1478.525 582.860 1479.290 583.000 ;
        RECT 1478.525 582.815 1478.815 582.860 ;
        RECT 1478.970 582.800 1479.290 582.860 ;
        RECT 1478.510 558.860 1478.830 558.920 ;
        RECT 1478.315 558.720 1478.830 558.860 ;
        RECT 1478.510 558.660 1478.830 558.720 ;
        RECT 1478.525 510.920 1478.815 510.965 ;
        RECT 1479.430 510.920 1479.750 510.980 ;
        RECT 1478.525 510.780 1479.750 510.920 ;
        RECT 1478.525 510.735 1478.815 510.780 ;
        RECT 1479.430 510.720 1479.750 510.780 ;
        RECT 1478.510 414.360 1478.830 414.420 ;
        RECT 1479.430 414.360 1479.750 414.420 ;
        RECT 1478.510 414.220 1479.750 414.360 ;
        RECT 1478.510 414.160 1478.830 414.220 ;
        RECT 1479.430 414.160 1479.750 414.220 ;
        RECT 1478.050 324.600 1478.370 324.660 ;
        RECT 1478.510 324.600 1478.830 324.660 ;
        RECT 1478.050 324.460 1478.830 324.600 ;
        RECT 1478.050 324.400 1478.370 324.460 ;
        RECT 1478.510 324.400 1478.830 324.460 ;
        RECT 1477.605 307.260 1477.895 307.305 ;
        RECT 1478.050 307.260 1478.370 307.320 ;
        RECT 1477.605 307.120 1478.370 307.260 ;
        RECT 1477.605 307.075 1477.895 307.120 ;
        RECT 1478.050 307.060 1478.370 307.120 ;
        RECT 1477.590 241.640 1477.910 241.700 ;
        RECT 1477.395 241.500 1477.910 241.640 ;
        RECT 1477.590 241.440 1477.910 241.500 ;
        RECT 1478.050 138.620 1478.370 138.680 ;
        RECT 1477.680 138.480 1478.370 138.620 ;
        RECT 1477.680 138.340 1477.820 138.480 ;
        RECT 1478.050 138.420 1478.370 138.480 ;
        RECT 1477.590 138.080 1477.910 138.340 ;
        RECT 1477.590 96.460 1477.910 96.520 ;
        RECT 1477.395 96.320 1477.910 96.460 ;
        RECT 1477.590 96.260 1477.910 96.320 ;
        RECT 813.810 61.100 814.130 61.160 ;
        RECT 1477.605 61.100 1477.895 61.145 ;
        RECT 813.810 60.960 1477.895 61.100 ;
        RECT 813.810 60.900 814.130 60.960 ;
        RECT 1477.605 60.915 1477.895 60.960 ;
      LAYER via ;
        RECT 1477.620 1641.900 1477.880 1642.160 ;
        RECT 1478.540 1641.900 1478.800 1642.160 ;
        RECT 1477.620 1521.200 1477.880 1521.460 ;
        RECT 1478.540 1521.200 1478.800 1521.460 ;
        RECT 1477.620 1462.720 1477.880 1462.980 ;
        RECT 1478.080 1462.380 1478.340 1462.640 ;
        RECT 1478.080 1414.780 1478.340 1415.040 ;
        RECT 1477.620 1414.100 1477.880 1414.360 ;
        RECT 1477.620 1345.420 1477.880 1345.680 ;
        RECT 1479.000 1345.420 1479.260 1345.680 ;
        RECT 1477.620 1290.000 1477.880 1290.260 ;
        RECT 1478.540 1290.000 1478.800 1290.260 ;
        RECT 1477.620 1110.820 1477.880 1111.080 ;
        RECT 1478.080 1110.820 1478.340 1111.080 ;
        RECT 1477.620 1014.260 1477.880 1014.520 ;
        RECT 1478.080 1014.260 1478.340 1014.520 ;
        RECT 1478.080 931.640 1478.340 931.900 ;
        RECT 1477.620 931.300 1477.880 931.560 ;
        RECT 1477.620 893.560 1477.880 893.820 ;
        RECT 1478.540 893.560 1478.800 893.820 ;
        RECT 1478.080 807.200 1478.340 807.460 ;
        RECT 1478.540 807.200 1478.800 807.460 ;
        RECT 1477.620 662.360 1477.880 662.620 ;
        RECT 1478.080 662.360 1478.340 662.620 ;
        RECT 1478.540 613.740 1478.800 614.000 ;
        RECT 1479.000 582.800 1479.260 583.060 ;
        RECT 1478.540 558.660 1478.800 558.920 ;
        RECT 1479.460 510.720 1479.720 510.980 ;
        RECT 1478.540 414.160 1478.800 414.420 ;
        RECT 1479.460 414.160 1479.720 414.420 ;
        RECT 1478.080 324.400 1478.340 324.660 ;
        RECT 1478.540 324.400 1478.800 324.660 ;
        RECT 1478.080 307.060 1478.340 307.320 ;
        RECT 1477.620 241.440 1477.880 241.700 ;
        RECT 1478.080 138.420 1478.340 138.680 ;
        RECT 1477.620 138.080 1477.880 138.340 ;
        RECT 1477.620 96.260 1477.880 96.520 ;
        RECT 813.840 60.900 814.100 61.160 ;
      LAYER met2 ;
        RECT 1483.065 1700.410 1483.345 1704.000 ;
        RECT 1481.360 1700.270 1483.345 1700.410 ;
        RECT 1481.360 1677.970 1481.500 1700.270 ;
        RECT 1483.065 1700.000 1483.345 1700.270 ;
        RECT 1477.680 1677.830 1481.500 1677.970 ;
        RECT 1477.680 1642.190 1477.820 1677.830 ;
        RECT 1477.620 1641.870 1477.880 1642.190 ;
        RECT 1478.540 1641.870 1478.800 1642.190 ;
        RECT 1478.600 1617.450 1478.740 1641.870 ;
        RECT 1478.140 1617.310 1478.740 1617.450 ;
        RECT 1478.140 1563.050 1478.280 1617.310 ;
        RECT 1478.140 1562.910 1478.740 1563.050 ;
        RECT 1478.600 1521.490 1478.740 1562.910 ;
        RECT 1477.620 1521.170 1477.880 1521.490 ;
        RECT 1478.540 1521.170 1478.800 1521.490 ;
        RECT 1477.680 1463.010 1477.820 1521.170 ;
        RECT 1477.620 1462.690 1477.880 1463.010 ;
        RECT 1478.080 1462.350 1478.340 1462.670 ;
        RECT 1478.140 1415.070 1478.280 1462.350 ;
        RECT 1478.080 1414.750 1478.340 1415.070 ;
        RECT 1477.620 1414.070 1477.880 1414.390 ;
        RECT 1477.680 1345.710 1477.820 1414.070 ;
        RECT 1477.620 1345.390 1477.880 1345.710 ;
        RECT 1479.000 1345.390 1479.260 1345.710 ;
        RECT 1479.060 1304.650 1479.200 1345.390 ;
        RECT 1479.060 1304.510 1479.660 1304.650 ;
        RECT 1479.520 1290.485 1479.660 1304.510 ;
        RECT 1477.620 1289.970 1477.880 1290.290 ;
        RECT 1478.530 1290.115 1478.810 1290.485 ;
        RECT 1479.450 1290.115 1479.730 1290.485 ;
        RECT 1478.540 1289.970 1478.800 1290.115 ;
        RECT 1477.680 1207.410 1477.820 1289.970 ;
        RECT 1477.680 1207.270 1478.280 1207.410 ;
        RECT 1477.680 1111.110 1477.820 1111.265 ;
        RECT 1478.140 1111.110 1478.280 1207.270 ;
        RECT 1477.620 1110.850 1477.880 1111.110 ;
        RECT 1478.080 1110.850 1478.340 1111.110 ;
        RECT 1477.620 1110.790 1478.340 1110.850 ;
        RECT 1477.680 1110.710 1478.280 1110.790 ;
        RECT 1477.680 1014.550 1477.820 1014.705 ;
        RECT 1478.140 1014.550 1478.280 1110.710 ;
        RECT 1477.620 1014.290 1477.880 1014.550 ;
        RECT 1478.080 1014.290 1478.340 1014.550 ;
        RECT 1477.620 1014.230 1478.340 1014.290 ;
        RECT 1477.680 1014.150 1478.280 1014.230 ;
        RECT 1478.140 931.930 1478.280 1014.150 ;
        RECT 1478.080 931.610 1478.340 931.930 ;
        RECT 1477.620 931.270 1477.880 931.590 ;
        RECT 1477.680 893.850 1477.820 931.270 ;
        RECT 1477.620 893.530 1477.880 893.850 ;
        RECT 1478.540 893.530 1478.800 893.850 ;
        RECT 1478.600 807.490 1478.740 893.530 ;
        RECT 1478.080 807.170 1478.340 807.490 ;
        RECT 1478.540 807.170 1478.800 807.490 ;
        RECT 1478.140 717.810 1478.280 807.170 ;
        RECT 1477.680 717.670 1478.280 717.810 ;
        RECT 1477.680 662.650 1477.820 717.670 ;
        RECT 1477.620 662.330 1477.880 662.650 ;
        RECT 1478.080 662.330 1478.340 662.650 ;
        RECT 1478.140 662.050 1478.280 662.330 ;
        RECT 1477.680 661.910 1478.280 662.050 ;
        RECT 1477.680 620.570 1477.820 661.910 ;
        RECT 1477.680 620.430 1478.740 620.570 ;
        RECT 1478.600 614.030 1478.740 620.430 ;
        RECT 1478.540 613.710 1478.800 614.030 ;
        RECT 1479.000 582.770 1479.260 583.090 ;
        RECT 1479.060 559.370 1479.200 582.770 ;
        RECT 1478.600 559.230 1479.200 559.370 ;
        RECT 1478.600 558.950 1478.740 559.230 ;
        RECT 1478.540 558.630 1478.800 558.950 ;
        RECT 1479.460 510.690 1479.720 511.010 ;
        RECT 1479.520 414.450 1479.660 510.690 ;
        RECT 1478.540 414.130 1478.800 414.450 ;
        RECT 1479.460 414.130 1479.720 414.450 ;
        RECT 1478.600 324.690 1478.740 414.130 ;
        RECT 1478.080 324.370 1478.340 324.690 ;
        RECT 1478.540 324.370 1478.800 324.690 ;
        RECT 1478.140 307.350 1478.280 324.370 ;
        RECT 1478.080 307.030 1478.340 307.350 ;
        RECT 1477.620 241.410 1477.880 241.730 ;
        RECT 1477.680 192.170 1477.820 241.410 ;
        RECT 1477.680 192.030 1478.280 192.170 ;
        RECT 1478.140 138.710 1478.280 192.030 ;
        RECT 1478.080 138.390 1478.340 138.710 ;
        RECT 1477.620 138.050 1477.880 138.370 ;
        RECT 1477.680 96.550 1477.820 138.050 ;
        RECT 1477.620 96.230 1477.880 96.550 ;
        RECT 813.840 60.870 814.100 61.190 ;
        RECT 813.900 3.130 814.040 60.870 ;
        RECT 811.600 2.990 814.040 3.130 ;
        RECT 811.600 2.400 811.740 2.990 ;
        RECT 811.390 -4.800 811.950 2.400 ;
      LAYER via2 ;
        RECT 1478.530 1290.160 1478.810 1290.440 ;
        RECT 1479.450 1290.160 1479.730 1290.440 ;
      LAYER met3 ;
        RECT 1478.505 1290.450 1478.835 1290.465 ;
        RECT 1479.425 1290.450 1479.755 1290.465 ;
        RECT 1478.505 1290.150 1479.755 1290.450 ;
        RECT 1478.505 1290.135 1478.835 1290.150 ;
        RECT 1479.425 1290.135 1479.755 1290.150 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2217.730 1688.340 2218.050 1688.400 ;
        RECT 2221.410 1688.340 2221.730 1688.400 ;
        RECT 2217.730 1688.200 2221.730 1688.340 ;
        RECT 2217.730 1688.140 2218.050 1688.200 ;
        RECT 2221.410 1688.140 2221.730 1688.200 ;
        RECT 2221.410 22.000 2221.730 22.060 ;
        RECT 2595.390 22.000 2595.710 22.060 ;
        RECT 2221.410 21.860 2595.710 22.000 ;
        RECT 2221.410 21.800 2221.730 21.860 ;
        RECT 2595.390 21.800 2595.710 21.860 ;
      LAYER via ;
        RECT 2217.760 1688.140 2218.020 1688.400 ;
        RECT 2221.440 1688.140 2221.700 1688.400 ;
        RECT 2221.440 21.800 2221.700 22.060 ;
        RECT 2595.420 21.800 2595.680 22.060 ;
      LAYER met2 ;
        RECT 2217.685 1700.000 2217.965 1704.000 ;
        RECT 2217.820 1688.430 2217.960 1700.000 ;
        RECT 2217.760 1688.110 2218.020 1688.430 ;
        RECT 2221.440 1688.110 2221.700 1688.430 ;
        RECT 2221.500 22.090 2221.640 1688.110 ;
        RECT 2221.440 21.770 2221.700 22.090 ;
        RECT 2595.420 21.770 2595.680 22.090 ;
        RECT 2595.480 2.400 2595.620 21.770 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2225.090 1688.340 2225.410 1688.400 ;
        RECT 2227.850 1688.340 2228.170 1688.400 ;
        RECT 2225.090 1688.200 2228.170 1688.340 ;
        RECT 2225.090 1688.140 2225.410 1688.200 ;
        RECT 2227.850 1688.140 2228.170 1688.200 ;
        RECT 2227.850 22.340 2228.170 22.400 ;
        RECT 2613.330 22.340 2613.650 22.400 ;
        RECT 2227.850 22.200 2613.650 22.340 ;
        RECT 2227.850 22.140 2228.170 22.200 ;
        RECT 2613.330 22.140 2613.650 22.200 ;
      LAYER via ;
        RECT 2225.120 1688.140 2225.380 1688.400 ;
        RECT 2227.880 1688.140 2228.140 1688.400 ;
        RECT 2227.880 22.140 2228.140 22.400 ;
        RECT 2613.360 22.140 2613.620 22.400 ;
      LAYER met2 ;
        RECT 2225.045 1700.000 2225.325 1704.000 ;
        RECT 2225.180 1688.430 2225.320 1700.000 ;
        RECT 2225.120 1688.110 2225.380 1688.430 ;
        RECT 2227.880 1688.110 2228.140 1688.430 ;
        RECT 2227.940 22.430 2228.080 1688.110 ;
        RECT 2227.880 22.110 2228.140 22.430 ;
        RECT 2613.360 22.110 2613.620 22.430 ;
        RECT 2613.420 2.400 2613.560 22.110 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2232.450 1688.340 2232.770 1688.400 ;
        RECT 2235.210 1688.340 2235.530 1688.400 ;
        RECT 2232.450 1688.200 2235.530 1688.340 ;
        RECT 2232.450 1688.140 2232.770 1688.200 ;
        RECT 2235.210 1688.140 2235.530 1688.200 ;
        RECT 2235.210 22.680 2235.530 22.740 ;
        RECT 2631.270 22.680 2631.590 22.740 ;
        RECT 2235.210 22.540 2631.590 22.680 ;
        RECT 2235.210 22.480 2235.530 22.540 ;
        RECT 2631.270 22.480 2631.590 22.540 ;
      LAYER via ;
        RECT 2232.480 1688.140 2232.740 1688.400 ;
        RECT 2235.240 1688.140 2235.500 1688.400 ;
        RECT 2235.240 22.480 2235.500 22.740 ;
        RECT 2631.300 22.480 2631.560 22.740 ;
      LAYER met2 ;
        RECT 2232.405 1700.000 2232.685 1704.000 ;
        RECT 2232.540 1688.430 2232.680 1700.000 ;
        RECT 2232.480 1688.110 2232.740 1688.430 ;
        RECT 2235.240 1688.110 2235.500 1688.430 ;
        RECT 2235.300 22.770 2235.440 1688.110 ;
        RECT 2235.240 22.450 2235.500 22.770 ;
        RECT 2631.300 22.450 2631.560 22.770 ;
        RECT 2631.360 2.400 2631.500 22.450 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2241.650 23.020 2241.970 23.080 ;
        RECT 2649.210 23.020 2649.530 23.080 ;
        RECT 2241.650 22.880 2649.530 23.020 ;
        RECT 2241.650 22.820 2241.970 22.880 ;
        RECT 2649.210 22.820 2649.530 22.880 ;
      LAYER via ;
        RECT 2241.680 22.820 2241.940 23.080 ;
        RECT 2649.240 22.820 2649.500 23.080 ;
      LAYER met2 ;
        RECT 2239.765 1700.410 2240.045 1704.000 ;
        RECT 2239.765 1700.270 2241.880 1700.410 ;
        RECT 2239.765 1700.000 2240.045 1700.270 ;
        RECT 2241.740 23.110 2241.880 1700.270 ;
        RECT 2241.680 22.790 2241.940 23.110 ;
        RECT 2649.240 22.790 2649.500 23.110 ;
        RECT 2649.300 2.400 2649.440 22.790 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2249.010 23.360 2249.330 23.420 ;
        RECT 2667.150 23.360 2667.470 23.420 ;
        RECT 2249.010 23.220 2667.470 23.360 ;
        RECT 2249.010 23.160 2249.330 23.220 ;
        RECT 2667.150 23.160 2667.470 23.220 ;
      LAYER via ;
        RECT 2249.040 23.160 2249.300 23.420 ;
        RECT 2667.180 23.160 2667.440 23.420 ;
      LAYER met2 ;
        RECT 2247.125 1700.410 2247.405 1704.000 ;
        RECT 2247.125 1700.270 2249.240 1700.410 ;
        RECT 2247.125 1700.000 2247.405 1700.270 ;
        RECT 2249.100 23.450 2249.240 1700.270 ;
        RECT 2249.040 23.130 2249.300 23.450 ;
        RECT 2667.180 23.130 2667.440 23.450 ;
        RECT 2667.240 2.400 2667.380 23.130 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2255.450 23.700 2255.770 23.760 ;
        RECT 2684.630 23.700 2684.950 23.760 ;
        RECT 2255.450 23.560 2684.950 23.700 ;
        RECT 2255.450 23.500 2255.770 23.560 ;
        RECT 2684.630 23.500 2684.950 23.560 ;
      LAYER via ;
        RECT 2255.480 23.500 2255.740 23.760 ;
        RECT 2684.660 23.500 2684.920 23.760 ;
      LAYER met2 ;
        RECT 2254.485 1700.410 2254.765 1704.000 ;
        RECT 2254.485 1700.270 2255.680 1700.410 ;
        RECT 2254.485 1700.000 2254.765 1700.270 ;
        RECT 2255.540 23.790 2255.680 1700.270 ;
        RECT 2255.480 23.470 2255.740 23.790 ;
        RECT 2684.660 23.470 2684.920 23.790 ;
        RECT 2684.720 2.400 2684.860 23.470 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2262.810 27.440 2263.130 27.500 ;
        RECT 2702.570 27.440 2702.890 27.500 ;
        RECT 2262.810 27.300 2702.890 27.440 ;
        RECT 2262.810 27.240 2263.130 27.300 ;
        RECT 2702.570 27.240 2702.890 27.300 ;
      LAYER via ;
        RECT 2262.840 27.240 2263.100 27.500 ;
        RECT 2702.600 27.240 2702.860 27.500 ;
      LAYER met2 ;
        RECT 2261.845 1700.410 2262.125 1704.000 ;
        RECT 2261.845 1700.270 2263.040 1700.410 ;
        RECT 2261.845 1700.000 2262.125 1700.270 ;
        RECT 2262.900 27.530 2263.040 1700.270 ;
        RECT 2262.840 27.210 2263.100 27.530 ;
        RECT 2702.600 27.210 2702.860 27.530 ;
        RECT 2702.660 2.400 2702.800 27.210 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2269.250 27.100 2269.570 27.160 ;
        RECT 2720.510 27.100 2720.830 27.160 ;
        RECT 2269.250 26.960 2720.830 27.100 ;
        RECT 2269.250 26.900 2269.570 26.960 ;
        RECT 2720.510 26.900 2720.830 26.960 ;
      LAYER via ;
        RECT 2269.280 26.900 2269.540 27.160 ;
        RECT 2720.540 26.900 2720.800 27.160 ;
      LAYER met2 ;
        RECT 2269.205 1700.000 2269.485 1704.000 ;
        RECT 2269.340 27.190 2269.480 1700.000 ;
        RECT 2269.280 26.870 2269.540 27.190 ;
        RECT 2720.540 26.870 2720.800 27.190 ;
        RECT 2720.600 2.400 2720.740 26.870 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2276.610 26.760 2276.930 26.820 ;
        RECT 2738.450 26.760 2738.770 26.820 ;
        RECT 2276.610 26.620 2738.770 26.760 ;
        RECT 2276.610 26.560 2276.930 26.620 ;
        RECT 2738.450 26.560 2738.770 26.620 ;
      LAYER via ;
        RECT 2276.640 26.560 2276.900 26.820 ;
        RECT 2738.480 26.560 2738.740 26.820 ;
      LAYER met2 ;
        RECT 2276.565 1700.000 2276.845 1704.000 ;
        RECT 2276.700 26.850 2276.840 1700.000 ;
        RECT 2276.640 26.530 2276.900 26.850 ;
        RECT 2738.480 26.530 2738.740 26.850 ;
        RECT 2738.540 2.400 2738.680 26.530 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2330.505 24.565 2330.675 26.435 ;
      LAYER mcon ;
        RECT 2330.505 26.265 2330.675 26.435 ;
      LAYER met1 ;
        RECT 2283.970 1688.340 2284.290 1688.400 ;
        RECT 2290.410 1688.340 2290.730 1688.400 ;
        RECT 2283.970 1688.200 2290.730 1688.340 ;
        RECT 2283.970 1688.140 2284.290 1688.200 ;
        RECT 2290.410 1688.140 2290.730 1688.200 ;
        RECT 2330.445 26.420 2330.735 26.465 ;
        RECT 2755.930 26.420 2756.250 26.480 ;
        RECT 2330.445 26.280 2756.250 26.420 ;
        RECT 2330.445 26.235 2330.735 26.280 ;
        RECT 2755.930 26.220 2756.250 26.280 ;
        RECT 2290.410 24.720 2290.730 24.780 ;
        RECT 2330.445 24.720 2330.735 24.765 ;
        RECT 2290.410 24.580 2330.735 24.720 ;
        RECT 2290.410 24.520 2290.730 24.580 ;
        RECT 2330.445 24.535 2330.735 24.580 ;
      LAYER via ;
        RECT 2284.000 1688.140 2284.260 1688.400 ;
        RECT 2290.440 1688.140 2290.700 1688.400 ;
        RECT 2755.960 26.220 2756.220 26.480 ;
        RECT 2290.440 24.520 2290.700 24.780 ;
      LAYER met2 ;
        RECT 2283.925 1700.000 2284.205 1704.000 ;
        RECT 2284.060 1688.430 2284.200 1700.000 ;
        RECT 2284.000 1688.110 2284.260 1688.430 ;
        RECT 2290.440 1688.110 2290.700 1688.430 ;
        RECT 2290.500 24.810 2290.640 1688.110 ;
        RECT 2755.960 26.190 2756.220 26.510 ;
        RECT 2290.440 24.490 2290.700 24.810 ;
        RECT 2756.020 2.400 2756.160 26.190 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 834.510 61.440 834.830 61.500 ;
        RECT 1490.930 61.440 1491.250 61.500 ;
        RECT 834.510 61.300 1491.250 61.440 ;
        RECT 834.510 61.240 834.830 61.300 ;
        RECT 1490.930 61.240 1491.250 61.300 ;
        RECT 829.450 2.960 829.770 3.020 ;
        RECT 834.510 2.960 834.830 3.020 ;
        RECT 829.450 2.820 834.830 2.960 ;
        RECT 829.450 2.760 829.770 2.820 ;
        RECT 834.510 2.760 834.830 2.820 ;
      LAYER via ;
        RECT 834.540 61.240 834.800 61.500 ;
        RECT 1490.960 61.240 1491.220 61.500 ;
        RECT 829.480 2.760 829.740 3.020 ;
        RECT 834.540 2.760 834.800 3.020 ;
      LAYER met2 ;
        RECT 1490.425 1700.410 1490.705 1704.000 ;
        RECT 1490.425 1700.270 1491.160 1700.410 ;
        RECT 1490.425 1700.000 1490.705 1700.270 ;
        RECT 1491.020 61.530 1491.160 1700.270 ;
        RECT 834.540 61.210 834.800 61.530 ;
        RECT 1490.960 61.210 1491.220 61.530 ;
        RECT 834.600 3.050 834.740 61.210 ;
        RECT 829.480 2.730 829.740 3.050 ;
        RECT 834.540 2.730 834.800 3.050 ;
        RECT 829.540 2.400 829.680 2.730 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2291.330 1683.920 2291.650 1683.980 ;
        RECT 2297.310 1683.920 2297.630 1683.980 ;
        RECT 2291.330 1683.780 2297.630 1683.920 ;
        RECT 2291.330 1683.720 2291.650 1683.780 ;
        RECT 2297.310 1683.720 2297.630 1683.780 ;
        RECT 2297.310 26.420 2297.630 26.480 ;
        RECT 2297.310 26.280 2330.200 26.420 ;
        RECT 2297.310 26.220 2297.630 26.280 ;
        RECT 2330.060 26.080 2330.200 26.280 ;
        RECT 2773.870 26.080 2774.190 26.140 ;
        RECT 2330.060 25.940 2774.190 26.080 ;
        RECT 2773.870 25.880 2774.190 25.940 ;
      LAYER via ;
        RECT 2291.360 1683.720 2291.620 1683.980 ;
        RECT 2297.340 1683.720 2297.600 1683.980 ;
        RECT 2297.340 26.220 2297.600 26.480 ;
        RECT 2773.900 25.880 2774.160 26.140 ;
      LAYER met2 ;
        RECT 2291.285 1700.000 2291.565 1704.000 ;
        RECT 2291.420 1684.010 2291.560 1700.000 ;
        RECT 2291.360 1683.690 2291.620 1684.010 ;
        RECT 2297.340 1683.690 2297.600 1684.010 ;
        RECT 2297.400 26.510 2297.540 1683.690 ;
        RECT 2297.340 26.190 2297.600 26.510 ;
        RECT 2773.900 25.850 2774.160 26.170 ;
        RECT 2773.960 2.400 2774.100 25.850 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2298.690 1683.920 2299.010 1683.980 ;
        RECT 2304.210 1683.920 2304.530 1683.980 ;
        RECT 2298.690 1683.780 2304.530 1683.920 ;
        RECT 2298.690 1683.720 2299.010 1683.780 ;
        RECT 2304.210 1683.720 2304.530 1683.780 ;
        RECT 2304.210 26.080 2304.530 26.140 ;
        RECT 2304.210 25.940 2329.740 26.080 ;
        RECT 2304.210 25.880 2304.530 25.940 ;
        RECT 2329.600 25.740 2329.740 25.940 ;
        RECT 2791.810 25.740 2792.130 25.800 ;
        RECT 2329.600 25.600 2792.130 25.740 ;
        RECT 2791.810 25.540 2792.130 25.600 ;
      LAYER via ;
        RECT 2298.720 1683.720 2298.980 1683.980 ;
        RECT 2304.240 1683.720 2304.500 1683.980 ;
        RECT 2304.240 25.880 2304.500 26.140 ;
        RECT 2791.840 25.540 2792.100 25.800 ;
      LAYER met2 ;
        RECT 2298.645 1700.000 2298.925 1704.000 ;
        RECT 2298.780 1684.010 2298.920 1700.000 ;
        RECT 2298.720 1683.690 2298.980 1684.010 ;
        RECT 2304.240 1683.690 2304.500 1684.010 ;
        RECT 2304.300 26.170 2304.440 1683.690 ;
        RECT 2304.240 25.850 2304.500 26.170 ;
        RECT 2791.840 25.510 2792.100 25.830 ;
        RECT 2791.900 2.400 2792.040 25.510 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2344.305 25.245 2347.695 25.415 ;
        RECT 2344.305 23.885 2344.475 25.245 ;
      LAYER mcon ;
        RECT 2347.525 25.245 2347.695 25.415 ;
      LAYER met1 ;
        RECT 2306.050 1683.920 2306.370 1683.980 ;
        RECT 2310.650 1683.920 2310.970 1683.980 ;
        RECT 2306.050 1683.780 2310.970 1683.920 ;
        RECT 2306.050 1683.720 2306.370 1683.780 ;
        RECT 2310.650 1683.720 2310.970 1683.780 ;
        RECT 2347.465 25.400 2347.755 25.445 ;
        RECT 2809.750 25.400 2810.070 25.460 ;
        RECT 2347.465 25.260 2810.070 25.400 ;
        RECT 2347.465 25.215 2347.755 25.260 ;
        RECT 2809.750 25.200 2810.070 25.260 ;
        RECT 2310.650 24.040 2310.970 24.100 ;
        RECT 2344.245 24.040 2344.535 24.085 ;
        RECT 2310.650 23.900 2344.535 24.040 ;
        RECT 2310.650 23.840 2310.970 23.900 ;
        RECT 2344.245 23.855 2344.535 23.900 ;
      LAYER via ;
        RECT 2306.080 1683.720 2306.340 1683.980 ;
        RECT 2310.680 1683.720 2310.940 1683.980 ;
        RECT 2809.780 25.200 2810.040 25.460 ;
        RECT 2310.680 23.840 2310.940 24.100 ;
      LAYER met2 ;
        RECT 2306.005 1700.000 2306.285 1704.000 ;
        RECT 2306.140 1684.010 2306.280 1700.000 ;
        RECT 2306.080 1683.690 2306.340 1684.010 ;
        RECT 2310.680 1683.690 2310.940 1684.010 ;
        RECT 2310.740 24.130 2310.880 1683.690 ;
        RECT 2809.780 25.170 2810.040 25.490 ;
        RECT 2310.680 23.810 2310.940 24.130 ;
        RECT 2809.840 2.400 2809.980 25.170 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2313.410 1683.920 2313.730 1683.980 ;
        RECT 2317.550 1683.920 2317.870 1683.980 ;
        RECT 2313.410 1683.780 2317.870 1683.920 ;
        RECT 2313.410 1683.720 2313.730 1683.780 ;
        RECT 2317.550 1683.720 2317.870 1683.780 ;
        RECT 2317.550 25.740 2317.870 25.800 ;
        RECT 2317.550 25.600 2329.280 25.740 ;
        RECT 2317.550 25.540 2317.870 25.600 ;
        RECT 2329.140 25.400 2329.280 25.600 ;
        RECT 2329.140 25.260 2347.220 25.400 ;
        RECT 2347.080 25.060 2347.220 25.260 ;
        RECT 2827.690 25.060 2828.010 25.120 ;
        RECT 2347.080 24.920 2828.010 25.060 ;
        RECT 2827.690 24.860 2828.010 24.920 ;
      LAYER via ;
        RECT 2313.440 1683.720 2313.700 1683.980 ;
        RECT 2317.580 1683.720 2317.840 1683.980 ;
        RECT 2317.580 25.540 2317.840 25.800 ;
        RECT 2827.720 24.860 2827.980 25.120 ;
      LAYER met2 ;
        RECT 2313.365 1700.000 2313.645 1704.000 ;
        RECT 2313.500 1684.010 2313.640 1700.000 ;
        RECT 2313.440 1683.690 2313.700 1684.010 ;
        RECT 2317.580 1683.690 2317.840 1684.010 ;
        RECT 2317.640 25.830 2317.780 1683.690 ;
        RECT 2317.580 25.510 2317.840 25.830 ;
        RECT 2827.720 24.830 2827.980 25.150 ;
        RECT 2827.780 2.400 2827.920 24.830 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2320.770 1683.920 2321.090 1683.980 ;
        RECT 2324.910 1683.920 2325.230 1683.980 ;
        RECT 2320.770 1683.780 2325.230 1683.920 ;
        RECT 2320.770 1683.720 2321.090 1683.780 ;
        RECT 2324.910 1683.720 2325.230 1683.780 ;
        RECT 2324.910 25.400 2325.230 25.460 ;
        RECT 2324.910 25.260 2328.820 25.400 ;
        RECT 2324.910 25.200 2325.230 25.260 ;
        RECT 2328.680 25.060 2328.820 25.260 ;
        RECT 2328.680 24.920 2346.760 25.060 ;
        RECT 2346.620 24.720 2346.760 24.920 ;
        RECT 2845.170 24.720 2845.490 24.780 ;
        RECT 2346.620 24.580 2845.490 24.720 ;
        RECT 2845.170 24.520 2845.490 24.580 ;
      LAYER via ;
        RECT 2320.800 1683.720 2321.060 1683.980 ;
        RECT 2324.940 1683.720 2325.200 1683.980 ;
        RECT 2324.940 25.200 2325.200 25.460 ;
        RECT 2845.200 24.520 2845.460 24.780 ;
      LAYER met2 ;
        RECT 2320.725 1700.000 2321.005 1704.000 ;
        RECT 2320.860 1684.010 2321.000 1700.000 ;
        RECT 2320.800 1683.690 2321.060 1684.010 ;
        RECT 2324.940 1683.690 2325.200 1684.010 ;
        RECT 2325.000 25.490 2325.140 1683.690 ;
        RECT 2324.940 25.170 2325.200 25.490 ;
        RECT 2845.200 24.490 2845.460 24.810 ;
        RECT 2845.260 2.400 2845.400 24.490 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2328.130 1689.020 2328.450 1689.080 ;
        RECT 2330.890 1689.020 2331.210 1689.080 ;
        RECT 2328.130 1688.880 2331.210 1689.020 ;
        RECT 2328.130 1688.820 2328.450 1688.880 ;
        RECT 2330.890 1688.820 2331.210 1688.880 ;
        RECT 2330.890 24.720 2331.210 24.780 ;
        RECT 2330.890 24.580 2346.300 24.720 ;
        RECT 2330.890 24.520 2331.210 24.580 ;
        RECT 2346.160 24.380 2346.300 24.580 ;
        RECT 2863.110 24.380 2863.430 24.440 ;
        RECT 2346.160 24.240 2863.430 24.380 ;
        RECT 2863.110 24.180 2863.430 24.240 ;
      LAYER via ;
        RECT 2328.160 1688.820 2328.420 1689.080 ;
        RECT 2330.920 1688.820 2331.180 1689.080 ;
        RECT 2330.920 24.520 2331.180 24.780 ;
        RECT 2863.140 24.180 2863.400 24.440 ;
      LAYER met2 ;
        RECT 2328.085 1700.000 2328.365 1704.000 ;
        RECT 2328.220 1689.110 2328.360 1700.000 ;
        RECT 2328.160 1688.790 2328.420 1689.110 ;
        RECT 2330.920 1688.790 2331.180 1689.110 ;
        RECT 2330.980 24.810 2331.120 1688.790 ;
        RECT 2330.920 24.490 2331.180 24.810 ;
        RECT 2863.140 24.150 2863.400 24.470 ;
        RECT 2863.200 2.400 2863.340 24.150 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2335.490 1689.020 2335.810 1689.080 ;
        RECT 2338.710 1689.020 2339.030 1689.080 ;
        RECT 2335.490 1688.880 2339.030 1689.020 ;
        RECT 2335.490 1688.820 2335.810 1688.880 ;
        RECT 2338.710 1688.820 2339.030 1688.880 ;
      LAYER via ;
        RECT 2335.520 1688.820 2335.780 1689.080 ;
        RECT 2338.740 1688.820 2339.000 1689.080 ;
      LAYER met2 ;
        RECT 2335.445 1700.000 2335.725 1704.000 ;
        RECT 2335.580 1689.110 2335.720 1700.000 ;
        RECT 2335.520 1688.790 2335.780 1689.110 ;
        RECT 2338.740 1688.790 2339.000 1689.110 ;
        RECT 2338.800 24.325 2338.940 1688.790 ;
        RECT 2338.730 23.955 2339.010 24.325 ;
        RECT 2881.070 23.955 2881.350 24.325 ;
        RECT 2881.140 2.400 2881.280 23.955 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
      LAYER via2 ;
        RECT 2338.730 24.000 2339.010 24.280 ;
        RECT 2881.070 24.000 2881.350 24.280 ;
      LAYER met3 ;
        RECT 2338.705 24.290 2339.035 24.305 ;
        RECT 2881.045 24.290 2881.375 24.305 ;
        RECT 2338.705 23.990 2881.375 24.290 ;
        RECT 2338.705 23.975 2339.035 23.990 ;
        RECT 2881.045 23.975 2881.375 23.990 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2344.690 24.040 2345.010 24.100 ;
        RECT 2898.990 24.040 2899.310 24.100 ;
        RECT 2344.690 23.900 2899.310 24.040 ;
        RECT 2344.690 23.840 2345.010 23.900 ;
        RECT 2898.990 23.840 2899.310 23.900 ;
      LAYER via ;
        RECT 2344.720 23.840 2344.980 24.100 ;
        RECT 2899.020 23.840 2899.280 24.100 ;
      LAYER met2 ;
        RECT 2342.805 1700.410 2343.085 1704.000 ;
        RECT 2342.805 1700.270 2344.920 1700.410 ;
        RECT 2342.805 1700.000 2343.085 1700.270 ;
        RECT 2344.780 24.130 2344.920 1700.270 ;
        RECT 2344.720 23.810 2344.980 24.130 ;
        RECT 2899.020 23.810 2899.280 24.130 ;
        RECT 2899.080 2.400 2899.220 23.810 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1497.830 1656.180 1498.150 1656.440 ;
        RECT 1497.920 1655.760 1498.060 1656.180 ;
        RECT 1497.830 1655.500 1498.150 1655.760 ;
        RECT 848.310 61.780 848.630 61.840 ;
        RECT 1497.830 61.780 1498.150 61.840 ;
        RECT 848.310 61.640 1498.150 61.780 ;
        RECT 848.310 61.580 848.630 61.640 ;
        RECT 1497.830 61.580 1498.150 61.640 ;
        RECT 846.930 2.960 847.250 3.020 ;
        RECT 848.310 2.960 848.630 3.020 ;
        RECT 846.930 2.820 848.630 2.960 ;
        RECT 846.930 2.760 847.250 2.820 ;
        RECT 848.310 2.760 848.630 2.820 ;
      LAYER via ;
        RECT 1497.860 1656.180 1498.120 1656.440 ;
        RECT 1497.860 1655.500 1498.120 1655.760 ;
        RECT 848.340 61.580 848.600 61.840 ;
        RECT 1497.860 61.580 1498.120 61.840 ;
        RECT 846.960 2.760 847.220 3.020 ;
        RECT 848.340 2.760 848.600 3.020 ;
      LAYER met2 ;
        RECT 1497.785 1700.000 1498.065 1704.000 ;
        RECT 1497.920 1656.470 1498.060 1700.000 ;
        RECT 1497.860 1656.150 1498.120 1656.470 ;
        RECT 1497.860 1655.470 1498.120 1655.790 ;
        RECT 1497.920 61.870 1498.060 1655.470 ;
        RECT 848.340 61.550 848.600 61.870 ;
        RECT 1497.860 61.550 1498.120 61.870 ;
        RECT 848.400 3.050 848.540 61.550 ;
        RECT 846.960 2.730 847.220 3.050 ;
        RECT 848.340 2.730 848.600 3.050 ;
        RECT 847.020 2.400 847.160 2.730 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 869.010 62.120 869.330 62.180 ;
        RECT 1504.730 62.120 1505.050 62.180 ;
        RECT 869.010 61.980 1505.050 62.120 ;
        RECT 869.010 61.920 869.330 61.980 ;
        RECT 1504.730 61.920 1505.050 61.980 ;
      LAYER via ;
        RECT 869.040 61.920 869.300 62.180 ;
        RECT 1504.760 61.920 1505.020 62.180 ;
      LAYER met2 ;
        RECT 1505.145 1700.410 1505.425 1704.000 ;
        RECT 1504.820 1700.270 1505.425 1700.410 ;
        RECT 1504.820 62.210 1504.960 1700.270 ;
        RECT 1505.145 1700.000 1505.425 1700.270 ;
        RECT 869.040 61.890 869.300 62.210 ;
        RECT 1504.760 61.890 1505.020 62.210 ;
        RECT 869.100 16.730 869.240 61.890 ;
        RECT 864.960 16.590 869.240 16.730 ;
        RECT 864.960 2.400 865.100 16.590 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 882.350 58.380 882.670 58.440 ;
        RECT 1511.630 58.380 1511.950 58.440 ;
        RECT 882.350 58.240 1511.950 58.380 ;
        RECT 882.350 58.180 882.670 58.240 ;
        RECT 1511.630 58.180 1511.950 58.240 ;
      LAYER via ;
        RECT 882.380 58.180 882.640 58.440 ;
        RECT 1511.660 58.180 1511.920 58.440 ;
      LAYER met2 ;
        RECT 1512.505 1700.410 1512.785 1704.000 ;
        RECT 1511.720 1700.270 1512.785 1700.410 ;
        RECT 1511.720 58.470 1511.860 1700.270 ;
        RECT 1512.505 1700.000 1512.785 1700.270 ;
        RECT 882.380 58.150 882.640 58.470 ;
        RECT 1511.660 58.150 1511.920 58.470 ;
        RECT 882.440 17.410 882.580 58.150 ;
        RECT 882.440 17.270 883.040 17.410 ;
        RECT 882.900 2.400 883.040 17.270 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 903.510 58.040 903.830 58.100 ;
        RECT 1518.530 58.040 1518.850 58.100 ;
        RECT 903.510 57.900 1518.850 58.040 ;
        RECT 903.510 57.840 903.830 57.900 ;
        RECT 1518.530 57.840 1518.850 57.900 ;
      LAYER via ;
        RECT 903.540 57.840 903.800 58.100 ;
        RECT 1518.560 57.840 1518.820 58.100 ;
      LAYER met2 ;
        RECT 1519.405 1700.410 1519.685 1704.000 ;
        RECT 1518.620 1700.270 1519.685 1700.410 ;
        RECT 1518.620 58.130 1518.760 1700.270 ;
        RECT 1519.405 1700.000 1519.685 1700.270 ;
        RECT 903.540 57.810 903.800 58.130 ;
        RECT 1518.560 57.810 1518.820 58.130 ;
        RECT 903.600 16.730 903.740 57.810 ;
        RECT 900.840 16.590 903.740 16.730 ;
        RECT 900.840 2.400 900.980 16.590 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 924.210 57.700 924.530 57.760 ;
        RECT 1525.430 57.700 1525.750 57.760 ;
        RECT 924.210 57.560 1525.750 57.700 ;
        RECT 924.210 57.500 924.530 57.560 ;
        RECT 1525.430 57.500 1525.750 57.560 ;
        RECT 918.690 2.960 919.010 3.020 ;
        RECT 923.750 2.960 924.070 3.020 ;
        RECT 918.690 2.820 924.070 2.960 ;
        RECT 918.690 2.760 919.010 2.820 ;
        RECT 923.750 2.760 924.070 2.820 ;
      LAYER via ;
        RECT 924.240 57.500 924.500 57.760 ;
        RECT 1525.460 57.500 1525.720 57.760 ;
        RECT 918.720 2.760 918.980 3.020 ;
        RECT 923.780 2.760 924.040 3.020 ;
      LAYER met2 ;
        RECT 1526.765 1700.410 1527.045 1704.000 ;
        RECT 1525.520 1700.270 1527.045 1700.410 ;
        RECT 1525.520 57.790 1525.660 1700.270 ;
        RECT 1526.765 1700.000 1527.045 1700.270 ;
        RECT 924.240 57.470 924.500 57.790 ;
        RECT 1525.460 57.470 1525.720 57.790 ;
        RECT 924.300 30.330 924.440 57.470 ;
        RECT 923.840 30.190 924.440 30.330 ;
        RECT 923.840 3.050 923.980 30.190 ;
        RECT 918.720 2.730 918.980 3.050 ;
        RECT 923.780 2.730 924.040 3.050 ;
        RECT 918.780 2.400 918.920 2.730 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1532.330 1666.580 1532.650 1666.640 ;
        RECT 1533.250 1666.580 1533.570 1666.640 ;
        RECT 1532.330 1666.440 1533.570 1666.580 ;
        RECT 1532.330 1666.380 1532.650 1666.440 ;
        RECT 1533.250 1666.380 1533.570 1666.440 ;
        RECT 938.010 57.360 938.330 57.420 ;
        RECT 1532.330 57.360 1532.650 57.420 ;
        RECT 938.010 57.220 1532.650 57.360 ;
        RECT 938.010 57.160 938.330 57.220 ;
        RECT 1532.330 57.160 1532.650 57.220 ;
        RECT 936.170 2.960 936.490 3.020 ;
        RECT 938.010 2.960 938.330 3.020 ;
        RECT 936.170 2.820 938.330 2.960 ;
        RECT 936.170 2.760 936.490 2.820 ;
        RECT 938.010 2.760 938.330 2.820 ;
      LAYER via ;
        RECT 1532.360 1666.380 1532.620 1666.640 ;
        RECT 1533.280 1666.380 1533.540 1666.640 ;
        RECT 938.040 57.160 938.300 57.420 ;
        RECT 1532.360 57.160 1532.620 57.420 ;
        RECT 936.200 2.760 936.460 3.020 ;
        RECT 938.040 2.760 938.300 3.020 ;
      LAYER met2 ;
        RECT 1534.125 1700.410 1534.405 1704.000 ;
        RECT 1533.340 1700.270 1534.405 1700.410 ;
        RECT 1533.340 1666.670 1533.480 1700.270 ;
        RECT 1534.125 1700.000 1534.405 1700.270 ;
        RECT 1532.360 1666.350 1532.620 1666.670 ;
        RECT 1533.280 1666.350 1533.540 1666.670 ;
        RECT 1532.420 57.450 1532.560 1666.350 ;
        RECT 938.040 57.130 938.300 57.450 ;
        RECT 1532.360 57.130 1532.620 57.450 ;
        RECT 938.100 3.050 938.240 57.130 ;
        RECT 936.200 2.730 936.460 3.050 ;
        RECT 938.040 2.730 938.300 3.050 ;
        RECT 936.260 2.400 936.400 2.730 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 958.710 57.020 959.030 57.080 ;
        RECT 1540.150 57.020 1540.470 57.080 ;
        RECT 958.710 56.880 1540.470 57.020 ;
        RECT 958.710 56.820 959.030 56.880 ;
        RECT 1540.150 56.820 1540.470 56.880 ;
      LAYER via ;
        RECT 958.740 56.820 959.000 57.080 ;
        RECT 1540.180 56.820 1540.440 57.080 ;
      LAYER met2 ;
        RECT 1541.485 1700.410 1541.765 1704.000 ;
        RECT 1540.240 1700.270 1541.765 1700.410 ;
        RECT 1540.240 57.110 1540.380 1700.270 ;
        RECT 1541.485 1700.000 1541.765 1700.270 ;
        RECT 958.740 56.790 959.000 57.110 ;
        RECT 1540.180 56.790 1540.440 57.110 ;
        RECT 958.800 16.730 958.940 56.790 ;
        RECT 954.200 16.590 958.940 16.730 ;
        RECT 954.200 2.400 954.340 16.590 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.510 56.680 972.830 56.740 ;
        RECT 1547.050 56.680 1547.370 56.740 ;
        RECT 972.510 56.540 1547.370 56.680 ;
        RECT 972.510 56.480 972.830 56.540 ;
        RECT 1547.050 56.480 1547.370 56.540 ;
      LAYER via ;
        RECT 972.540 56.480 972.800 56.740 ;
        RECT 1547.080 56.480 1547.340 56.740 ;
      LAYER met2 ;
        RECT 1548.845 1700.410 1549.125 1704.000 ;
        RECT 1547.140 1700.270 1549.125 1700.410 ;
        RECT 1547.140 56.770 1547.280 1700.270 ;
        RECT 1548.845 1700.000 1549.125 1700.270 ;
        RECT 972.540 56.450 972.800 56.770 ;
        RECT 1547.080 56.450 1547.340 56.770 ;
        RECT 972.600 17.410 972.740 56.450 ;
        RECT 972.140 17.270 972.740 17.410 ;
        RECT 972.140 2.400 972.280 17.270 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 650.970 26.760 651.290 26.820 ;
        RECT 1415.950 26.760 1416.270 26.820 ;
        RECT 650.970 26.620 1416.270 26.760 ;
        RECT 650.970 26.560 651.290 26.620 ;
        RECT 1415.950 26.560 1416.270 26.620 ;
      LAYER via ;
        RECT 651.000 26.560 651.260 26.820 ;
        RECT 1415.980 26.560 1416.240 26.820 ;
      LAYER met2 ;
        RECT 1416.825 1700.410 1417.105 1704.000 ;
        RECT 1416.040 1700.270 1417.105 1700.410 ;
        RECT 1416.040 26.850 1416.180 1700.270 ;
        RECT 1416.825 1700.000 1417.105 1700.270 ;
        RECT 651.000 26.530 651.260 26.850 ;
        RECT 1415.980 26.530 1416.240 26.850 ;
        RECT 651.060 2.400 651.200 26.530 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1554.485 1539.265 1554.655 1559.835 ;
        RECT 1553.565 1490.645 1553.735 1538.755 ;
        RECT 1554.485 1413.805 1554.655 1465.315 ;
        RECT 1554.485 1317.245 1554.655 1393.575 ;
        RECT 1554.485 1256.385 1554.655 1280.355 ;
        RECT 1553.565 1207.425 1553.735 1255.875 ;
        RECT 1554.025 1110.865 1554.195 1158.975 ;
        RECT 1554.025 1014.305 1554.195 1062.415 ;
        RECT 1554.025 737.885 1554.195 765.935 ;
        RECT 1554.025 607.325 1554.195 628.915 ;
        RECT 1554.025 448.205 1554.195 493.595 ;
        RECT 1554.025 379.525 1554.195 427.635 ;
        RECT 1554.025 303.365 1554.195 331.075 ;
        RECT 1554.485 83.045 1554.655 131.155 ;
      LAYER mcon ;
        RECT 1554.485 1559.665 1554.655 1559.835 ;
        RECT 1553.565 1538.585 1553.735 1538.755 ;
        RECT 1554.485 1465.145 1554.655 1465.315 ;
        RECT 1554.485 1393.405 1554.655 1393.575 ;
        RECT 1554.485 1280.185 1554.655 1280.355 ;
        RECT 1553.565 1255.705 1553.735 1255.875 ;
        RECT 1554.025 1158.805 1554.195 1158.975 ;
        RECT 1554.025 1062.245 1554.195 1062.415 ;
        RECT 1554.025 765.765 1554.195 765.935 ;
        RECT 1554.025 628.745 1554.195 628.915 ;
        RECT 1554.025 493.425 1554.195 493.595 ;
        RECT 1554.025 427.465 1554.195 427.635 ;
        RECT 1554.025 330.905 1554.195 331.075 ;
        RECT 1554.485 130.985 1554.655 131.155 ;
      LAYER met1 ;
        RECT 1553.950 1607.900 1554.270 1608.160 ;
        RECT 1554.040 1607.420 1554.180 1607.900 ;
        RECT 1554.410 1607.420 1554.730 1607.480 ;
        RECT 1554.040 1607.280 1554.730 1607.420 ;
        RECT 1554.410 1607.220 1554.730 1607.280 ;
        RECT 1554.410 1559.820 1554.730 1559.880 ;
        RECT 1554.215 1559.680 1554.730 1559.820 ;
        RECT 1554.410 1559.620 1554.730 1559.680 ;
        RECT 1553.490 1539.420 1553.810 1539.480 ;
        RECT 1554.425 1539.420 1554.715 1539.465 ;
        RECT 1553.490 1539.280 1554.715 1539.420 ;
        RECT 1553.490 1539.220 1553.810 1539.280 ;
        RECT 1554.425 1539.235 1554.715 1539.280 ;
        RECT 1553.490 1538.740 1553.810 1538.800 ;
        RECT 1553.295 1538.600 1553.810 1538.740 ;
        RECT 1553.490 1538.540 1553.810 1538.600 ;
        RECT 1553.505 1490.800 1553.795 1490.845 ;
        RECT 1554.410 1490.800 1554.730 1490.860 ;
        RECT 1553.505 1490.660 1554.730 1490.800 ;
        RECT 1553.505 1490.615 1553.795 1490.660 ;
        RECT 1554.410 1490.600 1554.730 1490.660 ;
        RECT 1554.410 1465.300 1554.730 1465.360 ;
        RECT 1554.215 1465.160 1554.730 1465.300 ;
        RECT 1554.410 1465.100 1554.730 1465.160 ;
        RECT 1554.410 1413.960 1554.730 1414.020 ;
        RECT 1554.215 1413.820 1554.730 1413.960 ;
        RECT 1554.410 1413.760 1554.730 1413.820 ;
        RECT 1554.410 1393.560 1554.730 1393.620 ;
        RECT 1554.215 1393.420 1554.730 1393.560 ;
        RECT 1554.410 1393.360 1554.730 1393.420 ;
        RECT 1554.410 1317.400 1554.730 1317.460 ;
        RECT 1554.215 1317.260 1554.730 1317.400 ;
        RECT 1554.410 1317.200 1554.730 1317.260 ;
        RECT 1554.410 1280.340 1554.730 1280.400 ;
        RECT 1554.215 1280.200 1554.730 1280.340 ;
        RECT 1554.410 1280.140 1554.730 1280.200 ;
        RECT 1553.490 1256.540 1553.810 1256.600 ;
        RECT 1554.425 1256.540 1554.715 1256.585 ;
        RECT 1553.490 1256.400 1554.715 1256.540 ;
        RECT 1553.490 1256.340 1553.810 1256.400 ;
        RECT 1554.425 1256.355 1554.715 1256.400 ;
        RECT 1553.490 1255.860 1553.810 1255.920 ;
        RECT 1553.295 1255.720 1553.810 1255.860 ;
        RECT 1553.490 1255.660 1553.810 1255.720 ;
        RECT 1553.505 1207.580 1553.795 1207.625 ;
        RECT 1554.410 1207.580 1554.730 1207.640 ;
        RECT 1553.505 1207.440 1554.730 1207.580 ;
        RECT 1553.505 1207.395 1553.795 1207.440 ;
        RECT 1554.410 1207.380 1554.730 1207.440 ;
        RECT 1554.410 1173.580 1554.730 1173.640 ;
        RECT 1554.040 1173.440 1554.730 1173.580 ;
        RECT 1554.040 1172.960 1554.180 1173.440 ;
        RECT 1554.410 1173.380 1554.730 1173.440 ;
        RECT 1553.950 1172.700 1554.270 1172.960 ;
        RECT 1553.950 1158.960 1554.270 1159.020 ;
        RECT 1553.755 1158.820 1554.270 1158.960 ;
        RECT 1553.950 1158.760 1554.270 1158.820 ;
        RECT 1553.965 1111.020 1554.255 1111.065 ;
        RECT 1554.410 1111.020 1554.730 1111.080 ;
        RECT 1553.965 1110.880 1554.730 1111.020 ;
        RECT 1553.965 1110.835 1554.255 1110.880 ;
        RECT 1554.410 1110.820 1554.730 1110.880 ;
        RECT 1554.410 1077.020 1554.730 1077.080 ;
        RECT 1554.040 1076.880 1554.730 1077.020 ;
        RECT 1554.040 1076.400 1554.180 1076.880 ;
        RECT 1554.410 1076.820 1554.730 1076.880 ;
        RECT 1553.950 1076.140 1554.270 1076.400 ;
        RECT 1553.950 1062.400 1554.270 1062.460 ;
        RECT 1553.755 1062.260 1554.270 1062.400 ;
        RECT 1553.950 1062.200 1554.270 1062.260 ;
        RECT 1553.965 1014.460 1554.255 1014.505 ;
        RECT 1554.410 1014.460 1554.730 1014.520 ;
        RECT 1553.965 1014.320 1554.730 1014.460 ;
        RECT 1553.965 1014.275 1554.255 1014.320 ;
        RECT 1554.410 1014.260 1554.730 1014.320 ;
        RECT 1554.410 980.460 1554.730 980.520 ;
        RECT 1554.040 980.320 1554.730 980.460 ;
        RECT 1554.040 979.840 1554.180 980.320 ;
        RECT 1554.410 980.260 1554.730 980.320 ;
        RECT 1553.950 979.580 1554.270 979.840 ;
        RECT 1554.410 917.900 1554.730 917.960 ;
        RECT 1555.330 917.900 1555.650 917.960 ;
        RECT 1554.410 917.760 1555.650 917.900 ;
        RECT 1554.410 917.700 1554.730 917.760 ;
        RECT 1555.330 917.700 1555.650 917.760 ;
        RECT 1554.410 883.900 1554.730 883.960 ;
        RECT 1554.040 883.760 1554.730 883.900 ;
        RECT 1554.040 883.280 1554.180 883.760 ;
        RECT 1554.410 883.700 1554.730 883.760 ;
        RECT 1553.950 883.020 1554.270 883.280 ;
        RECT 1553.950 835.080 1554.270 835.340 ;
        RECT 1554.040 834.600 1554.180 835.080 ;
        RECT 1554.410 834.600 1554.730 834.660 ;
        RECT 1554.040 834.460 1554.730 834.600 ;
        RECT 1554.410 834.400 1554.730 834.460 ;
        RECT 1553.950 765.920 1554.270 765.980 ;
        RECT 1553.755 765.780 1554.270 765.920 ;
        RECT 1553.950 765.720 1554.270 765.780 ;
        RECT 1553.950 738.040 1554.270 738.100 ;
        RECT 1553.755 737.900 1554.270 738.040 ;
        RECT 1553.950 737.840 1554.270 737.900 ;
        RECT 1554.410 690.440 1554.730 690.500 ;
        RECT 1554.040 690.300 1554.730 690.440 ;
        RECT 1554.040 689.820 1554.180 690.300 ;
        RECT 1554.410 690.240 1554.730 690.300 ;
        RECT 1553.950 689.560 1554.270 689.820 ;
        RECT 1553.950 628.900 1554.270 628.960 ;
        RECT 1553.755 628.760 1554.270 628.900 ;
        RECT 1553.950 628.700 1554.270 628.760 ;
        RECT 1553.950 607.480 1554.270 607.540 ;
        RECT 1553.755 607.340 1554.270 607.480 ;
        RECT 1553.950 607.280 1554.270 607.340 ;
        RECT 1553.950 559.200 1554.270 559.260 ;
        RECT 1554.870 559.200 1555.190 559.260 ;
        RECT 1553.950 559.060 1555.190 559.200 ;
        RECT 1553.950 559.000 1554.270 559.060 ;
        RECT 1554.870 559.000 1555.190 559.060 ;
        RECT 1554.870 511.260 1555.190 511.320 ;
        RECT 1554.500 511.120 1555.190 511.260 ;
        RECT 1554.500 510.980 1554.640 511.120 ;
        RECT 1554.870 511.060 1555.190 511.120 ;
        RECT 1554.410 510.720 1554.730 510.980 ;
        RECT 1553.965 493.580 1554.255 493.625 ;
        RECT 1554.410 493.580 1554.730 493.640 ;
        RECT 1553.965 493.440 1554.730 493.580 ;
        RECT 1553.965 493.395 1554.255 493.440 ;
        RECT 1554.410 493.380 1554.730 493.440 ;
        RECT 1553.950 448.360 1554.270 448.420 ;
        RECT 1553.755 448.220 1554.270 448.360 ;
        RECT 1553.950 448.160 1554.270 448.220 ;
        RECT 1553.950 427.620 1554.270 427.680 ;
        RECT 1553.755 427.480 1554.270 427.620 ;
        RECT 1553.950 427.420 1554.270 427.480 ;
        RECT 1553.950 379.680 1554.270 379.740 ;
        RECT 1553.755 379.540 1554.270 379.680 ;
        RECT 1553.950 379.480 1554.270 379.540 ;
        RECT 1553.950 331.060 1554.270 331.120 ;
        RECT 1553.755 330.920 1554.270 331.060 ;
        RECT 1553.950 330.860 1554.270 330.920 ;
        RECT 1553.950 303.520 1554.270 303.580 ;
        RECT 1553.755 303.380 1554.270 303.520 ;
        RECT 1553.950 303.320 1554.270 303.380 ;
        RECT 1553.950 282.780 1554.270 282.840 ;
        RECT 1554.410 282.780 1554.730 282.840 ;
        RECT 1553.950 282.640 1554.730 282.780 ;
        RECT 1553.950 282.580 1554.270 282.640 ;
        RECT 1554.410 282.580 1554.730 282.640 ;
        RECT 1554.410 227.700 1554.730 227.760 ;
        RECT 1555.330 227.700 1555.650 227.760 ;
        RECT 1554.410 227.560 1555.650 227.700 ;
        RECT 1554.410 227.500 1554.730 227.560 ;
        RECT 1555.330 227.500 1555.650 227.560 ;
        RECT 1554.410 131.140 1554.730 131.200 ;
        RECT 1554.215 131.000 1554.730 131.140 ;
        RECT 1554.410 130.940 1554.730 131.000 ;
        RECT 1554.410 83.200 1554.730 83.260 ;
        RECT 1554.215 83.060 1554.730 83.200 ;
        RECT 1554.410 83.000 1554.730 83.060 ;
        RECT 993.210 56.340 993.530 56.400 ;
        RECT 1554.410 56.340 1554.730 56.400 ;
        RECT 993.210 56.200 1554.730 56.340 ;
        RECT 993.210 56.140 993.530 56.200 ;
        RECT 1554.410 56.140 1554.730 56.200 ;
      LAYER via ;
        RECT 1553.980 1607.900 1554.240 1608.160 ;
        RECT 1554.440 1607.220 1554.700 1607.480 ;
        RECT 1554.440 1559.620 1554.700 1559.880 ;
        RECT 1553.520 1539.220 1553.780 1539.480 ;
        RECT 1553.520 1538.540 1553.780 1538.800 ;
        RECT 1554.440 1490.600 1554.700 1490.860 ;
        RECT 1554.440 1465.100 1554.700 1465.360 ;
        RECT 1554.440 1413.760 1554.700 1414.020 ;
        RECT 1554.440 1393.360 1554.700 1393.620 ;
        RECT 1554.440 1317.200 1554.700 1317.460 ;
        RECT 1554.440 1280.140 1554.700 1280.400 ;
        RECT 1553.520 1256.340 1553.780 1256.600 ;
        RECT 1553.520 1255.660 1553.780 1255.920 ;
        RECT 1554.440 1207.380 1554.700 1207.640 ;
        RECT 1554.440 1173.380 1554.700 1173.640 ;
        RECT 1553.980 1172.700 1554.240 1172.960 ;
        RECT 1553.980 1158.760 1554.240 1159.020 ;
        RECT 1554.440 1110.820 1554.700 1111.080 ;
        RECT 1554.440 1076.820 1554.700 1077.080 ;
        RECT 1553.980 1076.140 1554.240 1076.400 ;
        RECT 1553.980 1062.200 1554.240 1062.460 ;
        RECT 1554.440 1014.260 1554.700 1014.520 ;
        RECT 1554.440 980.260 1554.700 980.520 ;
        RECT 1553.980 979.580 1554.240 979.840 ;
        RECT 1554.440 917.700 1554.700 917.960 ;
        RECT 1555.360 917.700 1555.620 917.960 ;
        RECT 1554.440 883.700 1554.700 883.960 ;
        RECT 1553.980 883.020 1554.240 883.280 ;
        RECT 1553.980 835.080 1554.240 835.340 ;
        RECT 1554.440 834.400 1554.700 834.660 ;
        RECT 1553.980 765.720 1554.240 765.980 ;
        RECT 1553.980 737.840 1554.240 738.100 ;
        RECT 1554.440 690.240 1554.700 690.500 ;
        RECT 1553.980 689.560 1554.240 689.820 ;
        RECT 1553.980 628.700 1554.240 628.960 ;
        RECT 1553.980 607.280 1554.240 607.540 ;
        RECT 1553.980 559.000 1554.240 559.260 ;
        RECT 1554.900 559.000 1555.160 559.260 ;
        RECT 1554.900 511.060 1555.160 511.320 ;
        RECT 1554.440 510.720 1554.700 510.980 ;
        RECT 1554.440 493.380 1554.700 493.640 ;
        RECT 1553.980 448.160 1554.240 448.420 ;
        RECT 1553.980 427.420 1554.240 427.680 ;
        RECT 1553.980 379.480 1554.240 379.740 ;
        RECT 1553.980 330.860 1554.240 331.120 ;
        RECT 1553.980 303.320 1554.240 303.580 ;
        RECT 1553.980 282.580 1554.240 282.840 ;
        RECT 1554.440 282.580 1554.700 282.840 ;
        RECT 1554.440 227.500 1554.700 227.760 ;
        RECT 1555.360 227.500 1555.620 227.760 ;
        RECT 1554.440 130.940 1554.700 131.200 ;
        RECT 1554.440 83.000 1554.700 83.260 ;
        RECT 993.240 56.140 993.500 56.400 ;
        RECT 1554.440 56.140 1554.700 56.400 ;
      LAYER met2 ;
        RECT 1556.205 1700.410 1556.485 1704.000 ;
        RECT 1555.420 1700.270 1556.485 1700.410 ;
        RECT 1555.420 1656.210 1555.560 1700.270 ;
        RECT 1556.205 1700.000 1556.485 1700.270 ;
        RECT 1554.040 1656.070 1555.560 1656.210 ;
        RECT 1554.040 1608.190 1554.180 1656.070 ;
        RECT 1553.980 1607.870 1554.240 1608.190 ;
        RECT 1554.440 1607.190 1554.700 1607.510 ;
        RECT 1554.500 1559.910 1554.640 1607.190 ;
        RECT 1554.440 1559.590 1554.700 1559.910 ;
        RECT 1553.520 1539.190 1553.780 1539.510 ;
        RECT 1553.580 1538.830 1553.720 1539.190 ;
        RECT 1553.520 1538.510 1553.780 1538.830 ;
        RECT 1554.440 1490.570 1554.700 1490.890 ;
        RECT 1554.500 1465.390 1554.640 1490.570 ;
        RECT 1554.440 1465.070 1554.700 1465.390 ;
        RECT 1554.440 1413.730 1554.700 1414.050 ;
        RECT 1554.500 1393.650 1554.640 1413.730 ;
        RECT 1554.440 1393.330 1554.700 1393.650 ;
        RECT 1554.440 1317.170 1554.700 1317.490 ;
        RECT 1554.500 1280.430 1554.640 1317.170 ;
        RECT 1554.440 1280.110 1554.700 1280.430 ;
        RECT 1553.520 1256.310 1553.780 1256.630 ;
        RECT 1553.580 1255.950 1553.720 1256.310 ;
        RECT 1553.520 1255.630 1553.780 1255.950 ;
        RECT 1554.440 1207.350 1554.700 1207.670 ;
        RECT 1554.500 1173.670 1554.640 1207.350 ;
        RECT 1554.440 1173.350 1554.700 1173.670 ;
        RECT 1553.980 1172.670 1554.240 1172.990 ;
        RECT 1554.040 1159.050 1554.180 1172.670 ;
        RECT 1553.980 1158.730 1554.240 1159.050 ;
        RECT 1554.440 1110.790 1554.700 1111.110 ;
        RECT 1554.500 1077.110 1554.640 1110.790 ;
        RECT 1554.440 1076.790 1554.700 1077.110 ;
        RECT 1553.980 1076.110 1554.240 1076.430 ;
        RECT 1554.040 1062.490 1554.180 1076.110 ;
        RECT 1553.980 1062.170 1554.240 1062.490 ;
        RECT 1554.440 1014.230 1554.700 1014.550 ;
        RECT 1554.500 980.550 1554.640 1014.230 ;
        RECT 1554.440 980.230 1554.700 980.550 ;
        RECT 1553.980 979.550 1554.240 979.870 ;
        RECT 1554.040 966.125 1554.180 979.550 ;
        RECT 1553.970 965.755 1554.250 966.125 ;
        RECT 1555.350 965.755 1555.630 966.125 ;
        RECT 1555.420 917.990 1555.560 965.755 ;
        RECT 1554.440 917.670 1554.700 917.990 ;
        RECT 1555.360 917.670 1555.620 917.990 ;
        RECT 1554.500 883.990 1554.640 917.670 ;
        RECT 1554.440 883.670 1554.700 883.990 ;
        RECT 1553.980 882.990 1554.240 883.310 ;
        RECT 1554.040 835.370 1554.180 882.990 ;
        RECT 1553.980 835.050 1554.240 835.370 ;
        RECT 1554.440 834.370 1554.700 834.690 ;
        RECT 1554.500 766.885 1554.640 834.370 ;
        RECT 1554.430 766.515 1554.710 766.885 ;
        RECT 1553.970 765.835 1554.250 766.205 ;
        RECT 1553.980 765.690 1554.240 765.835 ;
        RECT 1553.980 737.810 1554.240 738.130 ;
        RECT 1554.040 717.810 1554.180 737.810 ;
        RECT 1554.040 717.670 1554.640 717.810 ;
        RECT 1554.500 690.530 1554.640 717.670 ;
        RECT 1554.440 690.210 1554.700 690.530 ;
        RECT 1553.980 689.530 1554.240 689.850 ;
        RECT 1554.040 628.990 1554.180 689.530 ;
        RECT 1553.980 628.670 1554.240 628.990 ;
        RECT 1553.980 607.250 1554.240 607.570 ;
        RECT 1554.040 559.290 1554.180 607.250 ;
        RECT 1553.980 558.970 1554.240 559.290 ;
        RECT 1554.900 558.970 1555.160 559.290 ;
        RECT 1554.960 511.350 1555.100 558.970 ;
        RECT 1554.900 511.030 1555.160 511.350 ;
        RECT 1554.440 510.690 1554.700 511.010 ;
        RECT 1554.500 493.670 1554.640 510.690 ;
        RECT 1554.440 493.350 1554.700 493.670 ;
        RECT 1553.980 448.130 1554.240 448.450 ;
        RECT 1554.040 427.710 1554.180 448.130 ;
        RECT 1553.980 427.390 1554.240 427.710 ;
        RECT 1553.980 379.450 1554.240 379.770 ;
        RECT 1554.040 379.285 1554.180 379.450 ;
        RECT 1552.130 378.915 1552.410 379.285 ;
        RECT 1553.970 378.915 1554.250 379.285 ;
        RECT 1552.200 331.685 1552.340 378.915 ;
        RECT 1552.130 331.315 1552.410 331.685 ;
        RECT 1553.970 331.315 1554.250 331.685 ;
        RECT 1554.040 331.150 1554.180 331.315 ;
        RECT 1553.980 330.830 1554.240 331.150 ;
        RECT 1553.980 303.290 1554.240 303.610 ;
        RECT 1554.040 282.870 1554.180 303.290 ;
        RECT 1553.980 282.550 1554.240 282.870 ;
        RECT 1554.440 282.550 1554.700 282.870 ;
        RECT 1554.500 227.790 1554.640 282.550 ;
        RECT 1554.440 227.470 1554.700 227.790 ;
        RECT 1555.360 227.470 1555.620 227.790 ;
        RECT 1555.420 138.450 1555.560 227.470 ;
        RECT 1554.500 138.310 1555.560 138.450 ;
        RECT 1554.500 131.230 1554.640 138.310 ;
        RECT 1554.440 130.910 1554.700 131.230 ;
        RECT 1554.440 82.970 1554.700 83.290 ;
        RECT 1554.500 56.430 1554.640 82.970 ;
        RECT 993.240 56.110 993.500 56.430 ;
        RECT 1554.440 56.110 1554.700 56.430 ;
        RECT 993.300 16.730 993.440 56.110 ;
        RECT 990.080 16.590 993.440 16.730 ;
        RECT 990.080 2.400 990.220 16.590 ;
        RECT 989.870 -4.800 990.430 2.400 ;
      LAYER via2 ;
        RECT 1553.970 965.800 1554.250 966.080 ;
        RECT 1555.350 965.800 1555.630 966.080 ;
        RECT 1554.430 766.560 1554.710 766.840 ;
        RECT 1553.970 765.880 1554.250 766.160 ;
        RECT 1552.130 378.960 1552.410 379.240 ;
        RECT 1553.970 378.960 1554.250 379.240 ;
        RECT 1552.130 331.360 1552.410 331.640 ;
        RECT 1553.970 331.360 1554.250 331.640 ;
      LAYER met3 ;
        RECT 1553.945 966.090 1554.275 966.105 ;
        RECT 1555.325 966.090 1555.655 966.105 ;
        RECT 1553.945 965.790 1555.655 966.090 ;
        RECT 1553.945 965.775 1554.275 965.790 ;
        RECT 1555.325 965.775 1555.655 965.790 ;
        RECT 1554.405 766.850 1554.735 766.865 ;
        RECT 1554.190 766.535 1554.735 766.850 ;
        RECT 1554.190 766.185 1554.490 766.535 ;
        RECT 1553.945 765.870 1554.490 766.185 ;
        RECT 1553.945 765.855 1554.275 765.870 ;
        RECT 1552.105 379.250 1552.435 379.265 ;
        RECT 1553.945 379.250 1554.275 379.265 ;
        RECT 1552.105 378.950 1554.275 379.250 ;
        RECT 1552.105 378.935 1552.435 378.950 ;
        RECT 1553.945 378.935 1554.275 378.950 ;
        RECT 1552.105 331.650 1552.435 331.665 ;
        RECT 1553.945 331.650 1554.275 331.665 ;
        RECT 1552.105 331.350 1554.275 331.650 ;
        RECT 1552.105 331.335 1552.435 331.350 ;
        RECT 1553.945 331.335 1554.275 331.350 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1356.610 1686.300 1356.930 1686.360 ;
        RECT 1562.230 1686.300 1562.550 1686.360 ;
        RECT 1356.610 1686.160 1562.550 1686.300 ;
        RECT 1356.610 1686.100 1356.930 1686.160 ;
        RECT 1562.230 1686.100 1562.550 1686.160 ;
        RECT 1007.470 22.000 1007.790 22.060 ;
        RECT 1355.690 22.000 1356.010 22.060 ;
        RECT 1007.470 21.860 1356.010 22.000 ;
        RECT 1007.470 21.800 1007.790 21.860 ;
        RECT 1355.690 21.800 1356.010 21.860 ;
      LAYER via ;
        RECT 1356.640 1686.100 1356.900 1686.360 ;
        RECT 1562.260 1686.100 1562.520 1686.360 ;
        RECT 1007.500 21.800 1007.760 22.060 ;
        RECT 1355.720 21.800 1355.980 22.060 ;
      LAYER met2 ;
        RECT 1563.565 1700.410 1563.845 1704.000 ;
        RECT 1562.320 1700.270 1563.845 1700.410 ;
        RECT 1562.320 1686.390 1562.460 1700.270 ;
        RECT 1563.565 1700.000 1563.845 1700.270 ;
        RECT 1356.640 1686.070 1356.900 1686.390 ;
        RECT 1562.260 1686.070 1562.520 1686.390 ;
        RECT 1356.700 1671.170 1356.840 1686.070 ;
        RECT 1355.780 1671.030 1356.840 1671.170 ;
        RECT 1355.780 22.090 1355.920 1671.030 ;
        RECT 1007.500 21.770 1007.760 22.090 ;
        RECT 1355.720 21.770 1355.980 22.090 ;
        RECT 1007.560 2.400 1007.700 21.770 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1363.970 1686.640 1364.290 1686.700 ;
        RECT 1570.970 1686.640 1571.290 1686.700 ;
        RECT 1363.970 1686.500 1571.290 1686.640 ;
        RECT 1363.970 1686.440 1364.290 1686.500 ;
        RECT 1570.970 1686.440 1571.290 1686.500 ;
        RECT 1025.410 21.660 1025.730 21.720 ;
        RECT 1362.590 21.660 1362.910 21.720 ;
        RECT 1025.410 21.520 1362.910 21.660 ;
        RECT 1025.410 21.460 1025.730 21.520 ;
        RECT 1362.590 21.460 1362.910 21.520 ;
      LAYER via ;
        RECT 1364.000 1686.440 1364.260 1686.700 ;
        RECT 1571.000 1686.440 1571.260 1686.700 ;
        RECT 1025.440 21.460 1025.700 21.720 ;
        RECT 1362.620 21.460 1362.880 21.720 ;
      LAYER met2 ;
        RECT 1570.925 1700.000 1571.205 1704.000 ;
        RECT 1571.060 1686.730 1571.200 1700.000 ;
        RECT 1364.000 1686.410 1364.260 1686.730 ;
        RECT 1571.000 1686.410 1571.260 1686.730 ;
        RECT 1364.060 1671.170 1364.200 1686.410 ;
        RECT 1362.680 1671.030 1364.200 1671.170 ;
        RECT 1362.680 21.750 1362.820 1671.030 ;
        RECT 1025.440 21.430 1025.700 21.750 ;
        RECT 1362.620 21.430 1362.880 21.750 ;
        RECT 1025.500 2.400 1025.640 21.430 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1573.270 1687.320 1573.590 1687.380 ;
        RECT 1576.950 1687.320 1577.270 1687.380 ;
        RECT 1573.270 1687.180 1577.270 1687.320 ;
        RECT 1573.270 1687.120 1573.590 1687.180 ;
        RECT 1576.950 1687.120 1577.270 1687.180 ;
      LAYER via ;
        RECT 1573.300 1687.120 1573.560 1687.380 ;
        RECT 1576.980 1687.120 1577.240 1687.380 ;
      LAYER met2 ;
        RECT 1578.285 1700.410 1578.565 1704.000 ;
        RECT 1577.040 1700.270 1578.565 1700.410 ;
        RECT 1577.040 1687.410 1577.180 1700.270 ;
        RECT 1578.285 1700.000 1578.565 1700.270 ;
        RECT 1573.300 1687.090 1573.560 1687.410 ;
        RECT 1576.980 1687.090 1577.240 1687.410 ;
        RECT 1573.360 24.325 1573.500 1687.090 ;
        RECT 1043.370 23.955 1043.650 24.325 ;
        RECT 1573.290 23.955 1573.570 24.325 ;
        RECT 1043.440 2.400 1043.580 23.955 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
      LAYER via2 ;
        RECT 1043.370 24.000 1043.650 24.280 ;
        RECT 1573.290 24.000 1573.570 24.280 ;
      LAYER met3 ;
        RECT 1043.345 24.290 1043.675 24.305 ;
        RECT 1573.265 24.290 1573.595 24.305 ;
        RECT 1043.345 23.990 1573.595 24.290 ;
        RECT 1043.345 23.975 1043.675 23.990 ;
        RECT 1573.265 23.975 1573.595 23.990 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1580.170 1686.640 1580.490 1686.700 ;
        RECT 1584.310 1686.640 1584.630 1686.700 ;
        RECT 1580.170 1686.500 1584.630 1686.640 ;
        RECT 1580.170 1686.440 1580.490 1686.500 ;
        RECT 1584.310 1686.440 1584.630 1686.500 ;
        RECT 1061.290 23.700 1061.610 23.760 ;
        RECT 1580.170 23.700 1580.490 23.760 ;
        RECT 1061.290 23.560 1580.490 23.700 ;
        RECT 1061.290 23.500 1061.610 23.560 ;
        RECT 1580.170 23.500 1580.490 23.560 ;
      LAYER via ;
        RECT 1580.200 1686.440 1580.460 1686.700 ;
        RECT 1584.340 1686.440 1584.600 1686.700 ;
        RECT 1061.320 23.500 1061.580 23.760 ;
        RECT 1580.200 23.500 1580.460 23.760 ;
      LAYER met2 ;
        RECT 1585.645 1700.410 1585.925 1704.000 ;
        RECT 1584.400 1700.270 1585.925 1700.410 ;
        RECT 1584.400 1686.730 1584.540 1700.270 ;
        RECT 1585.645 1700.000 1585.925 1700.270 ;
        RECT 1580.200 1686.410 1580.460 1686.730 ;
        RECT 1584.340 1686.410 1584.600 1686.730 ;
        RECT 1580.260 23.790 1580.400 1686.410 ;
        RECT 1061.320 23.470 1061.580 23.790 ;
        RECT 1580.200 23.470 1580.460 23.790 ;
        RECT 1061.380 2.400 1061.520 23.470 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1587.070 1687.320 1587.390 1687.380 ;
        RECT 1591.670 1687.320 1591.990 1687.380 ;
        RECT 1587.070 1687.180 1591.990 1687.320 ;
        RECT 1587.070 1687.120 1587.390 1687.180 ;
        RECT 1591.670 1687.120 1591.990 1687.180 ;
        RECT 1079.230 23.360 1079.550 23.420 ;
        RECT 1587.070 23.360 1587.390 23.420 ;
        RECT 1079.230 23.220 1587.390 23.360 ;
        RECT 1079.230 23.160 1079.550 23.220 ;
        RECT 1587.070 23.160 1587.390 23.220 ;
      LAYER via ;
        RECT 1587.100 1687.120 1587.360 1687.380 ;
        RECT 1591.700 1687.120 1591.960 1687.380 ;
        RECT 1079.260 23.160 1079.520 23.420 ;
        RECT 1587.100 23.160 1587.360 23.420 ;
      LAYER met2 ;
        RECT 1593.005 1700.410 1593.285 1704.000 ;
        RECT 1591.760 1700.270 1593.285 1700.410 ;
        RECT 1591.760 1687.410 1591.900 1700.270 ;
        RECT 1593.005 1700.000 1593.285 1700.270 ;
        RECT 1587.100 1687.090 1587.360 1687.410 ;
        RECT 1591.700 1687.090 1591.960 1687.410 ;
        RECT 1587.160 23.450 1587.300 1687.090 ;
        RECT 1079.260 23.130 1079.520 23.450 ;
        RECT 1587.100 23.130 1587.360 23.450 ;
        RECT 1079.320 2.400 1079.460 23.130 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1593.970 1686.640 1594.290 1686.700 ;
        RECT 1599.030 1686.640 1599.350 1686.700 ;
        RECT 1593.970 1686.500 1599.350 1686.640 ;
        RECT 1593.970 1686.440 1594.290 1686.500 ;
        RECT 1599.030 1686.440 1599.350 1686.500 ;
        RECT 1096.710 23.020 1097.030 23.080 ;
        RECT 1593.970 23.020 1594.290 23.080 ;
        RECT 1096.710 22.880 1594.290 23.020 ;
        RECT 1096.710 22.820 1097.030 22.880 ;
        RECT 1593.970 22.820 1594.290 22.880 ;
      LAYER via ;
        RECT 1594.000 1686.440 1594.260 1686.700 ;
        RECT 1599.060 1686.440 1599.320 1686.700 ;
        RECT 1096.740 22.820 1097.000 23.080 ;
        RECT 1594.000 22.820 1594.260 23.080 ;
      LAYER met2 ;
        RECT 1600.365 1700.410 1600.645 1704.000 ;
        RECT 1599.120 1700.270 1600.645 1700.410 ;
        RECT 1599.120 1686.730 1599.260 1700.270 ;
        RECT 1600.365 1700.000 1600.645 1700.270 ;
        RECT 1594.000 1686.410 1594.260 1686.730 ;
        RECT 1599.060 1686.410 1599.320 1686.730 ;
        RECT 1594.060 23.110 1594.200 1686.410 ;
        RECT 1096.740 22.790 1097.000 23.110 ;
        RECT 1594.000 22.790 1594.260 23.110 ;
        RECT 1096.800 2.400 1096.940 22.790 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1606.850 23.020 1607.170 23.080 ;
        RECT 1594.520 22.880 1607.170 23.020 ;
        RECT 1114.650 22.680 1114.970 22.740 ;
        RECT 1594.520 22.680 1594.660 22.880 ;
        RECT 1606.850 22.820 1607.170 22.880 ;
        RECT 1114.650 22.540 1594.660 22.680 ;
        RECT 1114.650 22.480 1114.970 22.540 ;
      LAYER via ;
        RECT 1114.680 22.480 1114.940 22.740 ;
        RECT 1606.880 22.820 1607.140 23.080 ;
      LAYER met2 ;
        RECT 1607.725 1700.000 1608.005 1704.000 ;
        RECT 1607.860 23.530 1608.000 1700.000 ;
        RECT 1606.940 23.390 1608.000 23.530 ;
        RECT 1606.940 23.110 1607.080 23.390 ;
        RECT 1606.880 22.790 1607.140 23.110 ;
        RECT 1114.680 22.450 1114.940 22.770 ;
        RECT 1114.740 2.400 1114.880 22.450 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1132.590 22.340 1132.910 22.400 ;
        RECT 1614.670 22.340 1614.990 22.400 ;
        RECT 1132.590 22.200 1614.990 22.340 ;
        RECT 1132.590 22.140 1132.910 22.200 ;
        RECT 1614.670 22.140 1614.990 22.200 ;
      LAYER via ;
        RECT 1132.620 22.140 1132.880 22.400 ;
        RECT 1614.700 22.140 1614.960 22.400 ;
      LAYER met2 ;
        RECT 1615.085 1700.410 1615.365 1704.000 ;
        RECT 1614.760 1700.270 1615.365 1700.410 ;
        RECT 1614.760 22.430 1614.900 1700.270 ;
        RECT 1615.085 1700.000 1615.365 1700.270 ;
        RECT 1132.620 22.110 1132.880 22.430 ;
        RECT 1614.700 22.110 1614.960 22.430 ;
        RECT 1132.680 2.400 1132.820 22.110 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1150.530 24.380 1150.850 24.440 ;
        RECT 1621.570 24.380 1621.890 24.440 ;
        RECT 1150.530 24.240 1621.890 24.380 ;
        RECT 1150.530 24.180 1150.850 24.240 ;
        RECT 1621.570 24.180 1621.890 24.240 ;
      LAYER via ;
        RECT 1150.560 24.180 1150.820 24.440 ;
        RECT 1621.600 24.180 1621.860 24.440 ;
      LAYER met2 ;
        RECT 1622.445 1700.410 1622.725 1704.000 ;
        RECT 1621.660 1700.270 1622.725 1700.410 ;
        RECT 1621.660 24.470 1621.800 1700.270 ;
        RECT 1622.445 1700.000 1622.725 1700.270 ;
        RECT 1150.560 24.150 1150.820 24.470 ;
        RECT 1621.600 24.150 1621.860 24.470 ;
        RECT 1150.620 2.400 1150.760 24.150 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1421.470 1684.600 1421.790 1684.660 ;
        RECT 1424.230 1684.600 1424.550 1684.660 ;
        RECT 1421.470 1684.460 1424.550 1684.600 ;
        RECT 1421.470 1684.400 1421.790 1684.460 ;
        RECT 1424.230 1684.400 1424.550 1684.460 ;
        RECT 668.910 27.100 669.230 27.160 ;
        RECT 1421.470 27.100 1421.790 27.160 ;
        RECT 668.910 26.960 1421.790 27.100 ;
        RECT 668.910 26.900 669.230 26.960 ;
        RECT 1421.470 26.900 1421.790 26.960 ;
      LAYER via ;
        RECT 1421.500 1684.400 1421.760 1684.660 ;
        RECT 1424.260 1684.400 1424.520 1684.660 ;
        RECT 668.940 26.900 669.200 27.160 ;
        RECT 1421.500 26.900 1421.760 27.160 ;
      LAYER met2 ;
        RECT 1424.185 1700.000 1424.465 1704.000 ;
        RECT 1424.320 1684.690 1424.460 1700.000 ;
        RECT 1421.500 1684.370 1421.760 1684.690 ;
        RECT 1424.260 1684.370 1424.520 1684.690 ;
        RECT 1421.560 27.190 1421.700 1684.370 ;
        RECT 668.940 26.870 669.200 27.190 ;
        RECT 1421.500 26.870 1421.760 27.190 ;
        RECT 669.000 2.400 669.140 26.870 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1168.470 24.040 1168.790 24.100 ;
        RECT 1628.470 24.040 1628.790 24.100 ;
        RECT 1168.470 23.900 1628.790 24.040 ;
        RECT 1168.470 23.840 1168.790 23.900 ;
        RECT 1628.470 23.840 1628.790 23.900 ;
      LAYER via ;
        RECT 1168.500 23.840 1168.760 24.100 ;
        RECT 1628.500 23.840 1628.760 24.100 ;
      LAYER met2 ;
        RECT 1629.805 1700.410 1630.085 1704.000 ;
        RECT 1628.560 1700.270 1630.085 1700.410 ;
        RECT 1628.560 24.130 1628.700 1700.270 ;
        RECT 1629.805 1700.000 1630.085 1700.270 ;
        RECT 1168.500 23.810 1168.760 24.130 ;
        RECT 1628.500 23.810 1628.760 24.130 ;
        RECT 1168.560 2.400 1168.700 23.810 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1608.230 25.400 1608.550 25.460 ;
        RECT 1635.370 25.400 1635.690 25.460 ;
        RECT 1608.230 25.260 1635.690 25.400 ;
        RECT 1608.230 25.200 1608.550 25.260 ;
        RECT 1635.370 25.200 1635.690 25.260 ;
        RECT 1185.950 24.720 1186.270 24.780 ;
        RECT 1608.230 24.720 1608.550 24.780 ;
        RECT 1185.950 24.580 1608.550 24.720 ;
        RECT 1185.950 24.520 1186.270 24.580 ;
        RECT 1608.230 24.520 1608.550 24.580 ;
      LAYER via ;
        RECT 1608.260 25.200 1608.520 25.460 ;
        RECT 1635.400 25.200 1635.660 25.460 ;
        RECT 1185.980 24.520 1186.240 24.780 ;
        RECT 1608.260 24.520 1608.520 24.780 ;
      LAYER met2 ;
        RECT 1637.165 1700.410 1637.445 1704.000 ;
        RECT 1635.460 1700.270 1637.445 1700.410 ;
        RECT 1635.460 25.490 1635.600 1700.270 ;
        RECT 1637.165 1700.000 1637.445 1700.270 ;
        RECT 1608.260 25.170 1608.520 25.490 ;
        RECT 1635.400 25.170 1635.660 25.490 ;
        RECT 1608.320 24.810 1608.460 25.170 ;
        RECT 1185.980 24.490 1186.240 24.810 ;
        RECT 1608.260 24.490 1608.520 24.810 ;
        RECT 1186.040 2.400 1186.180 24.490 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1203.890 25.060 1204.210 25.120 ;
        RECT 1643.650 25.060 1643.970 25.120 ;
        RECT 1203.890 24.920 1643.970 25.060 ;
        RECT 1203.890 24.860 1204.210 24.920 ;
        RECT 1643.650 24.860 1643.970 24.920 ;
      LAYER via ;
        RECT 1203.920 24.860 1204.180 25.120 ;
        RECT 1643.680 24.860 1643.940 25.120 ;
      LAYER met2 ;
        RECT 1644.525 1700.410 1644.805 1704.000 ;
        RECT 1643.740 1700.270 1644.805 1700.410 ;
        RECT 1643.740 25.150 1643.880 1700.270 ;
        RECT 1644.525 1700.000 1644.805 1700.270 ;
        RECT 1203.920 24.830 1204.180 25.150 ;
        RECT 1643.680 24.830 1643.940 25.150 ;
        RECT 1203.980 2.400 1204.120 24.830 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1607.845 24.735 1608.015 25.415 ;
        RECT 1635.905 24.735 1636.075 25.415 ;
        RECT 1607.845 24.565 1608.935 24.735 ;
        RECT 1634.985 24.565 1636.075 24.735 ;
      LAYER mcon ;
        RECT 1607.845 25.245 1608.015 25.415 ;
        RECT 1635.905 25.245 1636.075 25.415 ;
        RECT 1608.765 24.565 1608.935 24.735 ;
      LAYER met1 ;
        RECT 1649.170 1678.140 1649.490 1678.200 ;
        RECT 1650.550 1678.140 1650.870 1678.200 ;
        RECT 1649.170 1678.000 1650.870 1678.140 ;
        RECT 1649.170 1677.940 1649.490 1678.000 ;
        RECT 1650.550 1677.940 1650.870 1678.000 ;
        RECT 1221.830 25.400 1222.150 25.460 ;
        RECT 1607.785 25.400 1608.075 25.445 ;
        RECT 1221.830 25.260 1608.075 25.400 ;
        RECT 1221.830 25.200 1222.150 25.260 ;
        RECT 1607.785 25.215 1608.075 25.260 ;
        RECT 1635.845 25.400 1636.135 25.445 ;
        RECT 1649.170 25.400 1649.490 25.460 ;
        RECT 1635.845 25.260 1649.490 25.400 ;
        RECT 1635.845 25.215 1636.135 25.260 ;
        RECT 1649.170 25.200 1649.490 25.260 ;
        RECT 1608.705 24.720 1608.995 24.765 ;
        RECT 1634.925 24.720 1635.215 24.765 ;
        RECT 1608.705 24.580 1635.215 24.720 ;
        RECT 1608.705 24.535 1608.995 24.580 ;
        RECT 1634.925 24.535 1635.215 24.580 ;
      LAYER via ;
        RECT 1649.200 1677.940 1649.460 1678.200 ;
        RECT 1650.580 1677.940 1650.840 1678.200 ;
        RECT 1221.860 25.200 1222.120 25.460 ;
        RECT 1649.200 25.200 1649.460 25.460 ;
      LAYER met2 ;
        RECT 1651.885 1700.410 1652.165 1704.000 ;
        RECT 1650.640 1700.270 1652.165 1700.410 ;
        RECT 1650.640 1678.230 1650.780 1700.270 ;
        RECT 1651.885 1700.000 1652.165 1700.270 ;
        RECT 1649.200 1677.910 1649.460 1678.230 ;
        RECT 1650.580 1677.910 1650.840 1678.230 ;
        RECT 1649.260 25.490 1649.400 1677.910 ;
        RECT 1221.860 25.170 1222.120 25.490 ;
        RECT 1649.200 25.170 1649.460 25.490 ;
        RECT 1221.920 2.400 1222.060 25.170 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1656.070 1678.140 1656.390 1678.200 ;
        RECT 1657.910 1678.140 1658.230 1678.200 ;
        RECT 1656.070 1678.000 1658.230 1678.140 ;
        RECT 1656.070 1677.940 1656.390 1678.000 ;
        RECT 1657.910 1677.940 1658.230 1678.000 ;
        RECT 1239.770 25.740 1240.090 25.800 ;
        RECT 1656.070 25.740 1656.390 25.800 ;
        RECT 1239.770 25.600 1656.390 25.740 ;
        RECT 1239.770 25.540 1240.090 25.600 ;
        RECT 1656.070 25.540 1656.390 25.600 ;
      LAYER via ;
        RECT 1656.100 1677.940 1656.360 1678.200 ;
        RECT 1657.940 1677.940 1658.200 1678.200 ;
        RECT 1239.800 25.540 1240.060 25.800 ;
        RECT 1656.100 25.540 1656.360 25.800 ;
      LAYER met2 ;
        RECT 1659.245 1700.410 1659.525 1704.000 ;
        RECT 1658.000 1700.270 1659.525 1700.410 ;
        RECT 1658.000 1678.230 1658.140 1700.270 ;
        RECT 1659.245 1700.000 1659.525 1700.270 ;
        RECT 1656.100 1677.910 1656.360 1678.230 ;
        RECT 1657.940 1677.910 1658.200 1678.230 ;
        RECT 1656.160 25.830 1656.300 1677.910 ;
        RECT 1239.800 25.510 1240.060 25.830 ;
        RECT 1656.100 25.510 1656.360 25.830 ;
        RECT 1239.860 2.400 1240.000 25.510 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1662.970 1678.140 1663.290 1678.200 ;
        RECT 1665.270 1678.140 1665.590 1678.200 ;
        RECT 1662.970 1678.000 1665.590 1678.140 ;
        RECT 1662.970 1677.940 1663.290 1678.000 ;
        RECT 1665.270 1677.940 1665.590 1678.000 ;
        RECT 1257.250 26.080 1257.570 26.140 ;
        RECT 1662.970 26.080 1663.290 26.140 ;
        RECT 1257.250 25.940 1663.290 26.080 ;
        RECT 1257.250 25.880 1257.570 25.940 ;
        RECT 1662.970 25.880 1663.290 25.940 ;
      LAYER via ;
        RECT 1663.000 1677.940 1663.260 1678.200 ;
        RECT 1665.300 1677.940 1665.560 1678.200 ;
        RECT 1257.280 25.880 1257.540 26.140 ;
        RECT 1663.000 25.880 1663.260 26.140 ;
      LAYER met2 ;
        RECT 1666.605 1700.410 1666.885 1704.000 ;
        RECT 1665.360 1700.270 1666.885 1700.410 ;
        RECT 1665.360 1678.230 1665.500 1700.270 ;
        RECT 1666.605 1700.000 1666.885 1700.270 ;
        RECT 1663.000 1677.910 1663.260 1678.230 ;
        RECT 1665.300 1677.910 1665.560 1678.230 ;
        RECT 1663.060 26.170 1663.200 1677.910 ;
        RECT 1257.280 25.850 1257.540 26.170 ;
        RECT 1663.000 25.850 1663.260 26.170 ;
        RECT 1257.340 2.400 1257.480 25.850 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1669.870 1678.140 1670.190 1678.200 ;
        RECT 1672.630 1678.140 1672.950 1678.200 ;
        RECT 1669.870 1678.000 1672.950 1678.140 ;
        RECT 1669.870 1677.940 1670.190 1678.000 ;
        RECT 1672.630 1677.940 1672.950 1678.000 ;
        RECT 1593.510 23.700 1593.830 23.760 ;
        RECT 1593.510 23.560 1616.280 23.700 ;
        RECT 1593.510 23.500 1593.830 23.560 ;
        RECT 1616.140 23.360 1616.280 23.560 ;
        RECT 1669.870 23.360 1670.190 23.420 ;
        RECT 1616.140 23.220 1670.190 23.360 ;
        RECT 1669.870 23.160 1670.190 23.220 ;
        RECT 1275.190 17.240 1275.510 17.300 ;
        RECT 1593.510 17.240 1593.830 17.300 ;
        RECT 1275.190 17.100 1593.830 17.240 ;
        RECT 1275.190 17.040 1275.510 17.100 ;
        RECT 1593.510 17.040 1593.830 17.100 ;
      LAYER via ;
        RECT 1669.900 1677.940 1670.160 1678.200 ;
        RECT 1672.660 1677.940 1672.920 1678.200 ;
        RECT 1593.540 23.500 1593.800 23.760 ;
        RECT 1669.900 23.160 1670.160 23.420 ;
        RECT 1275.220 17.040 1275.480 17.300 ;
        RECT 1593.540 17.040 1593.800 17.300 ;
      LAYER met2 ;
        RECT 1673.965 1700.410 1674.245 1704.000 ;
        RECT 1672.720 1700.270 1674.245 1700.410 ;
        RECT 1672.720 1678.230 1672.860 1700.270 ;
        RECT 1673.965 1700.000 1674.245 1700.270 ;
        RECT 1669.900 1677.910 1670.160 1678.230 ;
        RECT 1672.660 1677.910 1672.920 1678.230 ;
        RECT 1593.540 23.470 1593.800 23.790 ;
        RECT 1593.600 17.330 1593.740 23.470 ;
        RECT 1669.960 23.450 1670.100 1677.910 ;
        RECT 1669.900 23.130 1670.160 23.450 ;
        RECT 1275.220 17.010 1275.480 17.330 ;
        RECT 1593.540 17.010 1593.800 17.330 ;
        RECT 1275.280 2.400 1275.420 17.010 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1676.770 1669.640 1677.090 1669.700 ;
        RECT 1679.990 1669.640 1680.310 1669.700 ;
        RECT 1676.770 1669.500 1680.310 1669.640 ;
        RECT 1676.770 1669.440 1677.090 1669.500 ;
        RECT 1679.990 1669.440 1680.310 1669.500 ;
        RECT 1601.790 22.680 1602.110 22.740 ;
        RECT 1676.770 22.680 1677.090 22.740 ;
        RECT 1601.790 22.540 1677.090 22.680 ;
        RECT 1601.790 22.480 1602.110 22.540 ;
        RECT 1676.770 22.480 1677.090 22.540 ;
        RECT 1293.130 17.580 1293.450 17.640 ;
        RECT 1601.790 17.580 1602.110 17.640 ;
        RECT 1293.130 17.440 1602.110 17.580 ;
        RECT 1293.130 17.380 1293.450 17.440 ;
        RECT 1601.790 17.380 1602.110 17.440 ;
      LAYER via ;
        RECT 1676.800 1669.440 1677.060 1669.700 ;
        RECT 1680.020 1669.440 1680.280 1669.700 ;
        RECT 1601.820 22.480 1602.080 22.740 ;
        RECT 1676.800 22.480 1677.060 22.740 ;
        RECT 1293.160 17.380 1293.420 17.640 ;
        RECT 1601.820 17.380 1602.080 17.640 ;
      LAYER met2 ;
        RECT 1681.325 1700.410 1681.605 1704.000 ;
        RECT 1680.080 1700.270 1681.605 1700.410 ;
        RECT 1680.080 1669.730 1680.220 1700.270 ;
        RECT 1681.325 1700.000 1681.605 1700.270 ;
        RECT 1676.800 1669.410 1677.060 1669.730 ;
        RECT 1680.020 1669.410 1680.280 1669.730 ;
        RECT 1676.860 22.770 1677.000 1669.410 ;
        RECT 1601.820 22.450 1602.080 22.770 ;
        RECT 1676.800 22.450 1677.060 22.770 ;
        RECT 1601.880 17.670 1602.020 22.450 ;
        RECT 1293.160 17.350 1293.420 17.670 ;
        RECT 1601.820 17.350 1602.080 17.670 ;
        RECT 1293.220 2.400 1293.360 17.350 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1685.585 1545.385 1685.755 1559.835 ;
        RECT 1685.585 1490.645 1685.755 1538.755 ;
        RECT 1685.585 1393.745 1685.755 1441.855 ;
        RECT 1686.505 1110.865 1686.675 1126.675 ;
        RECT 1685.585 931.345 1685.755 959.055 ;
        RECT 1685.585 807.245 1685.755 855.355 ;
        RECT 1685.125 524.365 1685.295 572.475 ;
        RECT 1686.045 476.085 1686.215 523.855 ;
        RECT 1685.585 241.485 1685.755 255.595 ;
        RECT 1603.245 17.085 1603.415 18.275 ;
      LAYER mcon ;
        RECT 1685.585 1559.665 1685.755 1559.835 ;
        RECT 1685.585 1538.585 1685.755 1538.755 ;
        RECT 1685.585 1441.685 1685.755 1441.855 ;
        RECT 1686.505 1126.505 1686.675 1126.675 ;
        RECT 1685.585 958.885 1685.755 959.055 ;
        RECT 1685.585 855.185 1685.755 855.355 ;
        RECT 1685.125 572.305 1685.295 572.475 ;
        RECT 1686.045 523.685 1686.215 523.855 ;
        RECT 1685.585 255.425 1685.755 255.595 ;
        RECT 1603.245 18.105 1603.415 18.275 ;
      LAYER met1 ;
        RECT 1685.510 1559.820 1685.830 1559.880 ;
        RECT 1685.315 1559.680 1685.830 1559.820 ;
        RECT 1685.510 1559.620 1685.830 1559.680 ;
        RECT 1685.525 1545.540 1685.815 1545.585 ;
        RECT 1685.970 1545.540 1686.290 1545.600 ;
        RECT 1685.525 1545.400 1686.290 1545.540 ;
        RECT 1685.525 1545.355 1685.815 1545.400 ;
        RECT 1685.970 1545.340 1686.290 1545.400 ;
        RECT 1685.510 1538.740 1685.830 1538.800 ;
        RECT 1685.315 1538.600 1685.830 1538.740 ;
        RECT 1685.510 1538.540 1685.830 1538.600 ;
        RECT 1685.525 1490.800 1685.815 1490.845 ;
        RECT 1686.430 1490.800 1686.750 1490.860 ;
        RECT 1685.525 1490.660 1686.750 1490.800 ;
        RECT 1685.525 1490.615 1685.815 1490.660 ;
        RECT 1686.430 1490.600 1686.750 1490.660 ;
        RECT 1685.510 1452.040 1685.830 1452.100 ;
        RECT 1686.430 1452.040 1686.750 1452.100 ;
        RECT 1685.510 1451.900 1686.750 1452.040 ;
        RECT 1685.510 1451.840 1685.830 1451.900 ;
        RECT 1686.430 1451.840 1686.750 1451.900 ;
        RECT 1685.510 1441.840 1685.830 1441.900 ;
        RECT 1685.315 1441.700 1685.830 1441.840 ;
        RECT 1685.510 1441.640 1685.830 1441.700 ;
        RECT 1685.525 1393.900 1685.815 1393.945 ;
        RECT 1685.970 1393.900 1686.290 1393.960 ;
        RECT 1685.525 1393.760 1686.290 1393.900 ;
        RECT 1685.525 1393.715 1685.815 1393.760 ;
        RECT 1685.970 1393.700 1686.290 1393.760 ;
        RECT 1685.970 1366.700 1686.290 1366.760 ;
        RECT 1685.600 1366.560 1686.290 1366.700 ;
        RECT 1685.600 1366.080 1685.740 1366.560 ;
        RECT 1685.970 1366.500 1686.290 1366.560 ;
        RECT 1685.510 1365.820 1685.830 1366.080 ;
        RECT 1685.510 1297.340 1685.830 1297.400 ;
        RECT 1686.430 1297.340 1686.750 1297.400 ;
        RECT 1685.510 1297.200 1686.750 1297.340 ;
        RECT 1685.510 1297.140 1685.830 1297.200 ;
        RECT 1686.430 1297.140 1686.750 1297.200 ;
        RECT 1685.510 1269.600 1685.830 1269.860 ;
        RECT 1685.600 1269.120 1685.740 1269.600 ;
        RECT 1686.430 1269.120 1686.750 1269.180 ;
        RECT 1685.600 1268.980 1686.750 1269.120 ;
        RECT 1686.430 1268.920 1686.750 1268.980 ;
        RECT 1686.430 1126.660 1686.750 1126.720 ;
        RECT 1686.235 1126.520 1686.750 1126.660 ;
        RECT 1686.430 1126.460 1686.750 1126.520 ;
        RECT 1686.430 1111.020 1686.750 1111.080 ;
        RECT 1686.235 1110.880 1686.750 1111.020 ;
        RECT 1686.430 1110.820 1686.750 1110.880 ;
        RECT 1685.970 1014.460 1686.290 1014.520 ;
        RECT 1686.430 1014.460 1686.750 1014.520 ;
        RECT 1685.970 1014.320 1686.750 1014.460 ;
        RECT 1685.970 1014.260 1686.290 1014.320 ;
        RECT 1686.430 1014.260 1686.750 1014.320 ;
        RECT 1685.970 980.460 1686.290 980.520 ;
        RECT 1685.600 980.320 1686.290 980.460 ;
        RECT 1685.600 979.840 1685.740 980.320 ;
        RECT 1685.970 980.260 1686.290 980.320 ;
        RECT 1685.510 979.580 1685.830 979.840 ;
        RECT 1685.510 959.040 1685.830 959.100 ;
        RECT 1685.315 958.900 1685.830 959.040 ;
        RECT 1685.510 958.840 1685.830 958.900 ;
        RECT 1685.510 931.500 1685.830 931.560 ;
        RECT 1685.315 931.360 1685.830 931.500 ;
        RECT 1685.510 931.300 1685.830 931.360 ;
        RECT 1685.510 862.620 1685.830 862.880 ;
        RECT 1685.600 862.200 1685.740 862.620 ;
        RECT 1685.510 861.940 1685.830 862.200 ;
        RECT 1685.510 855.340 1685.830 855.400 ;
        RECT 1685.315 855.200 1685.830 855.340 ;
        RECT 1685.510 855.140 1685.830 855.200 ;
        RECT 1685.525 807.400 1685.815 807.445 ;
        RECT 1686.430 807.400 1686.750 807.460 ;
        RECT 1685.525 807.260 1686.750 807.400 ;
        RECT 1685.525 807.215 1685.815 807.260 ;
        RECT 1686.430 807.200 1686.750 807.260 ;
        RECT 1686.430 766.260 1686.750 766.320 ;
        RECT 1686.060 766.120 1686.750 766.260 ;
        RECT 1686.060 765.980 1686.200 766.120 ;
        RECT 1686.430 766.060 1686.750 766.120 ;
        RECT 1685.970 765.720 1686.290 765.980 ;
        RECT 1685.510 676.160 1685.830 676.220 ;
        RECT 1685.970 676.160 1686.290 676.220 ;
        RECT 1685.510 676.020 1686.290 676.160 ;
        RECT 1685.510 675.960 1685.830 676.020 ;
        RECT 1685.970 675.960 1686.290 676.020 ;
        RECT 1685.510 627.880 1685.830 627.940 ;
        RECT 1686.430 627.880 1686.750 627.940 ;
        RECT 1685.510 627.740 1686.750 627.880 ;
        RECT 1685.510 627.680 1685.830 627.740 ;
        RECT 1686.430 627.680 1686.750 627.740 ;
        RECT 1685.065 572.460 1685.355 572.505 ;
        RECT 1685.970 572.460 1686.290 572.520 ;
        RECT 1685.065 572.320 1686.290 572.460 ;
        RECT 1685.065 572.275 1685.355 572.320 ;
        RECT 1685.970 572.260 1686.290 572.320 ;
        RECT 1685.050 524.520 1685.370 524.580 ;
        RECT 1684.855 524.380 1685.370 524.520 ;
        RECT 1685.050 524.320 1685.370 524.380 ;
        RECT 1685.050 523.840 1685.370 523.900 ;
        RECT 1685.985 523.840 1686.275 523.885 ;
        RECT 1685.050 523.700 1686.275 523.840 ;
        RECT 1685.050 523.640 1685.370 523.700 ;
        RECT 1685.985 523.655 1686.275 523.700 ;
        RECT 1685.970 476.240 1686.290 476.300 ;
        RECT 1685.775 476.100 1686.290 476.240 ;
        RECT 1685.970 476.040 1686.290 476.100 ;
        RECT 1685.970 304.000 1686.290 304.260 ;
        RECT 1686.060 303.240 1686.200 304.000 ;
        RECT 1685.970 302.980 1686.290 303.240 ;
        RECT 1685.525 255.580 1685.815 255.625 ;
        RECT 1685.970 255.580 1686.290 255.640 ;
        RECT 1685.525 255.440 1686.290 255.580 ;
        RECT 1685.525 255.395 1685.815 255.440 ;
        RECT 1685.970 255.380 1686.290 255.440 ;
        RECT 1685.510 241.640 1685.830 241.700 ;
        RECT 1685.315 241.500 1685.830 241.640 ;
        RECT 1685.510 241.440 1685.830 241.500 ;
        RECT 1613.750 23.020 1614.070 23.080 ;
        RECT 1685.970 23.020 1686.290 23.080 ;
        RECT 1613.750 22.880 1686.290 23.020 ;
        RECT 1613.750 22.820 1614.070 22.880 ;
        RECT 1685.970 22.820 1686.290 22.880 ;
        RECT 1311.070 18.260 1311.390 18.320 ;
        RECT 1603.185 18.260 1603.475 18.305 ;
        RECT 1311.070 18.120 1603.475 18.260 ;
        RECT 1311.070 18.060 1311.390 18.120 ;
        RECT 1603.185 18.075 1603.475 18.120 ;
        RECT 1603.185 17.240 1603.475 17.285 ;
        RECT 1613.750 17.240 1614.070 17.300 ;
        RECT 1603.185 17.100 1614.070 17.240 ;
        RECT 1603.185 17.055 1603.475 17.100 ;
        RECT 1613.750 17.040 1614.070 17.100 ;
      LAYER via ;
        RECT 1685.540 1559.620 1685.800 1559.880 ;
        RECT 1686.000 1545.340 1686.260 1545.600 ;
        RECT 1685.540 1538.540 1685.800 1538.800 ;
        RECT 1686.460 1490.600 1686.720 1490.860 ;
        RECT 1685.540 1451.840 1685.800 1452.100 ;
        RECT 1686.460 1451.840 1686.720 1452.100 ;
        RECT 1685.540 1441.640 1685.800 1441.900 ;
        RECT 1686.000 1393.700 1686.260 1393.960 ;
        RECT 1686.000 1366.500 1686.260 1366.760 ;
        RECT 1685.540 1365.820 1685.800 1366.080 ;
        RECT 1685.540 1297.140 1685.800 1297.400 ;
        RECT 1686.460 1297.140 1686.720 1297.400 ;
        RECT 1685.540 1269.600 1685.800 1269.860 ;
        RECT 1686.460 1268.920 1686.720 1269.180 ;
        RECT 1686.460 1126.460 1686.720 1126.720 ;
        RECT 1686.460 1110.820 1686.720 1111.080 ;
        RECT 1686.000 1014.260 1686.260 1014.520 ;
        RECT 1686.460 1014.260 1686.720 1014.520 ;
        RECT 1686.000 980.260 1686.260 980.520 ;
        RECT 1685.540 979.580 1685.800 979.840 ;
        RECT 1685.540 958.840 1685.800 959.100 ;
        RECT 1685.540 931.300 1685.800 931.560 ;
        RECT 1685.540 862.620 1685.800 862.880 ;
        RECT 1685.540 861.940 1685.800 862.200 ;
        RECT 1685.540 855.140 1685.800 855.400 ;
        RECT 1686.460 807.200 1686.720 807.460 ;
        RECT 1686.460 766.060 1686.720 766.320 ;
        RECT 1686.000 765.720 1686.260 765.980 ;
        RECT 1685.540 675.960 1685.800 676.220 ;
        RECT 1686.000 675.960 1686.260 676.220 ;
        RECT 1685.540 627.680 1685.800 627.940 ;
        RECT 1686.460 627.680 1686.720 627.940 ;
        RECT 1686.000 572.260 1686.260 572.520 ;
        RECT 1685.080 524.320 1685.340 524.580 ;
        RECT 1685.080 523.640 1685.340 523.900 ;
        RECT 1686.000 476.040 1686.260 476.300 ;
        RECT 1686.000 304.000 1686.260 304.260 ;
        RECT 1686.000 302.980 1686.260 303.240 ;
        RECT 1686.000 255.380 1686.260 255.640 ;
        RECT 1685.540 241.440 1685.800 241.700 ;
        RECT 1613.780 22.820 1614.040 23.080 ;
        RECT 1686.000 22.820 1686.260 23.080 ;
        RECT 1311.100 18.060 1311.360 18.320 ;
        RECT 1613.780 17.040 1614.040 17.300 ;
      LAYER met2 ;
        RECT 1688.685 1701.090 1688.965 1704.000 ;
        RECT 1686.980 1700.950 1688.965 1701.090 ;
        RECT 1686.980 1677.970 1687.120 1700.950 ;
        RECT 1688.685 1700.000 1688.965 1700.950 ;
        RECT 1685.600 1677.830 1687.120 1677.970 ;
        RECT 1685.600 1656.040 1685.740 1677.830 ;
        RECT 1685.600 1655.900 1686.200 1656.040 ;
        RECT 1686.060 1595.125 1686.200 1655.900 ;
        RECT 1685.990 1594.755 1686.270 1595.125 ;
        RECT 1685.530 1594.075 1685.810 1594.445 ;
        RECT 1685.600 1559.910 1685.740 1594.075 ;
        RECT 1685.540 1559.590 1685.800 1559.910 ;
        RECT 1686.000 1545.310 1686.260 1545.630 ;
        RECT 1686.060 1539.250 1686.200 1545.310 ;
        RECT 1685.600 1539.110 1686.200 1539.250 ;
        RECT 1685.600 1538.830 1685.740 1539.110 ;
        RECT 1685.540 1538.510 1685.800 1538.830 ;
        RECT 1686.460 1490.570 1686.720 1490.890 ;
        RECT 1686.520 1452.130 1686.660 1490.570 ;
        RECT 1685.540 1451.810 1685.800 1452.130 ;
        RECT 1686.460 1451.810 1686.720 1452.130 ;
        RECT 1685.600 1441.930 1685.740 1451.810 ;
        RECT 1685.540 1441.610 1685.800 1441.930 ;
        RECT 1686.000 1393.670 1686.260 1393.990 ;
        RECT 1686.060 1366.790 1686.200 1393.670 ;
        RECT 1686.000 1366.470 1686.260 1366.790 ;
        RECT 1685.540 1365.790 1685.800 1366.110 ;
        RECT 1685.600 1345.565 1685.740 1365.790 ;
        RECT 1685.530 1345.195 1685.810 1345.565 ;
        RECT 1686.450 1345.195 1686.730 1345.565 ;
        RECT 1686.520 1297.430 1686.660 1345.195 ;
        RECT 1685.540 1297.110 1685.800 1297.430 ;
        RECT 1686.460 1297.110 1686.720 1297.430 ;
        RECT 1685.600 1269.890 1685.740 1297.110 ;
        RECT 1685.540 1269.570 1685.800 1269.890 ;
        RECT 1686.460 1268.890 1686.720 1269.210 ;
        RECT 1686.520 1200.725 1686.660 1268.890 ;
        RECT 1685.530 1200.355 1685.810 1200.725 ;
        RECT 1686.450 1200.355 1686.730 1200.725 ;
        RECT 1685.600 1157.770 1685.740 1200.355 ;
        RECT 1685.600 1157.630 1686.660 1157.770 ;
        RECT 1686.520 1126.750 1686.660 1157.630 ;
        RECT 1686.460 1126.430 1686.720 1126.750 ;
        RECT 1686.460 1110.790 1686.720 1111.110 ;
        RECT 1686.520 1104.165 1686.660 1110.790 ;
        RECT 1685.530 1103.795 1685.810 1104.165 ;
        RECT 1686.450 1103.795 1686.730 1104.165 ;
        RECT 1685.600 1061.210 1685.740 1103.795 ;
        RECT 1685.600 1061.070 1686.660 1061.210 ;
        RECT 1686.520 1014.550 1686.660 1061.070 ;
        RECT 1686.000 1014.230 1686.260 1014.550 ;
        RECT 1686.460 1014.230 1686.720 1014.550 ;
        RECT 1686.060 980.550 1686.200 1014.230 ;
        RECT 1686.000 980.230 1686.260 980.550 ;
        RECT 1685.540 979.550 1685.800 979.870 ;
        RECT 1685.600 959.130 1685.740 979.550 ;
        RECT 1685.540 958.810 1685.800 959.130 ;
        RECT 1685.540 931.270 1685.800 931.590 ;
        RECT 1685.600 862.910 1685.740 931.270 ;
        RECT 1685.540 862.590 1685.800 862.910 ;
        RECT 1685.540 861.910 1685.800 862.230 ;
        RECT 1685.600 855.430 1685.740 861.910 ;
        RECT 1685.540 855.110 1685.800 855.430 ;
        RECT 1686.460 807.170 1686.720 807.490 ;
        RECT 1686.520 766.350 1686.660 807.170 ;
        RECT 1686.460 766.030 1686.720 766.350 ;
        RECT 1686.000 765.690 1686.260 766.010 ;
        RECT 1686.060 677.125 1686.200 765.690 ;
        RECT 1685.990 676.755 1686.270 677.125 ;
        RECT 1685.540 675.930 1685.800 676.250 ;
        RECT 1685.990 676.075 1686.270 676.445 ;
        RECT 1686.000 675.930 1686.260 676.075 ;
        RECT 1685.600 627.970 1685.740 675.930 ;
        RECT 1685.540 627.650 1685.800 627.970 ;
        RECT 1686.460 627.650 1686.720 627.970 ;
        RECT 1686.520 602.890 1686.660 627.650 ;
        RECT 1686.060 602.750 1686.660 602.890 ;
        RECT 1686.060 572.550 1686.200 602.750 ;
        RECT 1686.000 572.230 1686.260 572.550 ;
        RECT 1685.080 524.290 1685.340 524.610 ;
        RECT 1685.140 523.930 1685.280 524.290 ;
        RECT 1685.080 523.610 1685.340 523.930 ;
        RECT 1686.000 476.010 1686.260 476.330 ;
        RECT 1686.060 402.290 1686.200 476.010 ;
        RECT 1686.060 402.150 1686.660 402.290 ;
        RECT 1686.520 400.930 1686.660 402.150 ;
        RECT 1686.060 400.790 1686.660 400.930 ;
        RECT 1686.060 304.290 1686.200 400.790 ;
        RECT 1686.000 303.970 1686.260 304.290 ;
        RECT 1686.000 302.950 1686.260 303.270 ;
        RECT 1686.060 255.670 1686.200 302.950 ;
        RECT 1686.000 255.350 1686.260 255.670 ;
        RECT 1685.540 241.410 1685.800 241.730 ;
        RECT 1685.600 217.330 1685.740 241.410 ;
        RECT 1685.600 217.190 1686.200 217.330 ;
        RECT 1686.060 110.570 1686.200 217.190 ;
        RECT 1685.600 110.430 1686.200 110.570 ;
        RECT 1685.600 72.490 1685.740 110.430 ;
        RECT 1685.600 72.350 1686.200 72.490 ;
        RECT 1686.060 23.110 1686.200 72.350 ;
        RECT 1613.780 22.790 1614.040 23.110 ;
        RECT 1686.000 22.790 1686.260 23.110 ;
        RECT 1311.100 18.030 1311.360 18.350 ;
        RECT 1311.160 2.400 1311.300 18.030 ;
        RECT 1613.840 17.330 1613.980 22.790 ;
        RECT 1613.780 17.010 1614.040 17.330 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
      LAYER via2 ;
        RECT 1685.990 1594.800 1686.270 1595.080 ;
        RECT 1685.530 1594.120 1685.810 1594.400 ;
        RECT 1685.530 1345.240 1685.810 1345.520 ;
        RECT 1686.450 1345.240 1686.730 1345.520 ;
        RECT 1685.530 1200.400 1685.810 1200.680 ;
        RECT 1686.450 1200.400 1686.730 1200.680 ;
        RECT 1685.530 1103.840 1685.810 1104.120 ;
        RECT 1686.450 1103.840 1686.730 1104.120 ;
        RECT 1685.990 676.800 1686.270 677.080 ;
        RECT 1685.990 676.120 1686.270 676.400 ;
      LAYER met3 ;
        RECT 1685.965 1595.090 1686.295 1595.105 ;
        RECT 1684.830 1594.790 1686.295 1595.090 ;
        RECT 1684.830 1594.410 1685.130 1594.790 ;
        RECT 1685.965 1594.775 1686.295 1594.790 ;
        RECT 1685.505 1594.410 1685.835 1594.425 ;
        RECT 1684.830 1594.110 1685.835 1594.410 ;
        RECT 1685.505 1594.095 1685.835 1594.110 ;
        RECT 1685.505 1345.530 1685.835 1345.545 ;
        RECT 1686.425 1345.530 1686.755 1345.545 ;
        RECT 1685.505 1345.230 1686.755 1345.530 ;
        RECT 1685.505 1345.215 1685.835 1345.230 ;
        RECT 1686.425 1345.215 1686.755 1345.230 ;
        RECT 1685.505 1200.690 1685.835 1200.705 ;
        RECT 1686.425 1200.690 1686.755 1200.705 ;
        RECT 1685.505 1200.390 1686.755 1200.690 ;
        RECT 1685.505 1200.375 1685.835 1200.390 ;
        RECT 1686.425 1200.375 1686.755 1200.390 ;
        RECT 1685.505 1104.130 1685.835 1104.145 ;
        RECT 1686.425 1104.130 1686.755 1104.145 ;
        RECT 1685.505 1103.830 1686.755 1104.130 ;
        RECT 1685.505 1103.815 1685.835 1103.830 ;
        RECT 1686.425 1103.815 1686.755 1103.830 ;
        RECT 1685.965 677.090 1686.295 677.105 ;
        RECT 1685.965 676.790 1686.970 677.090 ;
        RECT 1685.965 676.775 1686.295 676.790 ;
        RECT 1685.965 676.410 1686.295 676.425 ;
        RECT 1686.670 676.410 1686.970 676.790 ;
        RECT 1685.965 676.110 1686.970 676.410 ;
        RECT 1685.965 676.095 1686.295 676.110 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1690.570 1678.140 1690.890 1678.200 ;
        RECT 1694.710 1678.140 1695.030 1678.200 ;
        RECT 1690.570 1678.000 1695.030 1678.140 ;
        RECT 1690.570 1677.940 1690.890 1678.000 ;
        RECT 1694.710 1677.940 1695.030 1678.000 ;
        RECT 1625.710 22.340 1626.030 22.400 ;
        RECT 1690.570 22.340 1690.890 22.400 ;
        RECT 1625.710 22.200 1690.890 22.340 ;
        RECT 1625.710 22.140 1626.030 22.200 ;
        RECT 1690.570 22.140 1690.890 22.200 ;
        RECT 1625.710 18.260 1626.030 18.320 ;
        RECT 1603.720 18.120 1626.030 18.260 ;
        RECT 1329.010 17.920 1329.330 17.980 ;
        RECT 1603.720 17.920 1603.860 18.120 ;
        RECT 1625.710 18.060 1626.030 18.120 ;
        RECT 1329.010 17.780 1603.860 17.920 ;
        RECT 1329.010 17.720 1329.330 17.780 ;
      LAYER via ;
        RECT 1690.600 1677.940 1690.860 1678.200 ;
        RECT 1694.740 1677.940 1695.000 1678.200 ;
        RECT 1625.740 22.140 1626.000 22.400 ;
        RECT 1690.600 22.140 1690.860 22.400 ;
        RECT 1329.040 17.720 1329.300 17.980 ;
        RECT 1625.740 18.060 1626.000 18.320 ;
      LAYER met2 ;
        RECT 1696.045 1700.410 1696.325 1704.000 ;
        RECT 1694.800 1700.270 1696.325 1700.410 ;
        RECT 1694.800 1678.230 1694.940 1700.270 ;
        RECT 1696.045 1700.000 1696.325 1700.270 ;
        RECT 1690.600 1677.910 1690.860 1678.230 ;
        RECT 1694.740 1677.910 1695.000 1678.230 ;
        RECT 1690.660 22.430 1690.800 1677.910 ;
        RECT 1625.740 22.110 1626.000 22.430 ;
        RECT 1690.600 22.110 1690.860 22.430 ;
        RECT 1625.800 18.350 1625.940 22.110 ;
        RECT 1625.740 18.030 1626.000 18.350 ;
        RECT 1329.040 17.690 1329.300 18.010 ;
        RECT 1329.100 2.400 1329.240 17.690 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1428.370 1678.140 1428.690 1678.200 ;
        RECT 1429.750 1678.140 1430.070 1678.200 ;
        RECT 1428.370 1678.000 1430.070 1678.140 ;
        RECT 1428.370 1677.940 1428.690 1678.000 ;
        RECT 1429.750 1677.940 1430.070 1678.000 ;
        RECT 686.390 27.440 686.710 27.500 ;
        RECT 1428.370 27.440 1428.690 27.500 ;
        RECT 686.390 27.300 1428.690 27.440 ;
        RECT 686.390 27.240 686.710 27.300 ;
        RECT 1428.370 27.240 1428.690 27.300 ;
      LAYER via ;
        RECT 1428.400 1677.940 1428.660 1678.200 ;
        RECT 1429.780 1677.940 1430.040 1678.200 ;
        RECT 686.420 27.240 686.680 27.500 ;
        RECT 1428.400 27.240 1428.660 27.500 ;
      LAYER met2 ;
        RECT 1431.545 1700.410 1431.825 1704.000 ;
        RECT 1429.840 1700.270 1431.825 1700.410 ;
        RECT 1429.840 1678.230 1429.980 1700.270 ;
        RECT 1431.545 1700.000 1431.825 1700.270 ;
        RECT 1428.400 1677.910 1428.660 1678.230 ;
        RECT 1429.780 1677.910 1430.040 1678.230 ;
        RECT 1428.460 27.530 1428.600 1677.910 ;
        RECT 686.420 27.210 686.680 27.530 ;
        RECT 1428.400 27.210 1428.660 27.530 ;
        RECT 686.480 2.400 686.620 27.210 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1698.925 621.265 1699.095 676.175 ;
        RECT 1698.925 589.985 1699.095 613.955 ;
        RECT 1698.925 282.965 1699.095 304.215 ;
        RECT 1698.925 210.205 1699.095 234.515 ;
        RECT 1698.465 144.925 1698.635 159.035 ;
        RECT 1698.465 48.365 1698.635 96.135 ;
        RECT 1366.345 15.045 1366.515 16.235 ;
        RECT 1414.185 15.045 1414.355 16.915 ;
      LAYER mcon ;
        RECT 1698.925 676.005 1699.095 676.175 ;
        RECT 1698.925 613.785 1699.095 613.955 ;
        RECT 1698.925 304.045 1699.095 304.215 ;
        RECT 1698.925 234.345 1699.095 234.515 ;
        RECT 1698.465 158.865 1698.635 159.035 ;
        RECT 1698.465 95.965 1698.635 96.135 ;
        RECT 1414.185 16.745 1414.355 16.915 ;
        RECT 1366.345 16.065 1366.515 16.235 ;
      LAYER met1 ;
        RECT 1698.850 1642.440 1699.170 1642.500 ;
        RECT 1701.610 1642.440 1701.930 1642.500 ;
        RECT 1698.850 1642.300 1701.930 1642.440 ;
        RECT 1698.850 1642.240 1699.170 1642.300 ;
        RECT 1701.610 1642.240 1701.930 1642.300 ;
        RECT 1698.850 934.900 1699.170 934.960 ;
        RECT 1699.770 934.900 1700.090 934.960 ;
        RECT 1698.850 934.760 1700.090 934.900 ;
        RECT 1698.850 934.700 1699.170 934.760 ;
        RECT 1699.770 934.700 1700.090 934.760 ;
        RECT 1698.850 676.160 1699.170 676.220 ;
        RECT 1698.655 676.020 1699.170 676.160 ;
        RECT 1698.850 675.960 1699.170 676.020 ;
        RECT 1698.390 621.420 1698.710 621.480 ;
        RECT 1698.865 621.420 1699.155 621.465 ;
        RECT 1698.390 621.280 1699.155 621.420 ;
        RECT 1698.390 621.220 1698.710 621.280 ;
        RECT 1698.865 621.235 1699.155 621.280 ;
        RECT 1698.850 613.940 1699.170 614.000 ;
        RECT 1698.655 613.800 1699.170 613.940 ;
        RECT 1698.850 613.740 1699.170 613.800 ;
        RECT 1698.850 590.140 1699.170 590.200 ;
        RECT 1698.655 590.000 1699.170 590.140 ;
        RECT 1698.850 589.940 1699.170 590.000 ;
        RECT 1698.850 400.560 1699.170 400.820 ;
        RECT 1698.940 400.140 1699.080 400.560 ;
        RECT 1698.850 399.880 1699.170 400.140 ;
        RECT 1698.850 304.200 1699.170 304.260 ;
        RECT 1698.655 304.060 1699.170 304.200 ;
        RECT 1698.850 304.000 1699.170 304.060 ;
        RECT 1698.850 283.120 1699.170 283.180 ;
        RECT 1698.655 282.980 1699.170 283.120 ;
        RECT 1698.850 282.920 1699.170 282.980 ;
        RECT 1698.850 234.500 1699.170 234.560 ;
        RECT 1698.655 234.360 1699.170 234.500 ;
        RECT 1698.850 234.300 1699.170 234.360 ;
        RECT 1698.850 210.360 1699.170 210.420 ;
        RECT 1698.655 210.220 1699.170 210.360 ;
        RECT 1698.850 210.160 1699.170 210.220 ;
        RECT 1698.405 159.020 1698.695 159.065 ;
        RECT 1698.850 159.020 1699.170 159.080 ;
        RECT 1698.405 158.880 1699.170 159.020 ;
        RECT 1698.405 158.835 1698.695 158.880 ;
        RECT 1698.850 158.820 1699.170 158.880 ;
        RECT 1698.390 145.080 1698.710 145.140 ;
        RECT 1698.195 144.940 1698.710 145.080 ;
        RECT 1698.390 144.880 1698.710 144.940 ;
        RECT 1698.390 96.800 1698.710 96.860 ;
        RECT 1698.850 96.800 1699.170 96.860 ;
        RECT 1698.390 96.660 1699.170 96.800 ;
        RECT 1698.390 96.600 1698.710 96.660 ;
        RECT 1698.850 96.600 1699.170 96.660 ;
        RECT 1698.405 96.120 1698.695 96.165 ;
        RECT 1698.850 96.120 1699.170 96.180 ;
        RECT 1698.405 95.980 1699.170 96.120 ;
        RECT 1698.405 95.935 1698.695 95.980 ;
        RECT 1698.850 95.920 1699.170 95.980 ;
        RECT 1698.390 48.520 1698.710 48.580 ;
        RECT 1698.195 48.380 1698.710 48.520 ;
        RECT 1698.390 48.320 1698.710 48.380 ;
        RECT 1449.070 32.540 1449.390 32.600 ;
        RECT 1698.390 32.540 1698.710 32.600 ;
        RECT 1449.070 32.400 1698.710 32.540 ;
        RECT 1449.070 32.340 1449.390 32.400 ;
        RECT 1698.390 32.340 1698.710 32.400 ;
        RECT 1414.125 16.900 1414.415 16.945 ;
        RECT 1449.070 16.900 1449.390 16.960 ;
        RECT 1414.125 16.760 1449.390 16.900 ;
        RECT 1414.125 16.715 1414.415 16.760 ;
        RECT 1449.070 16.700 1449.390 16.760 ;
        RECT 1346.490 16.220 1346.810 16.280 ;
        RECT 1366.285 16.220 1366.575 16.265 ;
        RECT 1346.490 16.080 1366.575 16.220 ;
        RECT 1346.490 16.020 1346.810 16.080 ;
        RECT 1366.285 16.035 1366.575 16.080 ;
        RECT 1366.285 15.200 1366.575 15.245 ;
        RECT 1414.125 15.200 1414.415 15.245 ;
        RECT 1366.285 15.060 1414.415 15.200 ;
        RECT 1366.285 15.015 1366.575 15.060 ;
        RECT 1414.125 15.015 1414.415 15.060 ;
      LAYER via ;
        RECT 1698.880 1642.240 1699.140 1642.500 ;
        RECT 1701.640 1642.240 1701.900 1642.500 ;
        RECT 1698.880 934.700 1699.140 934.960 ;
        RECT 1699.800 934.700 1700.060 934.960 ;
        RECT 1698.880 675.960 1699.140 676.220 ;
        RECT 1698.420 621.220 1698.680 621.480 ;
        RECT 1698.880 613.740 1699.140 614.000 ;
        RECT 1698.880 589.940 1699.140 590.200 ;
        RECT 1698.880 400.560 1699.140 400.820 ;
        RECT 1698.880 399.880 1699.140 400.140 ;
        RECT 1698.880 304.000 1699.140 304.260 ;
        RECT 1698.880 282.920 1699.140 283.180 ;
        RECT 1698.880 234.300 1699.140 234.560 ;
        RECT 1698.880 210.160 1699.140 210.420 ;
        RECT 1698.880 158.820 1699.140 159.080 ;
        RECT 1698.420 144.880 1698.680 145.140 ;
        RECT 1698.420 96.600 1698.680 96.860 ;
        RECT 1698.880 96.600 1699.140 96.860 ;
        RECT 1698.880 95.920 1699.140 96.180 ;
        RECT 1698.420 48.320 1698.680 48.580 ;
        RECT 1449.100 32.340 1449.360 32.600 ;
        RECT 1698.420 32.340 1698.680 32.600 ;
        RECT 1449.100 16.700 1449.360 16.960 ;
        RECT 1346.520 16.020 1346.780 16.280 ;
      LAYER met2 ;
        RECT 1703.405 1701.090 1703.685 1704.000 ;
        RECT 1701.700 1700.950 1703.685 1701.090 ;
        RECT 1701.700 1642.530 1701.840 1700.950 ;
        RECT 1703.405 1700.000 1703.685 1700.950 ;
        RECT 1698.880 1642.210 1699.140 1642.530 ;
        RECT 1701.640 1642.210 1701.900 1642.530 ;
        RECT 1698.940 1559.650 1699.080 1642.210 ;
        RECT 1698.480 1559.510 1699.080 1559.650 ;
        RECT 1698.480 1558.970 1698.620 1559.510 ;
        RECT 1698.480 1558.830 1699.080 1558.970 ;
        RECT 1698.940 1414.810 1699.080 1558.830 ;
        RECT 1698.480 1414.670 1699.080 1414.810 ;
        RECT 1698.480 1414.130 1698.620 1414.670 ;
        RECT 1698.480 1413.990 1699.080 1414.130 ;
        RECT 1698.940 1318.250 1699.080 1413.990 ;
        RECT 1698.480 1318.110 1699.080 1318.250 ;
        RECT 1698.480 1317.570 1698.620 1318.110 ;
        RECT 1698.480 1317.430 1699.080 1317.570 ;
        RECT 1698.940 1221.690 1699.080 1317.430 ;
        RECT 1698.480 1221.550 1699.080 1221.690 ;
        RECT 1698.480 1221.010 1698.620 1221.550 ;
        RECT 1698.480 1220.870 1699.080 1221.010 ;
        RECT 1698.940 1125.130 1699.080 1220.870 ;
        RECT 1698.480 1124.990 1699.080 1125.130 ;
        RECT 1698.480 1124.450 1698.620 1124.990 ;
        RECT 1698.480 1124.310 1699.080 1124.450 ;
        RECT 1698.940 1028.570 1699.080 1124.310 ;
        RECT 1698.480 1028.430 1699.080 1028.570 ;
        RECT 1698.480 1027.890 1698.620 1028.430 ;
        RECT 1698.480 1027.750 1699.080 1027.890 ;
        RECT 1698.940 934.990 1699.080 1027.750 ;
        RECT 1698.880 934.670 1699.140 934.990 ;
        RECT 1699.800 934.670 1700.060 934.990 ;
        RECT 1699.860 911.045 1700.000 934.670 ;
        RECT 1698.870 910.675 1699.150 911.045 ;
        RECT 1699.790 910.675 1700.070 911.045 ;
        RECT 1698.940 862.650 1699.080 910.675 ;
        RECT 1698.480 862.510 1699.080 862.650 ;
        RECT 1698.480 845.650 1698.620 862.510 ;
        RECT 1698.480 845.510 1699.540 845.650 ;
        RECT 1699.400 786.490 1699.540 845.510 ;
        RECT 1698.940 786.350 1699.540 786.490 ;
        RECT 1698.940 690.610 1699.080 786.350 ;
        RECT 1698.480 690.470 1699.080 690.610 ;
        RECT 1698.480 689.930 1698.620 690.470 ;
        RECT 1698.480 689.790 1699.080 689.930 ;
        RECT 1698.940 676.250 1699.080 689.790 ;
        RECT 1698.880 675.930 1699.140 676.250 ;
        RECT 1698.420 621.250 1698.680 621.510 ;
        RECT 1698.420 621.190 1699.080 621.250 ;
        RECT 1698.480 621.110 1699.080 621.190 ;
        RECT 1698.940 614.030 1699.080 621.110 ;
        RECT 1698.880 613.710 1699.140 614.030 ;
        RECT 1698.880 589.910 1699.140 590.230 ;
        RECT 1698.940 400.850 1699.080 589.910 ;
        RECT 1698.880 400.530 1699.140 400.850 ;
        RECT 1698.880 399.850 1699.140 400.170 ;
        RECT 1698.940 304.290 1699.080 399.850 ;
        RECT 1698.880 303.970 1699.140 304.290 ;
        RECT 1698.880 282.890 1699.140 283.210 ;
        RECT 1698.940 234.590 1699.080 282.890 ;
        RECT 1698.880 234.270 1699.140 234.590 ;
        RECT 1698.880 210.130 1699.140 210.450 ;
        RECT 1698.940 159.110 1699.080 210.130 ;
        RECT 1698.880 158.790 1699.140 159.110 ;
        RECT 1698.420 144.850 1698.680 145.170 ;
        RECT 1698.480 96.890 1698.620 144.850 ;
        RECT 1698.420 96.570 1698.680 96.890 ;
        RECT 1698.880 96.570 1699.140 96.890 ;
        RECT 1698.940 96.210 1699.080 96.570 ;
        RECT 1698.880 95.890 1699.140 96.210 ;
        RECT 1698.420 48.290 1698.680 48.610 ;
        RECT 1698.480 32.630 1698.620 48.290 ;
        RECT 1449.100 32.310 1449.360 32.630 ;
        RECT 1698.420 32.310 1698.680 32.630 ;
        RECT 1449.160 16.990 1449.300 32.310 ;
        RECT 1449.100 16.670 1449.360 16.990 ;
        RECT 1346.520 15.990 1346.780 16.310 ;
        RECT 1346.580 2.400 1346.720 15.990 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
      LAYER via2 ;
        RECT 1698.870 910.720 1699.150 911.000 ;
        RECT 1699.790 910.720 1700.070 911.000 ;
      LAYER met3 ;
        RECT 1698.845 911.010 1699.175 911.025 ;
        RECT 1699.765 911.010 1700.095 911.025 ;
        RECT 1698.845 910.710 1700.095 911.010 ;
        RECT 1698.845 910.695 1699.175 910.710 ;
        RECT 1699.765 910.695 1700.095 910.710 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1706.745 1594.005 1706.915 1642.115 ;
        RECT 1705.825 1497.445 1705.995 1545.555 ;
        RECT 1705.825 1400.885 1705.995 1448.995 ;
        RECT 1705.825 1304.325 1705.995 1352.435 ;
        RECT 1705.825 1076.185 1705.995 1103.895 ;
        RECT 1706.745 641.325 1706.915 693.515 ;
        RECT 1705.825 531.505 1705.995 579.615 ;
        RECT 1705.365 386.325 1705.535 434.775 ;
        RECT 1705.365 351.305 1705.535 385.815 ;
        RECT 1706.745 253.045 1706.915 282.795 ;
      LAYER mcon ;
        RECT 1706.745 1641.945 1706.915 1642.115 ;
        RECT 1705.825 1545.385 1705.995 1545.555 ;
        RECT 1705.825 1448.825 1705.995 1448.995 ;
        RECT 1705.825 1352.265 1705.995 1352.435 ;
        RECT 1705.825 1103.725 1705.995 1103.895 ;
        RECT 1706.745 693.345 1706.915 693.515 ;
        RECT 1705.825 579.445 1705.995 579.615 ;
        RECT 1705.365 434.605 1705.535 434.775 ;
        RECT 1705.365 385.645 1705.535 385.815 ;
        RECT 1706.745 282.625 1706.915 282.795 ;
      LAYER met1 ;
        RECT 1707.130 1656.720 1707.450 1656.780 ;
        RECT 1708.510 1656.720 1708.830 1656.780 ;
        RECT 1707.130 1656.580 1708.830 1656.720 ;
        RECT 1707.130 1656.520 1707.450 1656.580 ;
        RECT 1708.510 1656.520 1708.830 1656.580 ;
        RECT 1706.670 1642.100 1706.990 1642.160 ;
        RECT 1706.475 1641.960 1706.990 1642.100 ;
        RECT 1706.670 1641.900 1706.990 1641.960 ;
        RECT 1706.685 1594.160 1706.975 1594.205 ;
        RECT 1707.130 1594.160 1707.450 1594.220 ;
        RECT 1706.685 1594.020 1707.450 1594.160 ;
        RECT 1706.685 1593.975 1706.975 1594.020 ;
        RECT 1707.130 1593.960 1707.450 1594.020 ;
        RECT 1706.210 1559.480 1706.530 1559.540 ;
        RECT 1707.130 1559.480 1707.450 1559.540 ;
        RECT 1706.210 1559.340 1707.450 1559.480 ;
        RECT 1706.210 1559.280 1706.530 1559.340 ;
        RECT 1707.130 1559.280 1707.450 1559.340 ;
        RECT 1705.765 1545.540 1706.055 1545.585 ;
        RECT 1706.210 1545.540 1706.530 1545.600 ;
        RECT 1705.765 1545.400 1706.530 1545.540 ;
        RECT 1705.765 1545.355 1706.055 1545.400 ;
        RECT 1706.210 1545.340 1706.530 1545.400 ;
        RECT 1705.750 1497.600 1706.070 1497.660 ;
        RECT 1705.555 1497.460 1706.070 1497.600 ;
        RECT 1705.750 1497.400 1706.070 1497.460 ;
        RECT 1705.765 1448.980 1706.055 1449.025 ;
        RECT 1706.210 1448.980 1706.530 1449.040 ;
        RECT 1705.765 1448.840 1706.530 1448.980 ;
        RECT 1705.765 1448.795 1706.055 1448.840 ;
        RECT 1706.210 1448.780 1706.530 1448.840 ;
        RECT 1705.750 1401.040 1706.070 1401.100 ;
        RECT 1705.555 1400.900 1706.070 1401.040 ;
        RECT 1705.750 1400.840 1706.070 1400.900 ;
        RECT 1705.765 1352.420 1706.055 1352.465 ;
        RECT 1706.210 1352.420 1706.530 1352.480 ;
        RECT 1705.765 1352.280 1706.530 1352.420 ;
        RECT 1705.765 1352.235 1706.055 1352.280 ;
        RECT 1706.210 1352.220 1706.530 1352.280 ;
        RECT 1705.750 1304.480 1706.070 1304.540 ;
        RECT 1705.555 1304.340 1706.070 1304.480 ;
        RECT 1705.750 1304.280 1706.070 1304.340 ;
        RECT 1706.210 1221.860 1706.530 1221.920 ;
        RECT 1705.840 1221.720 1706.530 1221.860 ;
        RECT 1705.840 1221.240 1705.980 1221.720 ;
        RECT 1706.210 1221.660 1706.530 1221.720 ;
        RECT 1705.750 1220.980 1706.070 1221.240 ;
        RECT 1706.210 1152.500 1706.530 1152.560 ;
        RECT 1707.130 1152.500 1707.450 1152.560 ;
        RECT 1706.210 1152.360 1707.450 1152.500 ;
        RECT 1706.210 1152.300 1706.530 1152.360 ;
        RECT 1707.130 1152.300 1707.450 1152.360 ;
        RECT 1706.210 1125.300 1706.530 1125.360 ;
        RECT 1705.840 1125.160 1706.530 1125.300 ;
        RECT 1705.840 1124.680 1705.980 1125.160 ;
        RECT 1706.210 1125.100 1706.530 1125.160 ;
        RECT 1705.750 1124.420 1706.070 1124.680 ;
        RECT 1705.750 1103.880 1706.070 1103.940 ;
        RECT 1705.555 1103.740 1706.070 1103.880 ;
        RECT 1705.750 1103.680 1706.070 1103.740 ;
        RECT 1705.750 1076.340 1706.070 1076.400 ;
        RECT 1705.555 1076.200 1706.070 1076.340 ;
        RECT 1705.750 1076.140 1706.070 1076.200 ;
        RECT 1705.750 1014.460 1706.070 1014.520 ;
        RECT 1706.210 1014.460 1706.530 1014.520 ;
        RECT 1705.750 1014.320 1706.530 1014.460 ;
        RECT 1705.750 1014.260 1706.070 1014.320 ;
        RECT 1706.210 1014.260 1706.530 1014.320 ;
        RECT 1706.210 966.180 1706.530 966.240 ;
        RECT 1707.130 966.180 1707.450 966.240 ;
        RECT 1706.210 966.040 1707.450 966.180 ;
        RECT 1706.210 965.980 1706.530 966.040 ;
        RECT 1707.130 965.980 1707.450 966.040 ;
        RECT 1705.750 910.760 1706.070 910.820 ;
        RECT 1706.210 910.760 1706.530 910.820 ;
        RECT 1705.750 910.620 1706.530 910.760 ;
        RECT 1705.750 910.560 1706.070 910.620 ;
        RECT 1706.210 910.560 1706.530 910.620 ;
        RECT 1705.290 824.740 1705.610 824.800 ;
        RECT 1706.210 824.740 1706.530 824.800 ;
        RECT 1705.290 824.600 1706.530 824.740 ;
        RECT 1705.290 824.540 1705.610 824.600 ;
        RECT 1706.210 824.540 1706.530 824.600 ;
        RECT 1704.370 821.000 1704.690 821.060 ;
        RECT 1705.290 821.000 1705.610 821.060 ;
        RECT 1704.370 820.860 1705.610 821.000 ;
        RECT 1704.370 820.800 1704.690 820.860 ;
        RECT 1705.290 820.800 1705.610 820.860 ;
        RECT 1706.210 693.500 1706.530 693.560 ;
        RECT 1706.685 693.500 1706.975 693.545 ;
        RECT 1706.210 693.360 1706.975 693.500 ;
        RECT 1706.210 693.300 1706.530 693.360 ;
        RECT 1706.685 693.315 1706.975 693.360 ;
        RECT 1706.670 641.480 1706.990 641.540 ;
        RECT 1706.475 641.340 1706.990 641.480 ;
        RECT 1706.670 641.280 1706.990 641.340 ;
        RECT 1706.210 593.540 1706.530 593.600 ;
        RECT 1707.130 593.540 1707.450 593.600 ;
        RECT 1706.210 593.400 1707.450 593.540 ;
        RECT 1706.210 593.340 1706.530 593.400 ;
        RECT 1707.130 593.340 1707.450 593.400 ;
        RECT 1705.765 579.600 1706.055 579.645 ;
        RECT 1706.210 579.600 1706.530 579.660 ;
        RECT 1705.765 579.460 1706.530 579.600 ;
        RECT 1705.765 579.415 1706.055 579.460 ;
        RECT 1706.210 579.400 1706.530 579.460 ;
        RECT 1705.750 531.660 1706.070 531.720 ;
        RECT 1705.555 531.520 1706.070 531.660 ;
        RECT 1705.750 531.460 1706.070 531.520 ;
        RECT 1705.750 496.780 1706.070 497.040 ;
        RECT 1705.840 496.640 1705.980 496.780 ;
        RECT 1706.210 496.640 1706.530 496.700 ;
        RECT 1705.840 496.500 1706.530 496.640 ;
        RECT 1706.210 496.440 1706.530 496.500 ;
        RECT 1705.305 434.760 1705.595 434.805 ;
        RECT 1705.750 434.760 1706.070 434.820 ;
        RECT 1705.305 434.620 1706.070 434.760 ;
        RECT 1705.305 434.575 1705.595 434.620 ;
        RECT 1705.750 434.560 1706.070 434.620 ;
        RECT 1705.290 386.480 1705.610 386.540 ;
        RECT 1705.095 386.340 1705.610 386.480 ;
        RECT 1705.290 386.280 1705.610 386.340 ;
        RECT 1705.290 385.800 1705.610 385.860 ;
        RECT 1705.095 385.660 1705.610 385.800 ;
        RECT 1705.290 385.600 1705.610 385.660 ;
        RECT 1705.305 351.460 1705.595 351.505 ;
        RECT 1705.750 351.460 1706.070 351.520 ;
        RECT 1705.305 351.320 1706.070 351.460 ;
        RECT 1705.305 351.275 1705.595 351.320 ;
        RECT 1705.750 351.260 1706.070 351.320 ;
        RECT 1706.670 282.780 1706.990 282.840 ;
        RECT 1706.475 282.640 1706.990 282.780 ;
        RECT 1706.670 282.580 1706.990 282.640 ;
        RECT 1706.670 253.200 1706.990 253.260 ;
        RECT 1706.475 253.060 1706.990 253.200 ;
        RECT 1706.670 253.000 1706.990 253.060 ;
        RECT 1705.750 158.820 1706.070 159.080 ;
        RECT 1705.840 158.400 1705.980 158.820 ;
        RECT 1705.750 158.140 1706.070 158.400 ;
        RECT 1706.210 96.800 1706.530 96.860 ;
        RECT 1706.670 96.800 1706.990 96.860 ;
        RECT 1706.210 96.660 1706.990 96.800 ;
        RECT 1706.210 96.600 1706.530 96.660 ;
        RECT 1706.670 96.600 1706.990 96.660 ;
        RECT 1442.170 32.200 1442.490 32.260 ;
        RECT 1706.210 32.200 1706.530 32.260 ;
        RECT 1442.170 32.060 1706.530 32.200 ;
        RECT 1442.170 32.000 1442.490 32.060 ;
        RECT 1706.210 32.000 1706.530 32.060 ;
        RECT 1442.170 16.560 1442.490 16.620 ;
        RECT 1382.000 16.420 1442.490 16.560 ;
        RECT 1364.430 15.880 1364.750 15.940 ;
        RECT 1382.000 15.880 1382.140 16.420 ;
        RECT 1442.170 16.360 1442.490 16.420 ;
        RECT 1364.430 15.740 1382.140 15.880 ;
        RECT 1364.430 15.680 1364.750 15.740 ;
      LAYER via ;
        RECT 1707.160 1656.520 1707.420 1656.780 ;
        RECT 1708.540 1656.520 1708.800 1656.780 ;
        RECT 1706.700 1641.900 1706.960 1642.160 ;
        RECT 1707.160 1593.960 1707.420 1594.220 ;
        RECT 1706.240 1559.280 1706.500 1559.540 ;
        RECT 1707.160 1559.280 1707.420 1559.540 ;
        RECT 1706.240 1545.340 1706.500 1545.600 ;
        RECT 1705.780 1497.400 1706.040 1497.660 ;
        RECT 1706.240 1448.780 1706.500 1449.040 ;
        RECT 1705.780 1400.840 1706.040 1401.100 ;
        RECT 1706.240 1352.220 1706.500 1352.480 ;
        RECT 1705.780 1304.280 1706.040 1304.540 ;
        RECT 1706.240 1221.660 1706.500 1221.920 ;
        RECT 1705.780 1220.980 1706.040 1221.240 ;
        RECT 1706.240 1152.300 1706.500 1152.560 ;
        RECT 1707.160 1152.300 1707.420 1152.560 ;
        RECT 1706.240 1125.100 1706.500 1125.360 ;
        RECT 1705.780 1124.420 1706.040 1124.680 ;
        RECT 1705.780 1103.680 1706.040 1103.940 ;
        RECT 1705.780 1076.140 1706.040 1076.400 ;
        RECT 1705.780 1014.260 1706.040 1014.520 ;
        RECT 1706.240 1014.260 1706.500 1014.520 ;
        RECT 1706.240 965.980 1706.500 966.240 ;
        RECT 1707.160 965.980 1707.420 966.240 ;
        RECT 1705.780 910.560 1706.040 910.820 ;
        RECT 1706.240 910.560 1706.500 910.820 ;
        RECT 1705.320 824.540 1705.580 824.800 ;
        RECT 1706.240 824.540 1706.500 824.800 ;
        RECT 1704.400 820.800 1704.660 821.060 ;
        RECT 1705.320 820.800 1705.580 821.060 ;
        RECT 1706.240 693.300 1706.500 693.560 ;
        RECT 1706.700 641.280 1706.960 641.540 ;
        RECT 1706.240 593.340 1706.500 593.600 ;
        RECT 1707.160 593.340 1707.420 593.600 ;
        RECT 1706.240 579.400 1706.500 579.660 ;
        RECT 1705.780 531.460 1706.040 531.720 ;
        RECT 1705.780 496.780 1706.040 497.040 ;
        RECT 1706.240 496.440 1706.500 496.700 ;
        RECT 1705.780 434.560 1706.040 434.820 ;
        RECT 1705.320 386.280 1705.580 386.540 ;
        RECT 1705.320 385.600 1705.580 385.860 ;
        RECT 1705.780 351.260 1706.040 351.520 ;
        RECT 1706.700 282.580 1706.960 282.840 ;
        RECT 1706.700 253.000 1706.960 253.260 ;
        RECT 1705.780 158.820 1706.040 159.080 ;
        RECT 1705.780 158.140 1706.040 158.400 ;
        RECT 1706.240 96.600 1706.500 96.860 ;
        RECT 1706.700 96.600 1706.960 96.860 ;
        RECT 1442.200 32.000 1442.460 32.260 ;
        RECT 1706.240 32.000 1706.500 32.260 ;
        RECT 1364.460 15.680 1364.720 15.940 ;
        RECT 1442.200 16.360 1442.460 16.620 ;
      LAYER met2 ;
        RECT 1710.765 1700.410 1711.045 1704.000 ;
        RECT 1708.600 1700.270 1711.045 1700.410 ;
        RECT 1708.600 1656.810 1708.740 1700.270 ;
        RECT 1710.765 1700.000 1711.045 1700.270 ;
        RECT 1707.160 1656.490 1707.420 1656.810 ;
        RECT 1708.540 1656.490 1708.800 1656.810 ;
        RECT 1707.220 1642.610 1707.360 1656.490 ;
        RECT 1706.760 1642.470 1707.360 1642.610 ;
        RECT 1706.760 1642.190 1706.900 1642.470 ;
        RECT 1706.700 1641.870 1706.960 1642.190 ;
        RECT 1707.160 1593.930 1707.420 1594.250 ;
        RECT 1707.220 1559.570 1707.360 1593.930 ;
        RECT 1706.240 1559.250 1706.500 1559.570 ;
        RECT 1707.160 1559.250 1707.420 1559.570 ;
        RECT 1706.300 1545.630 1706.440 1559.250 ;
        RECT 1706.240 1545.310 1706.500 1545.630 ;
        RECT 1705.780 1497.370 1706.040 1497.690 ;
        RECT 1705.840 1497.090 1705.980 1497.370 ;
        RECT 1706.230 1497.090 1706.510 1497.205 ;
        RECT 1705.840 1496.950 1706.510 1497.090 ;
        RECT 1706.230 1496.835 1706.510 1496.950 ;
        RECT 1706.230 1449.235 1706.510 1449.605 ;
        RECT 1706.300 1449.070 1706.440 1449.235 ;
        RECT 1706.240 1448.750 1706.500 1449.070 ;
        RECT 1705.780 1400.810 1706.040 1401.130 ;
        RECT 1705.840 1400.530 1705.980 1400.810 ;
        RECT 1706.230 1400.530 1706.510 1400.645 ;
        RECT 1705.840 1400.390 1706.510 1400.530 ;
        RECT 1706.230 1400.275 1706.510 1400.390 ;
        RECT 1706.230 1352.675 1706.510 1353.045 ;
        RECT 1706.300 1352.510 1706.440 1352.675 ;
        RECT 1706.240 1352.190 1706.500 1352.510 ;
        RECT 1705.780 1304.250 1706.040 1304.570 ;
        RECT 1705.840 1303.970 1705.980 1304.250 ;
        RECT 1706.230 1303.970 1706.510 1304.085 ;
        RECT 1705.840 1303.830 1706.510 1303.970 ;
        RECT 1706.230 1303.715 1706.510 1303.830 ;
        RECT 1706.230 1256.115 1706.510 1256.485 ;
        RECT 1706.300 1221.950 1706.440 1256.115 ;
        RECT 1706.240 1221.630 1706.500 1221.950 ;
        RECT 1705.780 1220.950 1706.040 1221.270 ;
        RECT 1705.840 1200.725 1705.980 1220.950 ;
        RECT 1705.770 1200.355 1706.050 1200.725 ;
        RECT 1707.150 1200.355 1707.430 1200.725 ;
        RECT 1707.220 1152.590 1707.360 1200.355 ;
        RECT 1706.240 1152.270 1706.500 1152.590 ;
        RECT 1707.160 1152.270 1707.420 1152.590 ;
        RECT 1706.300 1125.390 1706.440 1152.270 ;
        RECT 1706.240 1125.070 1706.500 1125.390 ;
        RECT 1705.780 1124.390 1706.040 1124.710 ;
        RECT 1705.840 1103.970 1705.980 1124.390 ;
        RECT 1705.780 1103.650 1706.040 1103.970 ;
        RECT 1705.780 1076.110 1706.040 1076.430 ;
        RECT 1705.840 1055.770 1705.980 1076.110 ;
        RECT 1705.840 1055.630 1706.440 1055.770 ;
        RECT 1706.300 1014.550 1706.440 1055.630 ;
        RECT 1705.780 1014.405 1706.040 1014.550 ;
        RECT 1705.770 1014.035 1706.050 1014.405 ;
        RECT 1706.240 1014.230 1706.500 1014.550 ;
        RECT 1707.150 1014.035 1707.430 1014.405 ;
        RECT 1707.220 966.270 1707.360 1014.035 ;
        RECT 1706.240 965.950 1706.500 966.270 ;
        RECT 1707.160 965.950 1707.420 966.270 ;
        RECT 1706.300 931.330 1706.440 965.950 ;
        RECT 1705.840 931.190 1706.440 931.330 ;
        RECT 1705.840 910.850 1705.980 931.190 ;
        RECT 1705.780 910.530 1706.040 910.850 ;
        RECT 1706.240 910.530 1706.500 910.850 ;
        RECT 1706.300 824.830 1706.440 910.530 ;
        RECT 1705.320 824.510 1705.580 824.830 ;
        RECT 1706.240 824.510 1706.500 824.830 ;
        RECT 1705.380 821.090 1705.520 824.510 ;
        RECT 1704.400 820.770 1704.660 821.090 ;
        RECT 1705.320 820.770 1705.580 821.090 ;
        RECT 1704.460 773.005 1704.600 820.770 ;
        RECT 1704.390 772.635 1704.670 773.005 ;
        RECT 1706.690 772.635 1706.970 773.005 ;
        RECT 1706.760 738.210 1706.900 772.635 ;
        RECT 1706.300 738.070 1706.900 738.210 ;
        RECT 1706.300 693.590 1706.440 738.070 ;
        RECT 1706.240 693.270 1706.500 693.590 ;
        RECT 1706.700 641.250 1706.960 641.570 ;
        RECT 1706.760 628.050 1706.900 641.250 ;
        RECT 1706.760 627.910 1707.360 628.050 ;
        RECT 1707.220 593.630 1707.360 627.910 ;
        RECT 1706.240 593.310 1706.500 593.630 ;
        RECT 1707.160 593.310 1707.420 593.630 ;
        RECT 1706.300 579.690 1706.440 593.310 ;
        RECT 1706.240 579.370 1706.500 579.690 ;
        RECT 1705.780 531.430 1706.040 531.750 ;
        RECT 1705.840 497.070 1705.980 531.430 ;
        RECT 1705.780 496.750 1706.040 497.070 ;
        RECT 1706.240 496.410 1706.500 496.730 ;
        RECT 1706.300 448.530 1706.440 496.410 ;
        RECT 1705.840 448.390 1706.440 448.530 ;
        RECT 1705.840 434.850 1705.980 448.390 ;
        RECT 1705.780 434.530 1706.040 434.850 ;
        RECT 1705.320 386.250 1705.580 386.570 ;
        RECT 1705.380 385.890 1705.520 386.250 ;
        RECT 1705.320 385.570 1705.580 385.890 ;
        RECT 1705.780 351.230 1706.040 351.550 ;
        RECT 1705.840 307.770 1705.980 351.230 ;
        RECT 1705.840 307.630 1707.360 307.770 ;
        RECT 1707.220 283.290 1707.360 307.630 ;
        RECT 1706.760 283.150 1707.360 283.290 ;
        RECT 1706.760 282.870 1706.900 283.150 ;
        RECT 1706.700 282.550 1706.960 282.870 ;
        RECT 1706.700 252.970 1706.960 253.290 ;
        RECT 1706.760 192.850 1706.900 252.970 ;
        RECT 1705.840 192.710 1706.900 192.850 ;
        RECT 1705.840 159.110 1705.980 192.710 ;
        RECT 1705.780 158.790 1706.040 159.110 ;
        RECT 1705.780 158.110 1706.040 158.430 ;
        RECT 1705.840 144.685 1705.980 158.110 ;
        RECT 1705.770 144.315 1706.050 144.685 ;
        RECT 1706.690 144.315 1706.970 144.685 ;
        RECT 1706.760 96.890 1706.900 144.315 ;
        RECT 1706.240 96.570 1706.500 96.890 ;
        RECT 1706.700 96.570 1706.960 96.890 ;
        RECT 1706.300 32.290 1706.440 96.570 ;
        RECT 1442.200 31.970 1442.460 32.290 ;
        RECT 1706.240 31.970 1706.500 32.290 ;
        RECT 1442.260 16.650 1442.400 31.970 ;
        RECT 1442.200 16.330 1442.460 16.650 ;
        RECT 1364.460 15.650 1364.720 15.970 ;
        RECT 1364.520 2.400 1364.660 15.650 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
      LAYER via2 ;
        RECT 1706.230 1496.880 1706.510 1497.160 ;
        RECT 1706.230 1449.280 1706.510 1449.560 ;
        RECT 1706.230 1400.320 1706.510 1400.600 ;
        RECT 1706.230 1352.720 1706.510 1353.000 ;
        RECT 1706.230 1303.760 1706.510 1304.040 ;
        RECT 1706.230 1256.160 1706.510 1256.440 ;
        RECT 1705.770 1200.400 1706.050 1200.680 ;
        RECT 1707.150 1200.400 1707.430 1200.680 ;
        RECT 1705.770 1014.080 1706.050 1014.360 ;
        RECT 1707.150 1014.080 1707.430 1014.360 ;
        RECT 1704.390 772.680 1704.670 772.960 ;
        RECT 1706.690 772.680 1706.970 772.960 ;
        RECT 1705.770 144.360 1706.050 144.640 ;
        RECT 1706.690 144.360 1706.970 144.640 ;
      LAYER met3 ;
        RECT 1706.205 1497.170 1706.535 1497.185 ;
        RECT 1706.870 1497.170 1707.250 1497.180 ;
        RECT 1706.205 1496.870 1707.250 1497.170 ;
        RECT 1706.205 1496.855 1706.535 1496.870 ;
        RECT 1706.870 1496.860 1707.250 1496.870 ;
        RECT 1706.205 1449.570 1706.535 1449.585 ;
        RECT 1706.870 1449.570 1707.250 1449.580 ;
        RECT 1706.205 1449.270 1707.250 1449.570 ;
        RECT 1706.205 1449.255 1706.535 1449.270 ;
        RECT 1706.870 1449.260 1707.250 1449.270 ;
        RECT 1706.205 1400.610 1706.535 1400.625 ;
        RECT 1706.870 1400.610 1707.250 1400.620 ;
        RECT 1706.205 1400.310 1707.250 1400.610 ;
        RECT 1706.205 1400.295 1706.535 1400.310 ;
        RECT 1706.870 1400.300 1707.250 1400.310 ;
        RECT 1706.205 1353.010 1706.535 1353.025 ;
        RECT 1706.870 1353.010 1707.250 1353.020 ;
        RECT 1706.205 1352.710 1707.250 1353.010 ;
        RECT 1706.205 1352.695 1706.535 1352.710 ;
        RECT 1706.870 1352.700 1707.250 1352.710 ;
        RECT 1706.205 1304.050 1706.535 1304.065 ;
        RECT 1706.870 1304.050 1707.250 1304.060 ;
        RECT 1706.205 1303.750 1707.250 1304.050 ;
        RECT 1706.205 1303.735 1706.535 1303.750 ;
        RECT 1706.870 1303.740 1707.250 1303.750 ;
        RECT 1706.205 1256.450 1706.535 1256.465 ;
        RECT 1706.870 1256.450 1707.250 1256.460 ;
        RECT 1706.205 1256.150 1707.250 1256.450 ;
        RECT 1706.205 1256.135 1706.535 1256.150 ;
        RECT 1706.870 1256.140 1707.250 1256.150 ;
        RECT 1705.745 1200.690 1706.075 1200.705 ;
        RECT 1707.125 1200.690 1707.455 1200.705 ;
        RECT 1705.745 1200.390 1707.455 1200.690 ;
        RECT 1705.745 1200.375 1706.075 1200.390 ;
        RECT 1707.125 1200.375 1707.455 1200.390 ;
        RECT 1705.745 1014.370 1706.075 1014.385 ;
        RECT 1707.125 1014.370 1707.455 1014.385 ;
        RECT 1705.745 1014.070 1707.455 1014.370 ;
        RECT 1705.745 1014.055 1706.075 1014.070 ;
        RECT 1707.125 1014.055 1707.455 1014.070 ;
        RECT 1704.365 772.970 1704.695 772.985 ;
        RECT 1706.665 772.970 1706.995 772.985 ;
        RECT 1704.365 772.670 1706.995 772.970 ;
        RECT 1704.365 772.655 1704.695 772.670 ;
        RECT 1706.665 772.655 1706.995 772.670 ;
        RECT 1705.745 144.650 1706.075 144.665 ;
        RECT 1706.665 144.650 1706.995 144.665 ;
        RECT 1705.745 144.350 1706.995 144.650 ;
        RECT 1705.745 144.335 1706.075 144.350 ;
        RECT 1706.665 144.335 1706.995 144.350 ;
      LAYER via3 ;
        RECT 1706.900 1496.860 1707.220 1497.180 ;
        RECT 1706.900 1449.260 1707.220 1449.580 ;
        RECT 1706.900 1400.300 1707.220 1400.620 ;
        RECT 1706.900 1352.700 1707.220 1353.020 ;
        RECT 1706.900 1303.740 1707.220 1304.060 ;
        RECT 1706.900 1256.140 1707.220 1256.460 ;
      LAYER met4 ;
        RECT 1706.895 1496.855 1707.225 1497.185 ;
        RECT 1706.910 1449.585 1707.210 1496.855 ;
        RECT 1706.895 1449.255 1707.225 1449.585 ;
        RECT 1706.895 1400.295 1707.225 1400.625 ;
        RECT 1706.910 1353.025 1707.210 1400.295 ;
        RECT 1706.895 1352.695 1707.225 1353.025 ;
        RECT 1706.895 1303.735 1707.225 1304.065 ;
        RECT 1706.910 1256.465 1707.210 1303.735 ;
        RECT 1706.895 1256.135 1707.225 1256.465 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1442.630 31.860 1442.950 31.920 ;
        RECT 1718.170 31.860 1718.490 31.920 ;
        RECT 1442.630 31.720 1718.490 31.860 ;
        RECT 1442.630 31.660 1442.950 31.720 ;
        RECT 1718.170 31.660 1718.490 31.720 ;
        RECT 1382.370 16.220 1382.690 16.280 ;
        RECT 1442.630 16.220 1442.950 16.280 ;
        RECT 1382.370 16.080 1442.950 16.220 ;
        RECT 1382.370 16.020 1382.690 16.080 ;
        RECT 1442.630 16.020 1442.950 16.080 ;
      LAYER via ;
        RECT 1442.660 31.660 1442.920 31.920 ;
        RECT 1718.200 31.660 1718.460 31.920 ;
        RECT 1382.400 16.020 1382.660 16.280 ;
        RECT 1442.660 16.020 1442.920 16.280 ;
      LAYER met2 ;
        RECT 1718.125 1700.000 1718.405 1704.000 ;
        RECT 1718.260 31.950 1718.400 1700.000 ;
        RECT 1442.660 31.630 1442.920 31.950 ;
        RECT 1718.200 31.630 1718.460 31.950 ;
        RECT 1442.720 16.310 1442.860 31.630 ;
        RECT 1382.400 15.990 1382.660 16.310 ;
        RECT 1442.660 15.990 1442.920 16.310 ;
        RECT 1382.460 2.400 1382.600 15.990 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1400.310 31.180 1400.630 31.240 ;
        RECT 1725.990 31.180 1726.310 31.240 ;
        RECT 1400.310 31.040 1726.310 31.180 ;
        RECT 1400.310 30.980 1400.630 31.040 ;
        RECT 1725.990 30.980 1726.310 31.040 ;
      LAYER via ;
        RECT 1400.340 30.980 1400.600 31.240 ;
        RECT 1726.020 30.980 1726.280 31.240 ;
      LAYER met2 ;
        RECT 1725.485 1700.410 1725.765 1704.000 ;
        RECT 1725.485 1700.270 1726.220 1700.410 ;
        RECT 1725.485 1700.000 1725.765 1700.270 ;
        RECT 1726.080 31.270 1726.220 1700.270 ;
        RECT 1400.340 30.950 1400.600 31.270 ;
        RECT 1726.020 30.950 1726.280 31.270 ;
        RECT 1400.400 2.400 1400.540 30.950 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1418.250 26.420 1418.570 26.480 ;
        RECT 1732.890 26.420 1733.210 26.480 ;
        RECT 1418.250 26.280 1733.210 26.420 ;
        RECT 1418.250 26.220 1418.570 26.280 ;
        RECT 1732.890 26.220 1733.210 26.280 ;
      LAYER via ;
        RECT 1418.280 26.220 1418.540 26.480 ;
        RECT 1732.920 26.220 1733.180 26.480 ;
      LAYER met2 ;
        RECT 1732.845 1700.000 1733.125 1704.000 ;
        RECT 1732.980 26.510 1733.120 1700.000 ;
        RECT 1418.280 26.190 1418.540 26.510 ;
        RECT 1732.920 26.190 1733.180 26.510 ;
        RECT 1418.340 2.400 1418.480 26.190 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1435.730 26.760 1436.050 26.820 ;
        RECT 1739.790 26.760 1740.110 26.820 ;
        RECT 1435.730 26.620 1740.110 26.760 ;
        RECT 1435.730 26.560 1436.050 26.620 ;
        RECT 1739.790 26.560 1740.110 26.620 ;
      LAYER via ;
        RECT 1435.760 26.560 1436.020 26.820 ;
        RECT 1739.820 26.560 1740.080 26.820 ;
      LAYER met2 ;
        RECT 1740.205 1700.410 1740.485 1704.000 ;
        RECT 1739.880 1700.270 1740.485 1700.410 ;
        RECT 1739.880 26.850 1740.020 1700.270 ;
        RECT 1740.205 1700.000 1740.485 1700.270 ;
        RECT 1435.760 26.530 1436.020 26.850 ;
        RECT 1739.820 26.530 1740.080 26.850 ;
        RECT 1435.820 2.400 1435.960 26.530 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1453.670 27.100 1453.990 27.160 ;
        RECT 1746.690 27.100 1747.010 27.160 ;
        RECT 1453.670 26.960 1747.010 27.100 ;
        RECT 1453.670 26.900 1453.990 26.960 ;
        RECT 1746.690 26.900 1747.010 26.960 ;
      LAYER via ;
        RECT 1453.700 26.900 1453.960 27.160 ;
        RECT 1746.720 26.900 1746.980 27.160 ;
      LAYER met2 ;
        RECT 1747.565 1700.410 1747.845 1704.000 ;
        RECT 1746.780 1700.270 1747.845 1700.410 ;
        RECT 1746.780 27.190 1746.920 1700.270 ;
        RECT 1747.565 1700.000 1747.845 1700.270 ;
        RECT 1453.700 26.870 1453.960 27.190 ;
        RECT 1746.720 26.870 1746.980 27.190 ;
        RECT 1453.760 2.400 1453.900 26.870 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1471.610 31.520 1471.930 31.580 ;
        RECT 1753.130 31.520 1753.450 31.580 ;
        RECT 1471.610 31.380 1753.450 31.520 ;
        RECT 1471.610 31.320 1471.930 31.380 ;
        RECT 1753.130 31.320 1753.450 31.380 ;
      LAYER via ;
        RECT 1471.640 31.320 1471.900 31.580 ;
        RECT 1753.160 31.320 1753.420 31.580 ;
      LAYER met2 ;
        RECT 1754.925 1700.410 1755.205 1704.000 ;
        RECT 1753.220 1700.270 1755.205 1700.410 ;
        RECT 1753.220 31.610 1753.360 1700.270 ;
        RECT 1754.925 1700.000 1755.205 1700.270 ;
        RECT 1471.640 31.290 1471.900 31.610 ;
        RECT 1753.160 31.290 1753.420 31.610 ;
        RECT 1471.700 2.400 1471.840 31.290 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1489.090 27.440 1489.410 27.500 ;
        RECT 1760.490 27.440 1760.810 27.500 ;
        RECT 1489.090 27.300 1760.810 27.440 ;
        RECT 1489.090 27.240 1489.410 27.300 ;
        RECT 1760.490 27.240 1760.810 27.300 ;
      LAYER via ;
        RECT 1489.120 27.240 1489.380 27.500 ;
        RECT 1760.520 27.240 1760.780 27.500 ;
      LAYER met2 ;
        RECT 1762.285 1700.410 1762.565 1704.000 ;
        RECT 1760.580 1700.270 1762.565 1700.410 ;
        RECT 1760.580 27.530 1760.720 1700.270 ;
        RECT 1762.285 1700.000 1762.565 1700.270 ;
        RECT 1489.120 27.210 1489.380 27.530 ;
        RECT 1760.520 27.210 1760.780 27.530 ;
        RECT 1489.180 20.130 1489.320 27.210 ;
        RECT 1489.180 19.990 1489.780 20.130 ;
        RECT 1489.640 2.400 1489.780 19.990 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1752.745 21.845 1752.915 22.695 ;
      LAYER mcon ;
        RECT 1752.745 22.525 1752.915 22.695 ;
      LAYER met1 ;
        RECT 1752.685 22.680 1752.975 22.725 ;
        RECT 1767.390 22.680 1767.710 22.740 ;
        RECT 1752.685 22.540 1767.710 22.680 ;
        RECT 1752.685 22.495 1752.975 22.540 ;
        RECT 1767.390 22.480 1767.710 22.540 ;
        RECT 1507.030 22.000 1507.350 22.060 ;
        RECT 1752.685 22.000 1752.975 22.045 ;
        RECT 1507.030 21.860 1752.975 22.000 ;
        RECT 1507.030 21.800 1507.350 21.860 ;
        RECT 1752.685 21.815 1752.975 21.860 ;
      LAYER via ;
        RECT 1767.420 22.480 1767.680 22.740 ;
        RECT 1507.060 21.800 1507.320 22.060 ;
      LAYER met2 ;
        RECT 1769.645 1700.410 1769.925 1704.000 ;
        RECT 1767.480 1700.270 1769.925 1700.410 ;
        RECT 1767.480 22.770 1767.620 1700.270 ;
        RECT 1769.645 1700.000 1769.925 1700.270 ;
        RECT 1767.420 22.450 1767.680 22.770 ;
        RECT 1507.060 21.770 1507.320 22.090 ;
        RECT 1507.120 2.400 1507.260 21.770 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 710.310 59.740 710.630 59.800 ;
        RECT 1436.650 59.740 1436.970 59.800 ;
        RECT 710.310 59.600 1436.970 59.740 ;
        RECT 710.310 59.540 710.630 59.600 ;
        RECT 1436.650 59.540 1436.970 59.600 ;
        RECT 704.330 20.980 704.650 21.040 ;
        RECT 710.310 20.980 710.630 21.040 ;
        RECT 704.330 20.840 710.630 20.980 ;
        RECT 704.330 20.780 704.650 20.840 ;
        RECT 710.310 20.780 710.630 20.840 ;
      LAYER via ;
        RECT 710.340 59.540 710.600 59.800 ;
        RECT 1436.680 59.540 1436.940 59.800 ;
        RECT 704.360 20.780 704.620 21.040 ;
        RECT 710.340 20.780 710.600 21.040 ;
      LAYER met2 ;
        RECT 1438.905 1700.410 1439.185 1704.000 ;
        RECT 1436.740 1700.270 1439.185 1700.410 ;
        RECT 1436.740 59.830 1436.880 1700.270 ;
        RECT 1438.905 1700.000 1439.185 1700.270 ;
        RECT 710.340 59.510 710.600 59.830 ;
        RECT 1436.680 59.510 1436.940 59.830 ;
        RECT 710.400 21.070 710.540 59.510 ;
        RECT 704.360 20.750 704.620 21.070 ;
        RECT 710.340 20.750 710.600 21.070 ;
        RECT 704.420 2.400 704.560 20.750 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1524.970 21.660 1525.290 21.720 ;
        RECT 1774.750 21.660 1775.070 21.720 ;
        RECT 1524.970 21.520 1775.070 21.660 ;
        RECT 1524.970 21.460 1525.290 21.520 ;
        RECT 1774.750 21.460 1775.070 21.520 ;
      LAYER via ;
        RECT 1525.000 21.460 1525.260 21.720 ;
        RECT 1774.780 21.460 1775.040 21.720 ;
      LAYER met2 ;
        RECT 1777.005 1700.410 1777.285 1704.000 ;
        RECT 1774.840 1700.270 1777.285 1700.410 ;
        RECT 1774.840 21.750 1774.980 1700.270 ;
        RECT 1777.005 1700.000 1777.285 1700.270 ;
        RECT 1525.000 21.430 1525.260 21.750 ;
        RECT 1774.780 21.430 1775.040 21.750 ;
        RECT 1525.060 2.400 1525.200 21.430 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1780.730 1678.140 1781.050 1678.200 ;
        RECT 1783.030 1678.140 1783.350 1678.200 ;
        RECT 1780.730 1678.000 1783.350 1678.140 ;
        RECT 1780.730 1677.940 1781.050 1678.000 ;
        RECT 1783.030 1677.940 1783.350 1678.000 ;
        RECT 1542.910 21.320 1543.230 21.380 ;
        RECT 1780.730 21.320 1781.050 21.380 ;
        RECT 1542.910 21.180 1781.050 21.320 ;
        RECT 1542.910 21.120 1543.230 21.180 ;
        RECT 1780.730 21.120 1781.050 21.180 ;
      LAYER via ;
        RECT 1780.760 1677.940 1781.020 1678.200 ;
        RECT 1783.060 1677.940 1783.320 1678.200 ;
        RECT 1542.940 21.120 1543.200 21.380 ;
        RECT 1780.760 21.120 1781.020 21.380 ;
      LAYER met2 ;
        RECT 1784.365 1700.410 1784.645 1704.000 ;
        RECT 1783.120 1700.270 1784.645 1700.410 ;
        RECT 1783.120 1678.230 1783.260 1700.270 ;
        RECT 1784.365 1700.000 1784.645 1700.270 ;
        RECT 1780.760 1677.910 1781.020 1678.230 ;
        RECT 1783.060 1677.910 1783.320 1678.230 ;
        RECT 1780.820 21.410 1780.960 1677.910 ;
        RECT 1542.940 21.090 1543.200 21.410 ;
        RECT 1780.760 21.090 1781.020 21.410 ;
        RECT 1543.000 2.400 1543.140 21.090 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1788.165 689.605 1788.335 724.455 ;
        RECT 1787.705 620.925 1787.875 669.375 ;
        RECT 1788.165 496.485 1788.335 548.675 ;
        RECT 1788.165 386.325 1788.335 434.775 ;
        RECT 1788.165 241.485 1788.335 289.595 ;
      LAYER mcon ;
        RECT 1788.165 724.285 1788.335 724.455 ;
        RECT 1787.705 669.205 1787.875 669.375 ;
        RECT 1788.165 548.505 1788.335 548.675 ;
        RECT 1788.165 434.605 1788.335 434.775 ;
        RECT 1788.165 289.425 1788.335 289.595 ;
      LAYER met1 ;
        RECT 1788.090 1594.160 1788.410 1594.220 ;
        RECT 1788.550 1594.160 1788.870 1594.220 ;
        RECT 1788.090 1594.020 1788.870 1594.160 ;
        RECT 1788.090 1593.960 1788.410 1594.020 ;
        RECT 1788.550 1593.960 1788.870 1594.020 ;
        RECT 1787.630 1511.200 1787.950 1511.260 ;
        RECT 1788.550 1511.200 1788.870 1511.260 ;
        RECT 1787.630 1511.060 1788.870 1511.200 ;
        RECT 1787.630 1511.000 1787.950 1511.060 ;
        RECT 1788.550 1511.000 1788.870 1511.060 ;
        RECT 1787.630 1414.640 1787.950 1414.700 ;
        RECT 1788.550 1414.640 1788.870 1414.700 ;
        RECT 1787.630 1414.500 1788.870 1414.640 ;
        RECT 1787.630 1414.440 1787.950 1414.500 ;
        RECT 1788.550 1414.440 1788.870 1414.500 ;
        RECT 1787.630 1318.080 1787.950 1318.140 ;
        RECT 1788.550 1318.080 1788.870 1318.140 ;
        RECT 1787.630 1317.940 1788.870 1318.080 ;
        RECT 1787.630 1317.880 1787.950 1317.940 ;
        RECT 1788.550 1317.880 1788.870 1317.940 ;
        RECT 1787.630 1221.520 1787.950 1221.580 ;
        RECT 1788.550 1221.520 1788.870 1221.580 ;
        RECT 1787.630 1221.380 1788.870 1221.520 ;
        RECT 1787.630 1221.320 1787.950 1221.380 ;
        RECT 1788.550 1221.320 1788.870 1221.380 ;
        RECT 1787.630 1124.960 1787.950 1125.020 ;
        RECT 1788.550 1124.960 1788.870 1125.020 ;
        RECT 1787.630 1124.820 1788.870 1124.960 ;
        RECT 1787.630 1124.760 1787.950 1124.820 ;
        RECT 1788.550 1124.760 1788.870 1124.820 ;
        RECT 1787.630 1028.400 1787.950 1028.460 ;
        RECT 1788.550 1028.400 1788.870 1028.460 ;
        RECT 1787.630 1028.260 1788.870 1028.400 ;
        RECT 1787.630 1028.200 1787.950 1028.260 ;
        RECT 1788.550 1028.200 1788.870 1028.260 ;
        RECT 1787.630 931.840 1787.950 931.900 ;
        RECT 1788.550 931.840 1788.870 931.900 ;
        RECT 1787.630 931.700 1788.870 931.840 ;
        RECT 1787.630 931.640 1787.950 931.700 ;
        RECT 1788.550 931.640 1788.870 931.700 ;
        RECT 1787.170 869.620 1787.490 869.680 ;
        RECT 1788.550 869.620 1788.870 869.680 ;
        RECT 1787.170 869.480 1788.870 869.620 ;
        RECT 1787.170 869.420 1787.490 869.480 ;
        RECT 1788.550 869.420 1788.870 869.480 ;
        RECT 1787.630 835.280 1787.950 835.340 ;
        RECT 1788.550 835.280 1788.870 835.340 ;
        RECT 1787.630 835.140 1788.870 835.280 ;
        RECT 1787.630 835.080 1787.950 835.140 ;
        RECT 1788.550 835.080 1788.870 835.140 ;
        RECT 1788.090 786.800 1788.410 787.060 ;
        RECT 1788.180 786.320 1788.320 786.800 ;
        RECT 1788.550 786.320 1788.870 786.380 ;
        RECT 1788.180 786.180 1788.870 786.320 ;
        RECT 1788.550 786.120 1788.870 786.180 ;
        RECT 1787.630 738.380 1787.950 738.440 ;
        RECT 1788.550 738.380 1788.870 738.440 ;
        RECT 1787.630 738.240 1788.870 738.380 ;
        RECT 1787.630 738.180 1787.950 738.240 ;
        RECT 1788.550 738.180 1788.870 738.240 ;
        RECT 1788.090 724.440 1788.410 724.500 ;
        RECT 1787.895 724.300 1788.410 724.440 ;
        RECT 1788.090 724.240 1788.410 724.300 ;
        RECT 1788.090 689.760 1788.410 689.820 ;
        RECT 1787.895 689.620 1788.410 689.760 ;
        RECT 1788.090 689.560 1788.410 689.620 ;
        RECT 1787.630 676.160 1787.950 676.220 ;
        RECT 1788.550 676.160 1788.870 676.220 ;
        RECT 1787.630 676.020 1788.870 676.160 ;
        RECT 1787.630 675.960 1787.950 676.020 ;
        RECT 1788.550 675.960 1788.870 676.020 ;
        RECT 1787.630 669.360 1787.950 669.420 ;
        RECT 1787.435 669.220 1787.950 669.360 ;
        RECT 1787.630 669.160 1787.950 669.220 ;
        RECT 1787.645 621.080 1787.935 621.125 ;
        RECT 1788.090 621.080 1788.410 621.140 ;
        RECT 1787.645 620.940 1788.410 621.080 ;
        RECT 1787.645 620.895 1787.935 620.940 ;
        RECT 1788.090 620.880 1788.410 620.940 ;
        RECT 1788.105 548.660 1788.395 548.705 ;
        RECT 1788.550 548.660 1788.870 548.720 ;
        RECT 1788.105 548.520 1788.870 548.660 ;
        RECT 1788.105 548.475 1788.395 548.520 ;
        RECT 1788.550 548.460 1788.870 548.520 ;
        RECT 1788.090 496.640 1788.410 496.700 ;
        RECT 1787.895 496.500 1788.410 496.640 ;
        RECT 1788.090 496.440 1788.410 496.500 ;
        RECT 1787.630 448.700 1787.950 448.760 ;
        RECT 1788.550 448.700 1788.870 448.760 ;
        RECT 1787.630 448.560 1788.870 448.700 ;
        RECT 1787.630 448.500 1787.950 448.560 ;
        RECT 1788.550 448.500 1788.870 448.560 ;
        RECT 1788.090 434.760 1788.410 434.820 ;
        RECT 1787.895 434.620 1788.410 434.760 ;
        RECT 1788.090 434.560 1788.410 434.620 ;
        RECT 1788.105 386.480 1788.395 386.525 ;
        RECT 1788.550 386.480 1788.870 386.540 ;
        RECT 1788.105 386.340 1788.870 386.480 ;
        RECT 1788.105 386.295 1788.395 386.340 ;
        RECT 1788.550 386.280 1788.870 386.340 ;
        RECT 1788.550 338.540 1788.870 338.600 ;
        RECT 1788.180 338.400 1788.870 338.540 ;
        RECT 1788.180 338.260 1788.320 338.400 ;
        RECT 1788.550 338.340 1788.870 338.400 ;
        RECT 1788.090 338.000 1788.410 338.260 ;
        RECT 1788.105 289.580 1788.395 289.625 ;
        RECT 1788.550 289.580 1788.870 289.640 ;
        RECT 1788.105 289.440 1788.870 289.580 ;
        RECT 1788.105 289.395 1788.395 289.440 ;
        RECT 1788.550 289.380 1788.870 289.440 ;
        RECT 1788.090 241.640 1788.410 241.700 ;
        RECT 1787.895 241.500 1788.410 241.640 ;
        RECT 1788.090 241.440 1788.410 241.500 ;
        RECT 1788.550 145.420 1788.870 145.480 ;
        RECT 1788.180 145.280 1788.870 145.420 ;
        RECT 1788.180 145.140 1788.320 145.280 ;
        RECT 1788.550 145.220 1788.870 145.280 ;
        RECT 1788.090 144.880 1788.410 145.140 ;
        RECT 1560.850 20.980 1561.170 21.040 ;
        RECT 1787.630 20.980 1787.950 21.040 ;
        RECT 1560.850 20.840 1787.950 20.980 ;
        RECT 1560.850 20.780 1561.170 20.840 ;
        RECT 1787.630 20.780 1787.950 20.840 ;
      LAYER via ;
        RECT 1788.120 1593.960 1788.380 1594.220 ;
        RECT 1788.580 1593.960 1788.840 1594.220 ;
        RECT 1787.660 1511.000 1787.920 1511.260 ;
        RECT 1788.580 1511.000 1788.840 1511.260 ;
        RECT 1787.660 1414.440 1787.920 1414.700 ;
        RECT 1788.580 1414.440 1788.840 1414.700 ;
        RECT 1787.660 1317.880 1787.920 1318.140 ;
        RECT 1788.580 1317.880 1788.840 1318.140 ;
        RECT 1787.660 1221.320 1787.920 1221.580 ;
        RECT 1788.580 1221.320 1788.840 1221.580 ;
        RECT 1787.660 1124.760 1787.920 1125.020 ;
        RECT 1788.580 1124.760 1788.840 1125.020 ;
        RECT 1787.660 1028.200 1787.920 1028.460 ;
        RECT 1788.580 1028.200 1788.840 1028.460 ;
        RECT 1787.660 931.640 1787.920 931.900 ;
        RECT 1788.580 931.640 1788.840 931.900 ;
        RECT 1787.200 869.420 1787.460 869.680 ;
        RECT 1788.580 869.420 1788.840 869.680 ;
        RECT 1787.660 835.080 1787.920 835.340 ;
        RECT 1788.580 835.080 1788.840 835.340 ;
        RECT 1788.120 786.800 1788.380 787.060 ;
        RECT 1788.580 786.120 1788.840 786.380 ;
        RECT 1787.660 738.180 1787.920 738.440 ;
        RECT 1788.580 738.180 1788.840 738.440 ;
        RECT 1788.120 724.240 1788.380 724.500 ;
        RECT 1788.120 689.560 1788.380 689.820 ;
        RECT 1787.660 675.960 1787.920 676.220 ;
        RECT 1788.580 675.960 1788.840 676.220 ;
        RECT 1787.660 669.160 1787.920 669.420 ;
        RECT 1788.120 620.880 1788.380 621.140 ;
        RECT 1788.580 548.460 1788.840 548.720 ;
        RECT 1788.120 496.440 1788.380 496.700 ;
        RECT 1787.660 448.500 1787.920 448.760 ;
        RECT 1788.580 448.500 1788.840 448.760 ;
        RECT 1788.120 434.560 1788.380 434.820 ;
        RECT 1788.580 386.280 1788.840 386.540 ;
        RECT 1788.580 338.340 1788.840 338.600 ;
        RECT 1788.120 338.000 1788.380 338.260 ;
        RECT 1788.580 289.380 1788.840 289.640 ;
        RECT 1788.120 241.440 1788.380 241.700 ;
        RECT 1788.580 145.220 1788.840 145.480 ;
        RECT 1788.120 144.880 1788.380 145.140 ;
        RECT 1560.880 20.780 1561.140 21.040 ;
        RECT 1787.660 20.780 1787.920 21.040 ;
      LAYER met2 ;
        RECT 1791.725 1701.090 1792.005 1704.000 ;
        RECT 1789.560 1700.950 1792.005 1701.090 ;
        RECT 1789.560 1677.970 1789.700 1700.950 ;
        RECT 1791.725 1700.000 1792.005 1700.950 ;
        RECT 1788.640 1677.830 1789.700 1677.970 ;
        RECT 1788.640 1594.250 1788.780 1677.830 ;
        RECT 1788.120 1593.930 1788.380 1594.250 ;
        RECT 1788.580 1593.930 1788.840 1594.250 ;
        RECT 1788.180 1559.650 1788.320 1593.930 ;
        RECT 1788.180 1559.510 1788.780 1559.650 ;
        RECT 1788.640 1511.290 1788.780 1559.510 ;
        RECT 1787.660 1510.970 1787.920 1511.290 ;
        RECT 1788.580 1510.970 1788.840 1511.290 ;
        RECT 1787.720 1510.690 1787.860 1510.970 ;
        RECT 1787.720 1510.550 1788.320 1510.690 ;
        RECT 1788.180 1463.090 1788.320 1510.550 ;
        RECT 1788.180 1462.950 1788.780 1463.090 ;
        RECT 1788.640 1414.730 1788.780 1462.950 ;
        RECT 1787.660 1414.410 1787.920 1414.730 ;
        RECT 1788.580 1414.410 1788.840 1414.730 ;
        RECT 1787.720 1414.130 1787.860 1414.410 ;
        RECT 1787.720 1413.990 1788.320 1414.130 ;
        RECT 1788.180 1366.530 1788.320 1413.990 ;
        RECT 1788.180 1366.390 1788.780 1366.530 ;
        RECT 1788.640 1318.170 1788.780 1366.390 ;
        RECT 1787.660 1317.850 1787.920 1318.170 ;
        RECT 1788.580 1317.850 1788.840 1318.170 ;
        RECT 1787.720 1317.570 1787.860 1317.850 ;
        RECT 1787.720 1317.430 1788.320 1317.570 ;
        RECT 1788.180 1269.970 1788.320 1317.430 ;
        RECT 1788.180 1269.830 1788.780 1269.970 ;
        RECT 1788.640 1221.610 1788.780 1269.830 ;
        RECT 1787.660 1221.290 1787.920 1221.610 ;
        RECT 1788.580 1221.290 1788.840 1221.610 ;
        RECT 1787.720 1221.010 1787.860 1221.290 ;
        RECT 1787.720 1220.870 1788.320 1221.010 ;
        RECT 1788.180 1173.410 1788.320 1220.870 ;
        RECT 1788.180 1173.270 1788.780 1173.410 ;
        RECT 1788.640 1125.050 1788.780 1173.270 ;
        RECT 1787.660 1124.730 1787.920 1125.050 ;
        RECT 1788.580 1124.730 1788.840 1125.050 ;
        RECT 1787.720 1124.450 1787.860 1124.730 ;
        RECT 1787.720 1124.310 1788.320 1124.450 ;
        RECT 1788.180 1076.850 1788.320 1124.310 ;
        RECT 1788.180 1076.710 1788.780 1076.850 ;
        RECT 1788.640 1028.490 1788.780 1076.710 ;
        RECT 1787.660 1028.170 1787.920 1028.490 ;
        RECT 1788.580 1028.170 1788.840 1028.490 ;
        RECT 1787.720 1027.890 1787.860 1028.170 ;
        RECT 1787.720 1027.750 1788.320 1027.890 ;
        RECT 1788.180 980.290 1788.320 1027.750 ;
        RECT 1788.180 980.150 1788.780 980.290 ;
        RECT 1788.640 931.930 1788.780 980.150 ;
        RECT 1787.660 931.610 1787.920 931.930 ;
        RECT 1788.580 931.610 1788.840 931.930 ;
        RECT 1787.720 931.330 1787.860 931.610 ;
        RECT 1787.720 931.190 1788.320 931.330 ;
        RECT 1788.180 917.845 1788.320 931.190 ;
        RECT 1787.190 917.475 1787.470 917.845 ;
        RECT 1788.110 917.475 1788.390 917.845 ;
        RECT 1787.260 869.710 1787.400 917.475 ;
        RECT 1787.200 869.390 1787.460 869.710 ;
        RECT 1788.580 869.390 1788.840 869.710 ;
        RECT 1788.640 835.370 1788.780 869.390 ;
        RECT 1787.660 835.050 1787.920 835.370 ;
        RECT 1788.580 835.050 1788.840 835.370 ;
        RECT 1787.720 834.770 1787.860 835.050 ;
        RECT 1787.720 834.630 1788.320 834.770 ;
        RECT 1788.180 787.090 1788.320 834.630 ;
        RECT 1788.120 786.770 1788.380 787.090 ;
        RECT 1788.580 786.090 1788.840 786.410 ;
        RECT 1788.640 738.470 1788.780 786.090 ;
        RECT 1787.660 738.210 1787.920 738.470 ;
        RECT 1787.660 738.150 1788.320 738.210 ;
        RECT 1788.580 738.150 1788.840 738.470 ;
        RECT 1787.720 738.070 1788.320 738.150 ;
        RECT 1788.180 724.530 1788.320 738.070 ;
        RECT 1788.120 724.210 1788.380 724.530 ;
        RECT 1788.120 689.530 1788.380 689.850 ;
        RECT 1788.180 676.330 1788.320 689.530 ;
        RECT 1788.180 676.250 1788.780 676.330 ;
        RECT 1787.660 675.930 1787.920 676.250 ;
        RECT 1788.180 676.190 1788.840 676.250 ;
        RECT 1788.580 675.930 1788.840 676.190 ;
        RECT 1787.720 669.450 1787.860 675.930 ;
        RECT 1788.640 675.775 1788.780 675.930 ;
        RECT 1787.660 669.130 1787.920 669.450 ;
        RECT 1788.120 620.850 1788.380 621.170 ;
        RECT 1788.180 620.685 1788.320 620.850 ;
        RECT 1788.110 620.315 1788.390 620.685 ;
        RECT 1789.030 620.315 1789.310 620.685 ;
        RECT 1789.100 593.370 1789.240 620.315 ;
        RECT 1788.640 593.230 1789.240 593.370 ;
        RECT 1788.640 548.750 1788.780 593.230 ;
        RECT 1788.580 548.430 1788.840 548.750 ;
        RECT 1788.120 496.410 1788.380 496.730 ;
        RECT 1788.180 483.210 1788.320 496.410 ;
        RECT 1788.180 483.070 1788.780 483.210 ;
        RECT 1788.640 448.790 1788.780 483.070 ;
        RECT 1787.660 448.530 1787.920 448.790 ;
        RECT 1787.660 448.470 1788.320 448.530 ;
        RECT 1788.580 448.470 1788.840 448.790 ;
        RECT 1787.720 448.390 1788.320 448.470 ;
        RECT 1788.180 434.850 1788.320 448.390 ;
        RECT 1788.120 434.530 1788.380 434.850 ;
        RECT 1788.580 386.250 1788.840 386.570 ;
        RECT 1788.640 338.630 1788.780 386.250 ;
        RECT 1788.580 338.310 1788.840 338.630 ;
        RECT 1788.120 337.970 1788.380 338.290 ;
        RECT 1788.180 303.690 1788.320 337.970 ;
        RECT 1788.180 303.550 1788.780 303.690 ;
        RECT 1788.640 289.670 1788.780 303.550 ;
        RECT 1788.580 289.350 1788.840 289.670 ;
        RECT 1788.120 241.410 1788.380 241.730 ;
        RECT 1788.180 207.130 1788.320 241.410 ;
        RECT 1788.180 206.990 1788.780 207.130 ;
        RECT 1788.640 145.510 1788.780 206.990 ;
        RECT 1788.580 145.190 1788.840 145.510 ;
        RECT 1788.120 144.850 1788.380 145.170 ;
        RECT 1788.180 110.570 1788.320 144.850 ;
        RECT 1788.180 110.430 1788.780 110.570 ;
        RECT 1788.640 62.290 1788.780 110.430 ;
        RECT 1787.720 62.150 1788.780 62.290 ;
        RECT 1787.720 21.070 1787.860 62.150 ;
        RECT 1560.880 20.750 1561.140 21.070 ;
        RECT 1787.660 20.750 1787.920 21.070 ;
        RECT 1560.940 2.400 1561.080 20.750 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
      LAYER via2 ;
        RECT 1787.190 917.520 1787.470 917.800 ;
        RECT 1788.110 917.520 1788.390 917.800 ;
        RECT 1788.110 620.360 1788.390 620.640 ;
        RECT 1789.030 620.360 1789.310 620.640 ;
      LAYER met3 ;
        RECT 1787.165 917.810 1787.495 917.825 ;
        RECT 1788.085 917.810 1788.415 917.825 ;
        RECT 1787.165 917.510 1788.415 917.810 ;
        RECT 1787.165 917.495 1787.495 917.510 ;
        RECT 1788.085 917.495 1788.415 917.510 ;
        RECT 1788.085 620.650 1788.415 620.665 ;
        RECT 1789.005 620.650 1789.335 620.665 ;
        RECT 1788.085 620.350 1789.335 620.650 ;
        RECT 1788.085 620.335 1788.415 620.350 ;
        RECT 1789.005 620.335 1789.335 620.350 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1794.990 1678.140 1795.310 1678.200 ;
        RECT 1796.830 1678.140 1797.150 1678.200 ;
        RECT 1794.990 1678.000 1797.150 1678.140 ;
        RECT 1794.990 1677.940 1795.310 1678.000 ;
        RECT 1796.830 1677.940 1797.150 1678.000 ;
        RECT 1616.510 23.700 1616.830 23.760 ;
        RECT 1794.990 23.700 1795.310 23.760 ;
        RECT 1616.510 23.560 1795.310 23.700 ;
        RECT 1616.510 23.500 1616.830 23.560 ;
        RECT 1794.990 23.500 1795.310 23.560 ;
        RECT 1578.790 15.200 1579.110 15.260 ;
        RECT 1616.510 15.200 1616.830 15.260 ;
        RECT 1578.790 15.060 1616.830 15.200 ;
        RECT 1578.790 15.000 1579.110 15.060 ;
        RECT 1616.510 15.000 1616.830 15.060 ;
      LAYER via ;
        RECT 1795.020 1677.940 1795.280 1678.200 ;
        RECT 1796.860 1677.940 1797.120 1678.200 ;
        RECT 1616.540 23.500 1616.800 23.760 ;
        RECT 1795.020 23.500 1795.280 23.760 ;
        RECT 1578.820 15.000 1579.080 15.260 ;
        RECT 1616.540 15.000 1616.800 15.260 ;
      LAYER met2 ;
        RECT 1798.625 1700.410 1798.905 1704.000 ;
        RECT 1796.920 1700.270 1798.905 1700.410 ;
        RECT 1796.920 1678.230 1797.060 1700.270 ;
        RECT 1798.625 1700.000 1798.905 1700.270 ;
        RECT 1795.020 1677.910 1795.280 1678.230 ;
        RECT 1796.860 1677.910 1797.120 1678.230 ;
        RECT 1795.080 23.790 1795.220 1677.910 ;
        RECT 1616.540 23.470 1616.800 23.790 ;
        RECT 1795.020 23.470 1795.280 23.790 ;
        RECT 1616.600 15.290 1616.740 23.470 ;
        RECT 1578.820 14.970 1579.080 15.290 ;
        RECT 1616.540 14.970 1616.800 15.290 ;
        RECT 1578.880 2.400 1579.020 14.970 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1631.690 24.380 1632.010 24.440 ;
        RECT 1801.890 24.380 1802.210 24.440 ;
        RECT 1631.690 24.240 1802.210 24.380 ;
        RECT 1631.690 24.180 1632.010 24.240 ;
        RECT 1801.890 24.180 1802.210 24.240 ;
        RECT 1596.270 14.520 1596.590 14.580 ;
        RECT 1631.690 14.520 1632.010 14.580 ;
        RECT 1596.270 14.380 1632.010 14.520 ;
        RECT 1596.270 14.320 1596.590 14.380 ;
        RECT 1631.690 14.320 1632.010 14.380 ;
      LAYER via ;
        RECT 1631.720 24.180 1631.980 24.440 ;
        RECT 1801.920 24.180 1802.180 24.440 ;
        RECT 1596.300 14.320 1596.560 14.580 ;
        RECT 1631.720 14.320 1631.980 14.580 ;
      LAYER met2 ;
        RECT 1805.985 1700.410 1806.265 1704.000 ;
        RECT 1804.740 1700.270 1806.265 1700.410 ;
        RECT 1804.740 1687.490 1804.880 1700.270 ;
        RECT 1805.985 1700.000 1806.265 1700.270 ;
        RECT 1801.980 1687.350 1804.880 1687.490 ;
        RECT 1801.980 24.470 1802.120 1687.350 ;
        RECT 1631.720 24.150 1631.980 24.470 ;
        RECT 1801.920 24.150 1802.180 24.470 ;
        RECT 1631.780 14.610 1631.920 24.150 ;
        RECT 1596.300 14.290 1596.560 14.610 ;
        RECT 1631.720 14.290 1631.980 14.610 ;
        RECT 1596.360 2.400 1596.500 14.290 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1808.330 1688.680 1808.650 1688.740 ;
        RECT 1811.550 1688.680 1811.870 1688.740 ;
        RECT 1808.330 1688.540 1811.870 1688.680 ;
        RECT 1808.330 1688.480 1808.650 1688.540 ;
        RECT 1811.550 1688.480 1811.870 1688.540 ;
        RECT 1635.370 24.720 1635.690 24.780 ;
        RECT 1808.330 24.720 1808.650 24.780 ;
        RECT 1635.370 24.580 1808.650 24.720 ;
        RECT 1635.370 24.520 1635.690 24.580 ;
        RECT 1808.330 24.520 1808.650 24.580 ;
        RECT 1614.210 17.920 1614.530 17.980 ;
        RECT 1635.370 17.920 1635.690 17.980 ;
        RECT 1614.210 17.780 1635.690 17.920 ;
        RECT 1614.210 17.720 1614.530 17.780 ;
        RECT 1635.370 17.720 1635.690 17.780 ;
      LAYER via ;
        RECT 1808.360 1688.480 1808.620 1688.740 ;
        RECT 1811.580 1688.480 1811.840 1688.740 ;
        RECT 1635.400 24.520 1635.660 24.780 ;
        RECT 1808.360 24.520 1808.620 24.780 ;
        RECT 1614.240 17.720 1614.500 17.980 ;
        RECT 1635.400 17.720 1635.660 17.980 ;
      LAYER met2 ;
        RECT 1813.345 1700.410 1813.625 1704.000 ;
        RECT 1811.640 1700.270 1813.625 1700.410 ;
        RECT 1811.640 1688.770 1811.780 1700.270 ;
        RECT 1813.345 1700.000 1813.625 1700.270 ;
        RECT 1808.360 1688.450 1808.620 1688.770 ;
        RECT 1811.580 1688.450 1811.840 1688.770 ;
        RECT 1808.420 24.810 1808.560 1688.450 ;
        RECT 1635.400 24.490 1635.660 24.810 ;
        RECT 1808.360 24.490 1808.620 24.810 ;
        RECT 1635.460 18.010 1635.600 24.490 ;
        RECT 1614.240 17.690 1614.500 18.010 ;
        RECT 1635.400 17.690 1635.660 18.010 ;
        RECT 1614.300 2.400 1614.440 17.690 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1815.230 1688.680 1815.550 1688.740 ;
        RECT 1818.910 1688.680 1819.230 1688.740 ;
        RECT 1815.230 1688.540 1819.230 1688.680 ;
        RECT 1815.230 1688.480 1815.550 1688.540 ;
        RECT 1818.910 1688.480 1819.230 1688.540 ;
        RECT 1642.270 24.040 1642.590 24.100 ;
        RECT 1815.230 24.040 1815.550 24.100 ;
        RECT 1642.270 23.900 1815.550 24.040 ;
        RECT 1642.270 23.840 1642.590 23.900 ;
        RECT 1815.230 23.840 1815.550 23.900 ;
        RECT 1632.150 18.600 1632.470 18.660 ;
        RECT 1642.270 18.600 1642.590 18.660 ;
        RECT 1632.150 18.460 1642.590 18.600 ;
        RECT 1632.150 18.400 1632.470 18.460 ;
        RECT 1642.270 18.400 1642.590 18.460 ;
      LAYER via ;
        RECT 1815.260 1688.480 1815.520 1688.740 ;
        RECT 1818.940 1688.480 1819.200 1688.740 ;
        RECT 1642.300 23.840 1642.560 24.100 ;
        RECT 1815.260 23.840 1815.520 24.100 ;
        RECT 1632.180 18.400 1632.440 18.660 ;
        RECT 1642.300 18.400 1642.560 18.660 ;
      LAYER met2 ;
        RECT 1820.705 1700.410 1820.985 1704.000 ;
        RECT 1819.000 1700.270 1820.985 1700.410 ;
        RECT 1819.000 1688.770 1819.140 1700.270 ;
        RECT 1820.705 1700.000 1820.985 1700.270 ;
        RECT 1815.260 1688.450 1815.520 1688.770 ;
        RECT 1818.940 1688.450 1819.200 1688.770 ;
        RECT 1815.320 24.130 1815.460 1688.450 ;
        RECT 1642.300 23.810 1642.560 24.130 ;
        RECT 1815.260 23.810 1815.520 24.130 ;
        RECT 1642.360 18.690 1642.500 23.810 ;
        RECT 1632.180 18.370 1632.440 18.690 ;
        RECT 1642.300 18.370 1642.560 18.690 ;
        RECT 1632.240 2.400 1632.380 18.370 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1703.065 15.725 1703.695 15.895 ;
        RECT 1703.525 14.365 1703.695 15.725 ;
      LAYER met1 ;
        RECT 1828.110 1689.360 1828.430 1689.420 ;
        RECT 1776.680 1689.220 1828.430 1689.360 ;
        RECT 1742.090 1688.340 1742.410 1688.400 ;
        RECT 1776.680 1688.340 1776.820 1689.220 ;
        RECT 1828.110 1689.160 1828.430 1689.220 ;
        RECT 1742.090 1688.200 1776.820 1688.340 ;
        RECT 1742.090 1688.140 1742.410 1688.200 ;
        RECT 1728.750 16.560 1729.070 16.620 ;
        RECT 1742.090 16.560 1742.410 16.620 ;
        RECT 1728.750 16.420 1742.410 16.560 ;
        RECT 1728.750 16.360 1729.070 16.420 ;
        RECT 1742.090 16.360 1742.410 16.420 ;
        RECT 1679.530 15.880 1679.850 15.940 ;
        RECT 1703.005 15.880 1703.295 15.925 ;
        RECT 1679.530 15.740 1703.295 15.880 ;
        RECT 1679.530 15.680 1679.850 15.740 ;
        RECT 1703.005 15.695 1703.295 15.740 ;
        RECT 1703.465 14.520 1703.755 14.565 ;
        RECT 1704.370 14.520 1704.690 14.580 ;
        RECT 1703.465 14.380 1704.690 14.520 ;
        RECT 1703.465 14.335 1703.755 14.380 ;
        RECT 1704.370 14.320 1704.690 14.380 ;
        RECT 1650.090 14.180 1650.410 14.240 ;
        RECT 1677.690 14.180 1678.010 14.240 ;
        RECT 1650.090 14.040 1678.010 14.180 ;
        RECT 1650.090 13.980 1650.410 14.040 ;
        RECT 1677.690 13.980 1678.010 14.040 ;
      LAYER via ;
        RECT 1742.120 1688.140 1742.380 1688.400 ;
        RECT 1828.140 1689.160 1828.400 1689.420 ;
        RECT 1728.780 16.360 1729.040 16.620 ;
        RECT 1742.120 16.360 1742.380 16.620 ;
        RECT 1679.560 15.680 1679.820 15.940 ;
        RECT 1704.400 14.320 1704.660 14.580 ;
        RECT 1650.120 13.980 1650.380 14.240 ;
        RECT 1677.720 13.980 1677.980 14.240 ;
      LAYER met2 ;
        RECT 1828.065 1700.000 1828.345 1704.000 ;
        RECT 1828.200 1689.450 1828.340 1700.000 ;
        RECT 1828.140 1689.130 1828.400 1689.450 ;
        RECT 1742.120 1688.110 1742.380 1688.430 ;
        RECT 1742.180 16.650 1742.320 1688.110 ;
        RECT 1728.780 16.330 1729.040 16.650 ;
        RECT 1742.120 16.330 1742.380 16.650 ;
        RECT 1677.780 15.970 1679.760 16.050 ;
        RECT 1677.780 15.910 1679.820 15.970 ;
        RECT 1677.780 14.270 1677.920 15.910 ;
        RECT 1679.560 15.650 1679.820 15.910 ;
        RECT 1728.840 15.485 1728.980 16.330 ;
        RECT 1704.390 15.115 1704.670 15.485 ;
        RECT 1728.770 15.115 1729.050 15.485 ;
        RECT 1704.460 14.610 1704.600 15.115 ;
        RECT 1704.400 14.290 1704.660 14.610 ;
        RECT 1650.120 13.950 1650.380 14.270 ;
        RECT 1677.720 13.950 1677.980 14.270 ;
        RECT 1650.180 2.400 1650.320 13.950 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
      LAYER via2 ;
        RECT 1704.390 15.160 1704.670 15.440 ;
        RECT 1728.770 15.160 1729.050 15.440 ;
      LAYER met3 ;
        RECT 1704.365 15.450 1704.695 15.465 ;
        RECT 1728.745 15.450 1729.075 15.465 ;
        RECT 1704.365 15.150 1729.075 15.450 ;
        RECT 1704.365 15.135 1704.695 15.150 ;
        RECT 1728.745 15.135 1729.075 15.150 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1668.030 25.060 1668.350 25.120 ;
        RECT 1835.930 25.060 1836.250 25.120 ;
        RECT 1668.030 24.920 1836.250 25.060 ;
        RECT 1668.030 24.860 1668.350 24.920 ;
        RECT 1835.930 24.860 1836.250 24.920 ;
      LAYER via ;
        RECT 1668.060 24.860 1668.320 25.120 ;
        RECT 1835.960 24.860 1836.220 25.120 ;
      LAYER met2 ;
        RECT 1835.425 1700.410 1835.705 1704.000 ;
        RECT 1835.425 1700.270 1836.160 1700.410 ;
        RECT 1835.425 1700.000 1835.705 1700.270 ;
        RECT 1836.020 25.150 1836.160 1700.270 ;
        RECT 1668.060 24.830 1668.320 25.150 ;
        RECT 1835.960 24.830 1836.220 25.150 ;
        RECT 1668.120 2.400 1668.260 24.830 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1685.510 25.400 1685.830 25.460 ;
        RECT 1842.830 25.400 1843.150 25.460 ;
        RECT 1685.510 25.260 1843.150 25.400 ;
        RECT 1685.510 25.200 1685.830 25.260 ;
        RECT 1842.830 25.200 1843.150 25.260 ;
      LAYER via ;
        RECT 1685.540 25.200 1685.800 25.460 ;
        RECT 1842.860 25.200 1843.120 25.460 ;
      LAYER met2 ;
        RECT 1842.785 1700.000 1843.065 1704.000 ;
        RECT 1842.920 25.490 1843.060 1700.000 ;
        RECT 1685.540 25.170 1685.800 25.490 ;
        RECT 1842.860 25.170 1843.120 25.490 ;
        RECT 1685.600 2.400 1685.740 25.170 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1443.625 1531.785 1443.795 1538.755 ;
        RECT 1444.545 1373.345 1444.715 1421.455 ;
        RECT 1444.085 1207.425 1444.255 1295.655 ;
        RECT 1443.625 241.485 1443.795 285.175 ;
      LAYER mcon ;
        RECT 1443.625 1538.585 1443.795 1538.755 ;
        RECT 1444.545 1421.285 1444.715 1421.455 ;
        RECT 1444.085 1295.485 1444.255 1295.655 ;
        RECT 1443.625 285.005 1443.795 285.175 ;
      LAYER met1 ;
        RECT 1443.550 1628.500 1443.870 1628.560 ;
        RECT 1444.010 1628.500 1444.330 1628.560 ;
        RECT 1443.550 1628.360 1444.330 1628.500 ;
        RECT 1443.550 1628.300 1443.870 1628.360 ;
        RECT 1444.010 1628.300 1444.330 1628.360 ;
        RECT 1443.565 1538.740 1443.855 1538.785 ;
        RECT 1444.010 1538.740 1444.330 1538.800 ;
        RECT 1443.565 1538.600 1444.330 1538.740 ;
        RECT 1443.565 1538.555 1443.855 1538.600 ;
        RECT 1444.010 1538.540 1444.330 1538.600 ;
        RECT 1443.550 1531.940 1443.870 1532.000 ;
        RECT 1443.355 1531.800 1443.870 1531.940 ;
        RECT 1443.550 1531.740 1443.870 1531.800 ;
        RECT 1444.470 1490.600 1444.790 1490.860 ;
        RECT 1444.560 1490.180 1444.700 1490.600 ;
        RECT 1444.470 1489.920 1444.790 1490.180 ;
        RECT 1444.485 1421.440 1444.775 1421.485 ;
        RECT 1444.930 1421.440 1445.250 1421.500 ;
        RECT 1444.485 1421.300 1445.250 1421.440 ;
        RECT 1444.485 1421.255 1444.775 1421.300 ;
        RECT 1444.930 1421.240 1445.250 1421.300 ;
        RECT 1444.470 1373.500 1444.790 1373.560 ;
        RECT 1444.275 1373.360 1444.790 1373.500 ;
        RECT 1444.470 1373.300 1444.790 1373.360 ;
        RECT 1444.025 1295.640 1444.315 1295.685 ;
        RECT 1444.470 1295.640 1444.790 1295.700 ;
        RECT 1444.025 1295.500 1444.790 1295.640 ;
        RECT 1444.025 1295.455 1444.315 1295.500 ;
        RECT 1444.470 1295.440 1444.790 1295.500 ;
        RECT 1444.010 1207.580 1444.330 1207.640 ;
        RECT 1443.815 1207.440 1444.330 1207.580 ;
        RECT 1444.010 1207.380 1444.330 1207.440 ;
        RECT 1443.550 1152.500 1443.870 1152.560 ;
        RECT 1444.010 1152.500 1444.330 1152.560 ;
        RECT 1443.550 1152.360 1444.330 1152.500 ;
        RECT 1443.550 1152.300 1443.870 1152.360 ;
        RECT 1444.010 1152.300 1444.330 1152.360 ;
        RECT 1443.550 1124.760 1443.870 1125.020 ;
        RECT 1443.640 1124.280 1443.780 1124.760 ;
        RECT 1444.010 1124.280 1444.330 1124.340 ;
        RECT 1443.640 1124.140 1444.330 1124.280 ;
        RECT 1444.010 1124.080 1444.330 1124.140 ;
        RECT 1443.550 1028.200 1443.870 1028.460 ;
        RECT 1443.640 1028.060 1443.780 1028.200 ;
        RECT 1444.010 1028.060 1444.330 1028.120 ;
        RECT 1443.640 1027.920 1444.330 1028.060 ;
        RECT 1444.010 1027.860 1444.330 1027.920 ;
        RECT 1443.550 966.180 1443.870 966.240 ;
        RECT 1444.470 966.180 1444.790 966.240 ;
        RECT 1443.550 966.040 1444.790 966.180 ;
        RECT 1443.550 965.980 1443.870 966.040 ;
        RECT 1444.470 965.980 1444.790 966.040 ;
        RECT 1443.550 869.620 1443.870 869.680 ;
        RECT 1444.470 869.620 1444.790 869.680 ;
        RECT 1443.550 869.480 1444.790 869.620 ;
        RECT 1443.550 869.420 1443.870 869.480 ;
        RECT 1444.470 869.420 1444.790 869.480 ;
        RECT 1443.550 613.940 1443.870 614.000 ;
        RECT 1444.010 613.940 1444.330 614.000 ;
        RECT 1443.550 613.800 1444.330 613.940 ;
        RECT 1443.550 613.740 1443.870 613.800 ;
        RECT 1444.010 613.740 1444.330 613.800 ;
        RECT 1443.550 285.160 1443.870 285.220 ;
        RECT 1443.355 285.020 1443.870 285.160 ;
        RECT 1443.550 284.960 1443.870 285.020 ;
        RECT 1443.550 241.640 1443.870 241.700 ;
        RECT 1443.355 241.500 1443.870 241.640 ;
        RECT 1443.550 241.440 1443.870 241.500 ;
        RECT 1444.010 186.220 1444.330 186.280 ;
        RECT 1444.470 186.220 1444.790 186.280 ;
        RECT 1444.010 186.080 1444.790 186.220 ;
        RECT 1444.010 186.020 1444.330 186.080 ;
        RECT 1444.470 186.020 1444.790 186.080 ;
        RECT 724.110 60.080 724.430 60.140 ;
        RECT 1444.470 60.080 1444.790 60.140 ;
        RECT 724.110 59.940 1444.790 60.080 ;
        RECT 724.110 59.880 724.430 59.940 ;
        RECT 1444.470 59.880 1444.790 59.940 ;
      LAYER via ;
        RECT 1443.580 1628.300 1443.840 1628.560 ;
        RECT 1444.040 1628.300 1444.300 1628.560 ;
        RECT 1444.040 1538.540 1444.300 1538.800 ;
        RECT 1443.580 1531.740 1443.840 1532.000 ;
        RECT 1444.500 1490.600 1444.760 1490.860 ;
        RECT 1444.500 1489.920 1444.760 1490.180 ;
        RECT 1444.960 1421.240 1445.220 1421.500 ;
        RECT 1444.500 1373.300 1444.760 1373.560 ;
        RECT 1444.500 1295.440 1444.760 1295.700 ;
        RECT 1444.040 1207.380 1444.300 1207.640 ;
        RECT 1443.580 1152.300 1443.840 1152.560 ;
        RECT 1444.040 1152.300 1444.300 1152.560 ;
        RECT 1443.580 1124.760 1443.840 1125.020 ;
        RECT 1444.040 1124.080 1444.300 1124.340 ;
        RECT 1443.580 1028.200 1443.840 1028.460 ;
        RECT 1444.040 1027.860 1444.300 1028.120 ;
        RECT 1443.580 965.980 1443.840 966.240 ;
        RECT 1444.500 965.980 1444.760 966.240 ;
        RECT 1443.580 869.420 1443.840 869.680 ;
        RECT 1444.500 869.420 1444.760 869.680 ;
        RECT 1443.580 613.740 1443.840 614.000 ;
        RECT 1444.040 613.740 1444.300 614.000 ;
        RECT 1443.580 284.960 1443.840 285.220 ;
        RECT 1443.580 241.440 1443.840 241.700 ;
        RECT 1444.040 186.020 1444.300 186.280 ;
        RECT 1444.500 186.020 1444.760 186.280 ;
        RECT 724.140 59.880 724.400 60.140 ;
        RECT 1444.500 59.880 1444.760 60.140 ;
      LAYER met2 ;
        RECT 1446.265 1700.410 1446.545 1704.000 ;
        RECT 1445.020 1700.270 1446.545 1700.410 ;
        RECT 1445.020 1676.725 1445.160 1700.270 ;
        RECT 1446.265 1700.000 1446.545 1700.270 ;
        RECT 1443.570 1676.355 1443.850 1676.725 ;
        RECT 1444.950 1676.355 1445.230 1676.725 ;
        RECT 1443.640 1628.590 1443.780 1676.355 ;
        RECT 1443.580 1628.270 1443.840 1628.590 ;
        RECT 1444.040 1628.270 1444.300 1628.590 ;
        RECT 1444.100 1538.830 1444.240 1628.270 ;
        RECT 1444.040 1538.510 1444.300 1538.830 ;
        RECT 1443.580 1531.885 1443.840 1532.030 ;
        RECT 1443.570 1531.515 1443.850 1531.885 ;
        RECT 1444.490 1531.515 1444.770 1531.885 ;
        RECT 1444.560 1490.890 1444.700 1531.515 ;
        RECT 1444.500 1490.570 1444.760 1490.890 ;
        RECT 1444.500 1489.890 1444.760 1490.210 ;
        RECT 1444.560 1448.980 1444.700 1489.890 ;
        RECT 1444.560 1448.840 1445.160 1448.980 ;
        RECT 1445.020 1448.130 1445.160 1448.840 ;
        RECT 1444.560 1447.990 1445.160 1448.130 ;
        RECT 1444.560 1442.010 1444.700 1447.990 ;
        RECT 1444.560 1441.870 1445.160 1442.010 ;
        RECT 1445.020 1421.530 1445.160 1441.870 ;
        RECT 1444.960 1421.210 1445.220 1421.530 ;
        RECT 1444.500 1373.270 1444.760 1373.590 ;
        RECT 1444.560 1295.730 1444.700 1373.270 ;
        RECT 1444.500 1295.410 1444.760 1295.730 ;
        RECT 1444.040 1207.350 1444.300 1207.670 ;
        RECT 1444.100 1152.590 1444.240 1207.350 ;
        RECT 1443.580 1152.270 1443.840 1152.590 ;
        RECT 1444.040 1152.270 1444.300 1152.590 ;
        RECT 1443.640 1125.050 1443.780 1152.270 ;
        RECT 1443.580 1124.730 1443.840 1125.050 ;
        RECT 1444.040 1124.050 1444.300 1124.370 ;
        RECT 1444.100 1104.165 1444.240 1124.050 ;
        RECT 1444.030 1103.795 1444.310 1104.165 ;
        RECT 1443.570 1103.115 1443.850 1103.485 ;
        RECT 1443.640 1028.490 1443.780 1103.115 ;
        RECT 1443.580 1028.170 1443.840 1028.490 ;
        RECT 1444.040 1027.830 1444.300 1028.150 ;
        RECT 1444.100 990.490 1444.240 1027.830 ;
        RECT 1444.100 990.350 1444.700 990.490 ;
        RECT 1444.560 966.270 1444.700 990.350 ;
        RECT 1443.580 966.125 1443.840 966.270 ;
        RECT 1444.500 966.125 1444.760 966.270 ;
        RECT 1443.570 965.755 1443.850 966.125 ;
        RECT 1444.490 965.755 1444.770 966.125 ;
        RECT 1444.560 931.330 1444.700 965.755 ;
        RECT 1444.100 931.190 1444.700 931.330 ;
        RECT 1444.100 893.930 1444.240 931.190 ;
        RECT 1444.100 893.790 1444.700 893.930 ;
        RECT 1444.560 869.710 1444.700 893.790 ;
        RECT 1443.580 869.390 1443.840 869.710 ;
        RECT 1444.500 869.390 1444.760 869.710 ;
        RECT 1443.640 845.650 1443.780 869.390 ;
        RECT 1443.640 845.510 1444.240 845.650 ;
        RECT 1444.100 783.770 1444.240 845.510 ;
        RECT 1443.640 783.630 1444.240 783.770 ;
        RECT 1443.640 645.050 1443.780 783.630 ;
        RECT 1443.640 644.910 1444.240 645.050 ;
        RECT 1444.100 614.030 1444.240 644.910 ;
        RECT 1443.580 613.710 1443.840 614.030 ;
        RECT 1444.040 613.710 1444.300 614.030 ;
        RECT 1443.640 339.730 1443.780 613.710 ;
        RECT 1443.180 339.590 1443.780 339.730 ;
        RECT 1443.180 338.370 1443.320 339.590 ;
        RECT 1443.180 338.230 1443.780 338.370 ;
        RECT 1443.640 285.250 1443.780 338.230 ;
        RECT 1443.580 284.930 1443.840 285.250 ;
        RECT 1443.580 241.410 1443.840 241.730 ;
        RECT 1443.640 210.530 1443.780 241.410 ;
        RECT 1443.640 210.390 1444.700 210.530 ;
        RECT 1444.560 192.850 1444.700 210.390 ;
        RECT 1444.100 192.710 1444.700 192.850 ;
        RECT 1444.100 186.310 1444.240 192.710 ;
        RECT 1444.040 185.990 1444.300 186.310 ;
        RECT 1444.500 185.990 1444.760 186.310 ;
        RECT 1444.560 60.170 1444.700 185.990 ;
        RECT 724.140 59.850 724.400 60.170 ;
        RECT 1444.500 59.850 1444.760 60.170 ;
        RECT 724.200 17.410 724.340 59.850 ;
        RECT 722.360 17.270 724.340 17.410 ;
        RECT 722.360 2.400 722.500 17.270 ;
        RECT 722.150 -4.800 722.710 2.400 ;
      LAYER via2 ;
        RECT 1443.570 1676.400 1443.850 1676.680 ;
        RECT 1444.950 1676.400 1445.230 1676.680 ;
        RECT 1443.570 1531.560 1443.850 1531.840 ;
        RECT 1444.490 1531.560 1444.770 1531.840 ;
        RECT 1444.030 1103.840 1444.310 1104.120 ;
        RECT 1443.570 1103.160 1443.850 1103.440 ;
        RECT 1443.570 965.800 1443.850 966.080 ;
        RECT 1444.490 965.800 1444.770 966.080 ;
      LAYER met3 ;
        RECT 1443.545 1676.690 1443.875 1676.705 ;
        RECT 1444.925 1676.690 1445.255 1676.705 ;
        RECT 1443.545 1676.390 1445.255 1676.690 ;
        RECT 1443.545 1676.375 1443.875 1676.390 ;
        RECT 1444.925 1676.375 1445.255 1676.390 ;
        RECT 1443.545 1531.850 1443.875 1531.865 ;
        RECT 1444.465 1531.850 1444.795 1531.865 ;
        RECT 1443.545 1531.550 1444.795 1531.850 ;
        RECT 1443.545 1531.535 1443.875 1531.550 ;
        RECT 1444.465 1531.535 1444.795 1531.550 ;
        RECT 1444.005 1104.130 1444.335 1104.145 ;
        RECT 1443.790 1103.815 1444.335 1104.130 ;
        RECT 1443.790 1103.465 1444.090 1103.815 ;
        RECT 1443.545 1103.150 1444.090 1103.465 ;
        RECT 1443.545 1103.135 1443.875 1103.150 ;
        RECT 1443.545 966.090 1443.875 966.105 ;
        RECT 1444.465 966.090 1444.795 966.105 ;
        RECT 1443.545 965.790 1444.795 966.090 ;
        RECT 1443.545 965.775 1443.875 965.790 ;
        RECT 1444.465 965.775 1444.795 965.790 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1729.745 15.725 1729.915 16.915 ;
        RECT 1764.705 16.745 1764.875 19.975 ;
      LAYER mcon ;
        RECT 1764.705 19.805 1764.875 19.975 ;
        RECT 1729.745 16.745 1729.915 16.915 ;
      LAYER met1 ;
        RECT 1776.590 1689.700 1776.910 1689.760 ;
        RECT 1850.190 1689.700 1850.510 1689.760 ;
        RECT 1776.590 1689.560 1850.510 1689.700 ;
        RECT 1776.590 1689.500 1776.910 1689.560 ;
        RECT 1850.190 1689.500 1850.510 1689.560 ;
        RECT 1764.645 19.960 1764.935 20.005 ;
        RECT 1776.590 19.960 1776.910 20.020 ;
        RECT 1764.645 19.820 1776.910 19.960 ;
        RECT 1764.645 19.775 1764.935 19.820 ;
        RECT 1776.590 19.760 1776.910 19.820 ;
        RECT 1729.685 16.900 1729.975 16.945 ;
        RECT 1764.645 16.900 1764.935 16.945 ;
        RECT 1729.685 16.760 1764.935 16.900 ;
        RECT 1729.685 16.715 1729.975 16.760 ;
        RECT 1764.645 16.715 1764.935 16.760 ;
        RECT 1703.450 15.880 1703.770 15.940 ;
        RECT 1729.685 15.880 1729.975 15.925 ;
        RECT 1703.450 15.740 1729.975 15.880 ;
        RECT 1703.450 15.680 1703.770 15.740 ;
        RECT 1729.685 15.695 1729.975 15.740 ;
      LAYER via ;
        RECT 1776.620 1689.500 1776.880 1689.760 ;
        RECT 1850.220 1689.500 1850.480 1689.760 ;
        RECT 1776.620 19.760 1776.880 20.020 ;
        RECT 1703.480 15.680 1703.740 15.940 ;
      LAYER met2 ;
        RECT 1850.145 1700.000 1850.425 1704.000 ;
        RECT 1850.280 1689.790 1850.420 1700.000 ;
        RECT 1776.620 1689.470 1776.880 1689.790 ;
        RECT 1850.220 1689.470 1850.480 1689.790 ;
        RECT 1776.680 20.050 1776.820 1689.470 ;
        RECT 1776.620 19.730 1776.880 20.050 ;
        RECT 1703.480 15.650 1703.740 15.970 ;
        RECT 1703.540 2.400 1703.680 15.650 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1777.585 16.915 1777.755 18.275 ;
        RECT 1774.365 16.745 1777.755 16.915 ;
        RECT 1774.365 14.705 1774.535 16.745 ;
      LAYER mcon ;
        RECT 1777.585 18.105 1777.755 18.275 ;
      LAYER met1 ;
        RECT 1790.390 1690.380 1790.710 1690.440 ;
        RECT 1857.550 1690.380 1857.870 1690.440 ;
        RECT 1790.390 1690.240 1857.870 1690.380 ;
        RECT 1790.390 1690.180 1790.710 1690.240 ;
        RECT 1857.550 1690.180 1857.870 1690.240 ;
        RECT 1777.525 18.260 1777.815 18.305 ;
        RECT 1790.390 18.260 1790.710 18.320 ;
        RECT 1777.525 18.120 1790.710 18.260 ;
        RECT 1777.525 18.075 1777.815 18.120 ;
        RECT 1790.390 18.060 1790.710 18.120 ;
        RECT 1774.305 14.860 1774.595 14.905 ;
        RECT 1753.220 14.720 1774.595 14.860 ;
        RECT 1721.390 14.520 1721.710 14.580 ;
        RECT 1753.220 14.520 1753.360 14.720 ;
        RECT 1774.305 14.675 1774.595 14.720 ;
        RECT 1721.390 14.380 1753.360 14.520 ;
        RECT 1721.390 14.320 1721.710 14.380 ;
      LAYER via ;
        RECT 1790.420 1690.180 1790.680 1690.440 ;
        RECT 1857.580 1690.180 1857.840 1690.440 ;
        RECT 1790.420 18.060 1790.680 18.320 ;
        RECT 1721.420 14.320 1721.680 14.580 ;
      LAYER met2 ;
        RECT 1857.505 1700.000 1857.785 1704.000 ;
        RECT 1857.640 1690.470 1857.780 1700.000 ;
        RECT 1790.420 1690.150 1790.680 1690.470 ;
        RECT 1857.580 1690.150 1857.840 1690.470 ;
        RECT 1790.480 18.350 1790.620 1690.150 ;
        RECT 1790.420 18.030 1790.680 18.350 ;
        RECT 1721.420 14.290 1721.680 14.610 ;
        RECT 1721.480 2.400 1721.620 14.290 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1745.310 1687.320 1745.630 1687.380 ;
        RECT 1864.910 1687.320 1865.230 1687.380 ;
        RECT 1745.310 1687.180 1865.230 1687.320 ;
        RECT 1745.310 1687.120 1745.630 1687.180 ;
        RECT 1864.910 1687.120 1865.230 1687.180 ;
        RECT 1739.330 20.640 1739.650 20.700 ;
        RECT 1745.310 20.640 1745.630 20.700 ;
        RECT 1739.330 20.500 1745.630 20.640 ;
        RECT 1739.330 20.440 1739.650 20.500 ;
        RECT 1745.310 20.440 1745.630 20.500 ;
      LAYER via ;
        RECT 1745.340 1687.120 1745.600 1687.380 ;
        RECT 1864.940 1687.120 1865.200 1687.380 ;
        RECT 1739.360 20.440 1739.620 20.700 ;
        RECT 1745.340 20.440 1745.600 20.700 ;
      LAYER met2 ;
        RECT 1864.865 1700.000 1865.145 1704.000 ;
        RECT 1865.000 1687.410 1865.140 1700.000 ;
        RECT 1745.340 1687.090 1745.600 1687.410 ;
        RECT 1864.940 1687.090 1865.200 1687.410 ;
        RECT 1745.400 20.730 1745.540 1687.090 ;
        RECT 1739.360 20.410 1739.620 20.730 ;
        RECT 1745.340 20.410 1745.600 20.730 ;
        RECT 1739.420 2.400 1739.560 20.410 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1759.110 1685.620 1759.430 1685.680 ;
        RECT 1872.270 1685.620 1872.590 1685.680 ;
        RECT 1759.110 1685.480 1872.590 1685.620 ;
        RECT 1759.110 1685.420 1759.430 1685.480 ;
        RECT 1872.270 1685.420 1872.590 1685.480 ;
        RECT 1756.810 20.640 1757.130 20.700 ;
        RECT 1759.110 20.640 1759.430 20.700 ;
        RECT 1756.810 20.500 1759.430 20.640 ;
        RECT 1756.810 20.440 1757.130 20.500 ;
        RECT 1759.110 20.440 1759.430 20.500 ;
      LAYER via ;
        RECT 1759.140 1685.420 1759.400 1685.680 ;
        RECT 1872.300 1685.420 1872.560 1685.680 ;
        RECT 1756.840 20.440 1757.100 20.700 ;
        RECT 1759.140 20.440 1759.400 20.700 ;
      LAYER met2 ;
        RECT 1872.225 1700.000 1872.505 1704.000 ;
        RECT 1872.360 1685.710 1872.500 1700.000 ;
        RECT 1759.140 1685.390 1759.400 1685.710 ;
        RECT 1872.300 1685.390 1872.560 1685.710 ;
        RECT 1759.200 20.730 1759.340 1685.390 ;
        RECT 1756.840 20.410 1757.100 20.730 ;
        RECT 1759.140 20.410 1759.400 20.730 ;
        RECT 1756.900 2.400 1757.040 20.410 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1819.905 1686.145 1820.075 1688.355 ;
      LAYER mcon ;
        RECT 1819.905 1688.185 1820.075 1688.355 ;
      LAYER met1 ;
        RECT 1879.630 1688.680 1879.950 1688.740 ;
        RECT 1862.240 1688.540 1879.950 1688.680 ;
        RECT 1819.845 1688.340 1820.135 1688.385 ;
        RECT 1862.240 1688.340 1862.380 1688.540 ;
        RECT 1879.630 1688.480 1879.950 1688.540 ;
        RECT 1819.845 1688.200 1862.380 1688.340 ;
        RECT 1819.845 1688.155 1820.135 1688.200 ;
        RECT 1779.810 1686.300 1780.130 1686.360 ;
        RECT 1819.845 1686.300 1820.135 1686.345 ;
        RECT 1779.810 1686.160 1820.135 1686.300 ;
        RECT 1779.810 1686.100 1780.130 1686.160 ;
        RECT 1819.845 1686.115 1820.135 1686.160 ;
        RECT 1774.750 14.860 1775.070 14.920 ;
        RECT 1779.810 14.860 1780.130 14.920 ;
        RECT 1774.750 14.720 1780.130 14.860 ;
        RECT 1774.750 14.660 1775.070 14.720 ;
        RECT 1779.810 14.660 1780.130 14.720 ;
      LAYER via ;
        RECT 1879.660 1688.480 1879.920 1688.740 ;
        RECT 1779.840 1686.100 1780.100 1686.360 ;
        RECT 1774.780 14.660 1775.040 14.920 ;
        RECT 1779.840 14.660 1780.100 14.920 ;
      LAYER met2 ;
        RECT 1879.585 1700.000 1879.865 1704.000 ;
        RECT 1879.720 1688.770 1879.860 1700.000 ;
        RECT 1879.660 1688.450 1879.920 1688.770 ;
        RECT 1779.840 1686.070 1780.100 1686.390 ;
        RECT 1779.900 14.950 1780.040 1686.070 ;
        RECT 1774.780 14.630 1775.040 14.950 ;
        RECT 1779.840 14.630 1780.100 14.950 ;
        RECT 1774.840 2.400 1774.980 14.630 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1793.610 1689.020 1793.930 1689.080 ;
        RECT 1886.990 1689.020 1887.310 1689.080 ;
        RECT 1793.610 1688.880 1804.420 1689.020 ;
        RECT 1793.610 1688.820 1793.930 1688.880 ;
        RECT 1804.280 1688.340 1804.420 1688.880 ;
        RECT 1861.780 1688.880 1887.310 1689.020 ;
        RECT 1861.780 1688.680 1861.920 1688.880 ;
        RECT 1886.990 1688.820 1887.310 1688.880 ;
        RECT 1819.460 1688.540 1861.920 1688.680 ;
        RECT 1819.460 1688.340 1819.600 1688.540 ;
        RECT 1804.280 1688.200 1819.600 1688.340 ;
        RECT 1792.690 2.960 1793.010 3.020 ;
        RECT 1793.610 2.960 1793.930 3.020 ;
        RECT 1792.690 2.820 1793.930 2.960 ;
        RECT 1792.690 2.760 1793.010 2.820 ;
        RECT 1793.610 2.760 1793.930 2.820 ;
      LAYER via ;
        RECT 1793.640 1688.820 1793.900 1689.080 ;
        RECT 1887.020 1688.820 1887.280 1689.080 ;
        RECT 1792.720 2.760 1792.980 3.020 ;
        RECT 1793.640 2.760 1793.900 3.020 ;
      LAYER met2 ;
        RECT 1886.945 1700.000 1887.225 1704.000 ;
        RECT 1887.080 1689.110 1887.220 1700.000 ;
        RECT 1793.640 1688.790 1793.900 1689.110 ;
        RECT 1887.020 1688.790 1887.280 1689.110 ;
        RECT 1793.700 3.050 1793.840 1688.790 ;
        RECT 1792.720 2.730 1792.980 3.050 ;
        RECT 1793.640 2.730 1793.900 3.050 ;
        RECT 1792.780 2.400 1792.920 2.730 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1861.305 1688.865 1861.475 1690.395 ;
      LAYER mcon ;
        RECT 1861.305 1690.225 1861.475 1690.395 ;
      LAYER met1 ;
        RECT 1861.245 1690.380 1861.535 1690.425 ;
        RECT 1894.350 1690.380 1894.670 1690.440 ;
        RECT 1861.245 1690.240 1894.670 1690.380 ;
        RECT 1861.245 1690.195 1861.535 1690.240 ;
        RECT 1894.350 1690.180 1894.670 1690.240 ;
        RECT 1814.310 1689.020 1814.630 1689.080 ;
        RECT 1861.245 1689.020 1861.535 1689.065 ;
        RECT 1814.310 1688.880 1861.535 1689.020 ;
        RECT 1814.310 1688.820 1814.630 1688.880 ;
        RECT 1861.245 1688.835 1861.535 1688.880 ;
        RECT 1810.630 20.640 1810.950 20.700 ;
        RECT 1814.310 20.640 1814.630 20.700 ;
        RECT 1810.630 20.500 1814.630 20.640 ;
        RECT 1810.630 20.440 1810.950 20.500 ;
        RECT 1814.310 20.440 1814.630 20.500 ;
      LAYER via ;
        RECT 1894.380 1690.180 1894.640 1690.440 ;
        RECT 1814.340 1688.820 1814.600 1689.080 ;
        RECT 1810.660 20.440 1810.920 20.700 ;
        RECT 1814.340 20.440 1814.600 20.700 ;
      LAYER met2 ;
        RECT 1894.305 1700.000 1894.585 1704.000 ;
        RECT 1894.440 1690.470 1894.580 1700.000 ;
        RECT 1894.380 1690.150 1894.640 1690.470 ;
        RECT 1814.340 1688.790 1814.600 1689.110 ;
        RECT 1814.400 20.730 1814.540 1688.790 ;
        RECT 1810.660 20.410 1810.920 20.730 ;
        RECT 1814.340 20.410 1814.600 20.730 ;
        RECT 1810.720 2.400 1810.860 20.410 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1834.625 435.285 1834.795 436.135 ;
      LAYER mcon ;
        RECT 1834.625 435.965 1834.795 436.135 ;
      LAYER met1 ;
        RECT 1834.550 1686.640 1834.870 1686.700 ;
        RECT 1901.710 1686.640 1902.030 1686.700 ;
        RECT 1834.550 1686.500 1902.030 1686.640 ;
        RECT 1834.550 1686.440 1834.870 1686.500 ;
        RECT 1901.710 1686.440 1902.030 1686.500 ;
        RECT 1834.090 1256.540 1834.410 1256.600 ;
        RECT 1834.090 1256.400 1834.780 1256.540 ;
        RECT 1834.090 1256.340 1834.410 1256.400 ;
        RECT 1834.640 1256.260 1834.780 1256.400 ;
        RECT 1834.550 1256.000 1834.870 1256.260 ;
        RECT 1834.550 436.120 1834.870 436.180 ;
        RECT 1834.355 435.980 1834.870 436.120 ;
        RECT 1834.550 435.920 1834.870 435.980 ;
        RECT 1834.550 435.440 1834.870 435.500 ;
        RECT 1834.355 435.300 1834.870 435.440 ;
        RECT 1834.550 435.240 1834.870 435.300 ;
        RECT 1834.550 193.500 1834.870 193.760 ;
        RECT 1834.640 193.080 1834.780 193.500 ;
        RECT 1834.550 192.820 1834.870 193.080 ;
        RECT 1834.550 62.260 1834.870 62.520 ;
        RECT 1834.640 61.840 1834.780 62.260 ;
        RECT 1834.550 61.580 1834.870 61.840 ;
        RECT 1828.570 23.360 1828.890 23.420 ;
        RECT 1834.550 23.360 1834.870 23.420 ;
        RECT 1828.570 23.220 1834.870 23.360 ;
        RECT 1828.570 23.160 1828.890 23.220 ;
        RECT 1834.550 23.160 1834.870 23.220 ;
      LAYER via ;
        RECT 1834.580 1686.440 1834.840 1686.700 ;
        RECT 1901.740 1686.440 1902.000 1686.700 ;
        RECT 1834.120 1256.340 1834.380 1256.600 ;
        RECT 1834.580 1256.000 1834.840 1256.260 ;
        RECT 1834.580 435.920 1834.840 436.180 ;
        RECT 1834.580 435.240 1834.840 435.500 ;
        RECT 1834.580 193.500 1834.840 193.760 ;
        RECT 1834.580 192.820 1834.840 193.080 ;
        RECT 1834.580 62.260 1834.840 62.520 ;
        RECT 1834.580 61.580 1834.840 61.840 ;
        RECT 1828.600 23.160 1828.860 23.420 ;
        RECT 1834.580 23.160 1834.840 23.420 ;
      LAYER met2 ;
        RECT 1901.665 1700.000 1901.945 1704.000 ;
        RECT 1901.800 1686.730 1901.940 1700.000 ;
        RECT 1834.580 1686.410 1834.840 1686.730 ;
        RECT 1901.740 1686.410 1902.000 1686.730 ;
        RECT 1834.640 1257.730 1834.780 1686.410 ;
        RECT 1834.180 1257.590 1834.780 1257.730 ;
        RECT 1834.180 1256.630 1834.320 1257.590 ;
        RECT 1834.120 1256.310 1834.380 1256.630 ;
        RECT 1834.580 1255.970 1834.840 1256.290 ;
        RECT 1834.640 436.210 1834.780 1255.970 ;
        RECT 1834.580 435.890 1834.840 436.210 ;
        RECT 1834.580 435.210 1834.840 435.530 ;
        RECT 1834.640 242.605 1834.780 435.210 ;
        RECT 1834.570 242.235 1834.850 242.605 ;
        RECT 1834.570 241.555 1834.850 241.925 ;
        RECT 1834.640 193.790 1834.780 241.555 ;
        RECT 1834.580 193.470 1834.840 193.790 ;
        RECT 1834.580 192.790 1834.840 193.110 ;
        RECT 1834.640 62.550 1834.780 192.790 ;
        RECT 1834.580 62.230 1834.840 62.550 ;
        RECT 1834.580 61.550 1834.840 61.870 ;
        RECT 1834.640 23.450 1834.780 61.550 ;
        RECT 1828.600 23.130 1828.860 23.450 ;
        RECT 1834.580 23.130 1834.840 23.450 ;
        RECT 1828.660 2.400 1828.800 23.130 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
      LAYER via2 ;
        RECT 1834.570 242.280 1834.850 242.560 ;
        RECT 1834.570 241.600 1834.850 241.880 ;
      LAYER met3 ;
        RECT 1834.545 242.570 1834.875 242.585 ;
        RECT 1834.545 242.255 1835.090 242.570 ;
        RECT 1834.790 241.905 1835.090 242.255 ;
        RECT 1834.545 241.590 1835.090 241.905 ;
        RECT 1834.545 241.575 1834.875 241.590 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1909.070 1688.340 1909.390 1688.400 ;
        RECT 1869.140 1688.200 1909.390 1688.340 ;
        RECT 1848.810 1686.980 1849.130 1687.040 ;
        RECT 1869.140 1686.980 1869.280 1688.200 ;
        RECT 1909.070 1688.140 1909.390 1688.200 ;
        RECT 1848.810 1686.840 1869.280 1686.980 ;
        RECT 1848.810 1686.780 1849.130 1686.840 ;
        RECT 1846.050 20.640 1846.370 20.700 ;
        RECT 1848.810 20.640 1849.130 20.700 ;
        RECT 1846.050 20.500 1849.130 20.640 ;
        RECT 1846.050 20.440 1846.370 20.500 ;
        RECT 1848.810 20.440 1849.130 20.500 ;
      LAYER via ;
        RECT 1848.840 1686.780 1849.100 1687.040 ;
        RECT 1909.100 1688.140 1909.360 1688.400 ;
        RECT 1846.080 20.440 1846.340 20.700 ;
        RECT 1848.840 20.440 1849.100 20.700 ;
      LAYER met2 ;
        RECT 1909.025 1700.000 1909.305 1704.000 ;
        RECT 1909.160 1688.430 1909.300 1700.000 ;
        RECT 1909.100 1688.110 1909.360 1688.430 ;
        RECT 1848.840 1686.750 1849.100 1687.070 ;
        RECT 1848.900 20.730 1849.040 1686.750 ;
        RECT 1846.080 20.410 1846.340 20.730 ;
        RECT 1848.840 20.410 1849.100 20.730 ;
        RECT 1846.140 2.400 1846.280 20.410 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1869.510 1688.000 1869.830 1688.060 ;
        RECT 1916.430 1688.000 1916.750 1688.060 ;
        RECT 1869.510 1687.860 1916.750 1688.000 ;
        RECT 1869.510 1687.800 1869.830 1687.860 ;
        RECT 1916.430 1687.800 1916.750 1687.860 ;
        RECT 1863.990 19.280 1864.310 19.340 ;
        RECT 1869.510 19.280 1869.830 19.340 ;
        RECT 1863.990 19.140 1869.830 19.280 ;
        RECT 1863.990 19.080 1864.310 19.140 ;
        RECT 1869.510 19.080 1869.830 19.140 ;
      LAYER via ;
        RECT 1869.540 1687.800 1869.800 1688.060 ;
        RECT 1916.460 1687.800 1916.720 1688.060 ;
        RECT 1864.020 19.080 1864.280 19.340 ;
        RECT 1869.540 19.080 1869.800 19.340 ;
      LAYER met2 ;
        RECT 1916.385 1700.000 1916.665 1704.000 ;
        RECT 1916.520 1688.090 1916.660 1700.000 ;
        RECT 1869.540 1687.770 1869.800 1688.090 ;
        RECT 1916.460 1687.770 1916.720 1688.090 ;
        RECT 1869.600 19.370 1869.740 1687.770 ;
        RECT 1864.020 19.050 1864.280 19.370 ;
        RECT 1869.540 19.050 1869.800 19.370 ;
        RECT 1864.080 2.400 1864.220 19.050 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1450.985 1055.445 1451.155 1097.095 ;
        RECT 1450.065 952.425 1450.235 1000.535 ;
        RECT 1450.065 862.665 1450.235 910.775 ;
        RECT 1450.065 520.965 1450.235 558.875 ;
        RECT 1450.065 468.945 1450.235 489.855 ;
      LAYER mcon ;
        RECT 1450.985 1096.925 1451.155 1097.095 ;
        RECT 1450.065 1000.365 1450.235 1000.535 ;
        RECT 1450.065 910.605 1450.235 910.775 ;
        RECT 1450.065 558.705 1450.235 558.875 ;
        RECT 1450.065 489.685 1450.235 489.855 ;
      LAYER met1 ;
        RECT 1450.450 1587.020 1450.770 1587.080 ;
        RECT 1450.910 1587.020 1451.230 1587.080 ;
        RECT 1450.450 1586.880 1451.230 1587.020 ;
        RECT 1450.450 1586.820 1450.770 1586.880 ;
        RECT 1450.910 1586.820 1451.230 1586.880 ;
        RECT 1449.990 1473.120 1450.310 1473.180 ;
        RECT 1450.910 1473.120 1451.230 1473.180 ;
        RECT 1449.990 1472.980 1451.230 1473.120 ;
        RECT 1449.990 1472.920 1450.310 1472.980 ;
        RECT 1450.910 1472.920 1451.230 1472.980 ;
        RECT 1449.990 1448.980 1450.310 1449.040 ;
        RECT 1450.910 1448.980 1451.230 1449.040 ;
        RECT 1449.990 1448.840 1451.230 1448.980 ;
        RECT 1449.990 1448.780 1450.310 1448.840 ;
        RECT 1450.910 1448.780 1451.230 1448.840 ;
        RECT 1450.450 1345.620 1450.770 1345.680 ;
        RECT 1450.910 1345.620 1451.230 1345.680 ;
        RECT 1450.450 1345.480 1451.230 1345.620 ;
        RECT 1450.450 1345.420 1450.770 1345.480 ;
        RECT 1450.910 1345.420 1451.230 1345.480 ;
        RECT 1449.990 1256.200 1450.310 1256.260 ;
        RECT 1450.450 1256.200 1450.770 1256.260 ;
        RECT 1449.990 1256.060 1450.770 1256.200 ;
        RECT 1449.990 1256.000 1450.310 1256.060 ;
        RECT 1450.450 1256.000 1450.770 1256.060 ;
        RECT 1449.990 1207.580 1450.310 1207.640 ;
        RECT 1450.910 1207.580 1451.230 1207.640 ;
        RECT 1449.990 1207.440 1451.230 1207.580 ;
        RECT 1449.990 1207.380 1450.310 1207.440 ;
        RECT 1450.910 1207.380 1451.230 1207.440 ;
        RECT 1451.830 1104.560 1452.150 1104.620 ;
        RECT 1451.000 1104.420 1452.150 1104.560 ;
        RECT 1451.000 1104.280 1451.140 1104.420 ;
        RECT 1451.830 1104.360 1452.150 1104.420 ;
        RECT 1450.910 1104.020 1451.230 1104.280 ;
        RECT 1450.910 1097.080 1451.230 1097.140 ;
        RECT 1450.715 1096.940 1451.230 1097.080 ;
        RECT 1450.910 1096.880 1451.230 1096.940 ;
        RECT 1450.910 1055.600 1451.230 1055.660 ;
        RECT 1450.715 1055.460 1451.230 1055.600 ;
        RECT 1450.910 1055.400 1451.230 1055.460 ;
        RECT 1450.005 1000.520 1450.295 1000.565 ;
        RECT 1450.910 1000.520 1451.230 1000.580 ;
        RECT 1450.005 1000.380 1451.230 1000.520 ;
        RECT 1450.005 1000.335 1450.295 1000.380 ;
        RECT 1450.910 1000.320 1451.230 1000.380 ;
        RECT 1449.990 952.580 1450.310 952.640 ;
        RECT 1449.795 952.440 1450.310 952.580 ;
        RECT 1449.990 952.380 1450.310 952.440 ;
        RECT 1449.990 941.500 1450.310 941.760 ;
        RECT 1450.080 941.080 1450.220 941.500 ;
        RECT 1449.990 940.820 1450.310 941.080 ;
        RECT 1449.990 910.760 1450.310 910.820 ;
        RECT 1449.795 910.620 1450.310 910.760 ;
        RECT 1449.990 910.560 1450.310 910.620 ;
        RECT 1449.990 862.820 1450.310 862.880 ;
        RECT 1449.795 862.680 1450.310 862.820 ;
        RECT 1449.990 862.620 1450.310 862.680 ;
        RECT 1449.990 765.920 1450.310 765.980 ;
        RECT 1450.450 765.920 1450.770 765.980 ;
        RECT 1449.990 765.780 1450.770 765.920 ;
        RECT 1449.990 765.720 1450.310 765.780 ;
        RECT 1450.450 765.720 1450.770 765.780 ;
        RECT 1449.530 662.560 1449.850 662.620 ;
        RECT 1450.450 662.560 1450.770 662.620 ;
        RECT 1449.530 662.420 1450.770 662.560 ;
        RECT 1449.530 662.360 1449.850 662.420 ;
        RECT 1450.450 662.360 1450.770 662.420 ;
        RECT 1449.530 621.080 1449.850 621.140 ;
        RECT 1449.990 621.080 1450.310 621.140 ;
        RECT 1449.530 620.940 1450.310 621.080 ;
        RECT 1449.530 620.880 1449.850 620.940 ;
        RECT 1449.990 620.880 1450.310 620.940 ;
        RECT 1450.005 558.860 1450.295 558.905 ;
        RECT 1450.450 558.860 1450.770 558.920 ;
        RECT 1450.005 558.720 1450.770 558.860 ;
        RECT 1450.005 558.675 1450.295 558.720 ;
        RECT 1450.450 558.660 1450.770 558.720 ;
        RECT 1449.990 521.120 1450.310 521.180 ;
        RECT 1449.795 520.980 1450.310 521.120 ;
        RECT 1449.990 520.920 1450.310 520.980 ;
        RECT 1449.990 489.840 1450.310 489.900 ;
        RECT 1449.795 489.700 1450.310 489.840 ;
        RECT 1449.990 489.640 1450.310 489.700 ;
        RECT 1449.990 469.100 1450.310 469.160 ;
        RECT 1449.795 468.960 1450.310 469.100 ;
        RECT 1449.990 468.900 1450.310 468.960 ;
        RECT 1450.450 420.960 1450.770 421.220 ;
        RECT 1450.540 420.480 1450.680 420.960 ;
        RECT 1450.910 420.480 1451.230 420.540 ;
        RECT 1450.540 420.340 1451.230 420.480 ;
        RECT 1450.910 420.280 1451.230 420.340 ;
        RECT 744.810 60.420 745.130 60.480 ;
        RECT 1449.990 60.420 1450.310 60.480 ;
        RECT 744.810 60.280 1450.310 60.420 ;
        RECT 744.810 60.220 745.130 60.280 ;
        RECT 1449.990 60.220 1450.310 60.280 ;
      LAYER via ;
        RECT 1450.480 1586.820 1450.740 1587.080 ;
        RECT 1450.940 1586.820 1451.200 1587.080 ;
        RECT 1450.020 1472.920 1450.280 1473.180 ;
        RECT 1450.940 1472.920 1451.200 1473.180 ;
        RECT 1450.020 1448.780 1450.280 1449.040 ;
        RECT 1450.940 1448.780 1451.200 1449.040 ;
        RECT 1450.480 1345.420 1450.740 1345.680 ;
        RECT 1450.940 1345.420 1451.200 1345.680 ;
        RECT 1450.020 1256.000 1450.280 1256.260 ;
        RECT 1450.480 1256.000 1450.740 1256.260 ;
        RECT 1450.020 1207.380 1450.280 1207.640 ;
        RECT 1450.940 1207.380 1451.200 1207.640 ;
        RECT 1451.860 1104.360 1452.120 1104.620 ;
        RECT 1450.940 1104.020 1451.200 1104.280 ;
        RECT 1450.940 1096.880 1451.200 1097.140 ;
        RECT 1450.940 1055.400 1451.200 1055.660 ;
        RECT 1450.940 1000.320 1451.200 1000.580 ;
        RECT 1450.020 952.380 1450.280 952.640 ;
        RECT 1450.020 941.500 1450.280 941.760 ;
        RECT 1450.020 940.820 1450.280 941.080 ;
        RECT 1450.020 910.560 1450.280 910.820 ;
        RECT 1450.020 862.620 1450.280 862.880 ;
        RECT 1450.020 765.720 1450.280 765.980 ;
        RECT 1450.480 765.720 1450.740 765.980 ;
        RECT 1449.560 662.360 1449.820 662.620 ;
        RECT 1450.480 662.360 1450.740 662.620 ;
        RECT 1449.560 620.880 1449.820 621.140 ;
        RECT 1450.020 620.880 1450.280 621.140 ;
        RECT 1450.480 558.660 1450.740 558.920 ;
        RECT 1450.020 520.920 1450.280 521.180 ;
        RECT 1450.020 489.640 1450.280 489.900 ;
        RECT 1450.020 468.900 1450.280 469.160 ;
        RECT 1450.480 420.960 1450.740 421.220 ;
        RECT 1450.940 420.280 1451.200 420.540 ;
        RECT 744.840 60.220 745.100 60.480 ;
        RECT 1450.020 60.220 1450.280 60.480 ;
      LAYER met2 ;
        RECT 1453.625 1701.090 1453.905 1704.000 ;
        RECT 1451.460 1700.950 1453.905 1701.090 ;
        RECT 1451.460 1677.970 1451.600 1700.950 ;
        RECT 1453.625 1700.000 1453.905 1700.950 ;
        RECT 1450.540 1677.830 1451.600 1677.970 ;
        RECT 1450.540 1587.110 1450.680 1677.830 ;
        RECT 1450.480 1586.790 1450.740 1587.110 ;
        RECT 1450.940 1586.790 1451.200 1587.110 ;
        RECT 1451.000 1473.210 1451.140 1586.790 ;
        RECT 1450.020 1472.890 1450.280 1473.210 ;
        RECT 1450.940 1472.890 1451.200 1473.210 ;
        RECT 1450.080 1449.070 1450.220 1472.890 ;
        RECT 1450.020 1448.750 1450.280 1449.070 ;
        RECT 1450.940 1448.750 1451.200 1449.070 ;
        RECT 1451.000 1345.710 1451.140 1448.750 ;
        RECT 1450.480 1345.390 1450.740 1345.710 ;
        RECT 1450.940 1345.390 1451.200 1345.710 ;
        RECT 1450.540 1256.290 1450.680 1345.390 ;
        RECT 1450.020 1255.970 1450.280 1256.290 ;
        RECT 1450.480 1255.970 1450.740 1256.290 ;
        RECT 1450.080 1207.670 1450.220 1255.970 ;
        RECT 1450.020 1207.350 1450.280 1207.670 ;
        RECT 1450.940 1207.350 1451.200 1207.670 ;
        RECT 1451.000 1176.810 1451.140 1207.350 ;
        RECT 1451.000 1176.670 1452.060 1176.810 ;
        RECT 1451.920 1104.650 1452.060 1176.670 ;
        RECT 1451.860 1104.330 1452.120 1104.650 ;
        RECT 1450.940 1104.165 1451.200 1104.310 ;
        RECT 1450.930 1103.795 1451.210 1104.165 ;
        RECT 1450.930 1103.115 1451.210 1103.485 ;
        RECT 1451.000 1097.170 1451.140 1103.115 ;
        RECT 1450.940 1096.850 1451.200 1097.170 ;
        RECT 1450.940 1055.370 1451.200 1055.690 ;
        RECT 1451.000 1048.970 1451.140 1055.370 ;
        RECT 1451.000 1048.830 1451.600 1048.970 ;
        RECT 1451.460 1021.090 1451.600 1048.830 ;
        RECT 1451.000 1020.950 1451.600 1021.090 ;
        RECT 1451.000 1000.610 1451.140 1020.950 ;
        RECT 1450.940 1000.290 1451.200 1000.610 ;
        RECT 1450.020 952.350 1450.280 952.670 ;
        RECT 1450.080 941.790 1450.220 952.350 ;
        RECT 1450.020 941.470 1450.280 941.790 ;
        RECT 1450.020 940.790 1450.280 941.110 ;
        RECT 1450.080 910.850 1450.220 940.790 ;
        RECT 1450.020 910.530 1450.280 910.850 ;
        RECT 1450.020 862.590 1450.280 862.910 ;
        RECT 1450.080 766.010 1450.220 862.590 ;
        RECT 1450.020 765.690 1450.280 766.010 ;
        RECT 1450.480 765.690 1450.740 766.010 ;
        RECT 1450.540 662.650 1450.680 765.690 ;
        RECT 1449.560 662.330 1449.820 662.650 ;
        RECT 1450.480 662.330 1450.740 662.650 ;
        RECT 1449.620 621.170 1449.760 662.330 ;
        RECT 1449.560 620.850 1449.820 621.170 ;
        RECT 1450.020 620.850 1450.280 621.170 ;
        RECT 1450.080 599.490 1450.220 620.850 ;
        RECT 1449.620 599.350 1450.220 599.490 ;
        RECT 1449.620 572.290 1449.760 599.350 ;
        RECT 1449.620 572.150 1450.680 572.290 ;
        RECT 1450.540 558.950 1450.680 572.150 ;
        RECT 1450.480 558.630 1450.740 558.950 ;
        RECT 1450.020 520.890 1450.280 521.210 ;
        RECT 1450.080 489.930 1450.220 520.890 ;
        RECT 1450.020 489.610 1450.280 489.930 ;
        RECT 1450.020 468.870 1450.280 469.190 ;
        RECT 1450.080 441.730 1450.220 468.870 ;
        RECT 1450.080 441.590 1450.680 441.730 ;
        RECT 1450.540 421.250 1450.680 441.590 ;
        RECT 1450.480 420.930 1450.740 421.250 ;
        RECT 1450.940 420.250 1451.200 420.570 ;
        RECT 1451.000 303.805 1451.140 420.250 ;
        RECT 1450.010 303.435 1450.290 303.805 ;
        RECT 1450.930 303.435 1451.210 303.805 ;
        RECT 1450.080 60.510 1450.220 303.435 ;
        RECT 744.840 60.190 745.100 60.510 ;
        RECT 1450.020 60.190 1450.280 60.510 ;
        RECT 744.900 17.410 745.040 60.190 ;
        RECT 740.300 17.270 745.040 17.410 ;
        RECT 740.300 2.400 740.440 17.270 ;
        RECT 740.090 -4.800 740.650 2.400 ;
      LAYER via2 ;
        RECT 1450.930 1103.840 1451.210 1104.120 ;
        RECT 1450.930 1103.160 1451.210 1103.440 ;
        RECT 1450.010 303.480 1450.290 303.760 ;
        RECT 1450.930 303.480 1451.210 303.760 ;
      LAYER met3 ;
        RECT 1450.905 1104.130 1451.235 1104.145 ;
        RECT 1450.905 1103.815 1451.450 1104.130 ;
        RECT 1451.150 1103.465 1451.450 1103.815 ;
        RECT 1450.905 1103.150 1451.450 1103.465 ;
        RECT 1450.905 1103.135 1451.235 1103.150 ;
        RECT 1449.985 303.770 1450.315 303.785 ;
        RECT 1450.905 303.770 1451.235 303.785 ;
        RECT 1449.985 303.470 1451.235 303.770 ;
        RECT 1449.985 303.455 1450.315 303.470 ;
        RECT 1450.905 303.455 1451.235 303.470 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1908.150 1684.260 1908.470 1684.320 ;
        RECT 1923.790 1684.260 1924.110 1684.320 ;
        RECT 1908.150 1684.120 1924.110 1684.260 ;
        RECT 1908.150 1684.060 1908.470 1684.120 ;
        RECT 1923.790 1684.060 1924.110 1684.120 ;
        RECT 1881.930 15.200 1882.250 15.260 ;
        RECT 1908.150 15.200 1908.470 15.260 ;
        RECT 1881.930 15.060 1908.470 15.200 ;
        RECT 1881.930 15.000 1882.250 15.060 ;
        RECT 1908.150 15.000 1908.470 15.060 ;
      LAYER via ;
        RECT 1908.180 1684.060 1908.440 1684.320 ;
        RECT 1923.820 1684.060 1924.080 1684.320 ;
        RECT 1881.960 15.000 1882.220 15.260 ;
        RECT 1908.180 15.000 1908.440 15.260 ;
      LAYER met2 ;
        RECT 1923.745 1700.000 1924.025 1704.000 ;
        RECT 1923.880 1684.350 1924.020 1700.000 ;
        RECT 1908.180 1684.030 1908.440 1684.350 ;
        RECT 1923.820 1684.030 1924.080 1684.350 ;
        RECT 1908.240 15.290 1908.380 1684.030 ;
        RECT 1881.960 14.970 1882.220 15.290 ;
        RECT 1908.180 14.970 1908.440 15.290 ;
        RECT 1882.020 2.400 1882.160 14.970 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1904.010 1684.600 1904.330 1684.660 ;
        RECT 1931.150 1684.600 1931.470 1684.660 ;
        RECT 1904.010 1684.460 1931.470 1684.600 ;
        RECT 1904.010 1684.400 1904.330 1684.460 ;
        RECT 1931.150 1684.400 1931.470 1684.460 ;
        RECT 1899.870 17.580 1900.190 17.640 ;
        RECT 1904.010 17.580 1904.330 17.640 ;
        RECT 1899.870 17.440 1904.330 17.580 ;
        RECT 1899.870 17.380 1900.190 17.440 ;
        RECT 1904.010 17.380 1904.330 17.440 ;
      LAYER via ;
        RECT 1904.040 1684.400 1904.300 1684.660 ;
        RECT 1931.180 1684.400 1931.440 1684.660 ;
        RECT 1899.900 17.380 1900.160 17.640 ;
        RECT 1904.040 17.380 1904.300 17.640 ;
      LAYER met2 ;
        RECT 1931.105 1700.000 1931.385 1704.000 ;
        RECT 1931.240 1684.690 1931.380 1700.000 ;
        RECT 1904.040 1684.370 1904.300 1684.690 ;
        RECT 1931.180 1684.370 1931.440 1684.690 ;
        RECT 1904.100 17.670 1904.240 1684.370 ;
        RECT 1899.900 17.350 1900.160 17.670 ;
        RECT 1904.040 17.350 1904.300 17.670 ;
        RECT 1899.960 2.400 1900.100 17.350 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1921.490 1688.340 1921.810 1688.400 ;
        RECT 1938.510 1688.340 1938.830 1688.400 ;
        RECT 1921.490 1688.200 1938.830 1688.340 ;
        RECT 1921.490 1688.140 1921.810 1688.200 ;
        RECT 1938.510 1688.140 1938.830 1688.200 ;
        RECT 1917.810 20.300 1918.130 20.360 ;
        RECT 1921.490 20.300 1921.810 20.360 ;
        RECT 1917.810 20.160 1921.810 20.300 ;
        RECT 1917.810 20.100 1918.130 20.160 ;
        RECT 1921.490 20.100 1921.810 20.160 ;
      LAYER via ;
        RECT 1921.520 1688.140 1921.780 1688.400 ;
        RECT 1938.540 1688.140 1938.800 1688.400 ;
        RECT 1917.840 20.100 1918.100 20.360 ;
        RECT 1921.520 20.100 1921.780 20.360 ;
      LAYER met2 ;
        RECT 1938.465 1700.000 1938.745 1704.000 ;
        RECT 1938.600 1688.430 1938.740 1700.000 ;
        RECT 1921.520 1688.110 1921.780 1688.430 ;
        RECT 1938.540 1688.110 1938.800 1688.430 ;
        RECT 1921.580 20.390 1921.720 1688.110 ;
        RECT 1917.840 20.070 1918.100 20.390 ;
        RECT 1921.520 20.070 1921.780 20.390 ;
        RECT 1917.900 2.400 1918.040 20.070 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1942.190 1689.360 1942.510 1689.420 ;
        RECT 1945.870 1689.360 1946.190 1689.420 ;
        RECT 1942.190 1689.220 1946.190 1689.360 ;
        RECT 1942.190 1689.160 1942.510 1689.220 ;
        RECT 1945.870 1689.160 1946.190 1689.220 ;
        RECT 1942.190 14.180 1942.510 14.240 ;
        RECT 1935.380 14.040 1942.510 14.180 ;
        RECT 1935.380 13.900 1935.520 14.040 ;
        RECT 1942.190 13.980 1942.510 14.040 ;
        RECT 1935.290 13.640 1935.610 13.900 ;
      LAYER via ;
        RECT 1942.220 1689.160 1942.480 1689.420 ;
        RECT 1945.900 1689.160 1946.160 1689.420 ;
        RECT 1942.220 13.980 1942.480 14.240 ;
        RECT 1935.320 13.640 1935.580 13.900 ;
      LAYER met2 ;
        RECT 1945.825 1700.000 1946.105 1704.000 ;
        RECT 1945.960 1689.450 1946.100 1700.000 ;
        RECT 1942.220 1689.130 1942.480 1689.450 ;
        RECT 1945.900 1689.130 1946.160 1689.450 ;
        RECT 1942.280 14.270 1942.420 1689.130 ;
        RECT 1942.220 13.950 1942.480 14.270 ;
        RECT 1935.320 13.610 1935.580 13.930 ;
        RECT 1935.380 2.400 1935.520 13.610 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1953.185 1700.410 1953.465 1704.000 ;
        RECT 1952.860 1700.270 1953.465 1700.410 ;
        RECT 1952.860 7.210 1953.000 1700.270 ;
        RECT 1953.185 1700.000 1953.465 1700.270 ;
        RECT 1952.860 7.070 1953.460 7.210 ;
        RECT 1953.320 2.400 1953.460 7.070 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1968.025 1538.925 1968.195 1587.035 ;
        RECT 1968.025 1400.885 1968.195 1490.475 ;
        RECT 1968.025 1304.325 1968.195 1393.575 ;
        RECT 1967.565 965.345 1967.735 1024.675 ;
        RECT 1967.565 917.405 1967.735 959.055 ;
        RECT 1968.025 766.105 1968.195 814.215 ;
        RECT 1968.025 710.685 1968.195 742.475 ;
        RECT 1968.025 552.245 1968.195 600.355 ;
        RECT 1968.025 434.265 1968.195 503.455 ;
        RECT 1968.485 324.445 1968.655 372.555 ;
        RECT 1968.025 138.125 1968.195 186.235 ;
        RECT 1971.245 2.805 1971.415 5.355 ;
      LAYER mcon ;
        RECT 1968.025 1586.865 1968.195 1587.035 ;
        RECT 1968.025 1490.305 1968.195 1490.475 ;
        RECT 1968.025 1393.405 1968.195 1393.575 ;
        RECT 1967.565 1024.505 1967.735 1024.675 ;
        RECT 1967.565 958.885 1967.735 959.055 ;
        RECT 1968.025 814.045 1968.195 814.215 ;
        RECT 1968.025 742.305 1968.195 742.475 ;
        RECT 1968.025 600.185 1968.195 600.355 ;
        RECT 1968.025 503.285 1968.195 503.455 ;
        RECT 1968.485 372.385 1968.655 372.555 ;
        RECT 1968.025 186.065 1968.195 186.235 ;
        RECT 1971.245 5.185 1971.415 5.355 ;
      LAYER met1 ;
        RECT 1960.590 1684.600 1960.910 1684.660 ;
        RECT 1967.950 1684.600 1968.270 1684.660 ;
        RECT 1960.590 1684.460 1968.270 1684.600 ;
        RECT 1960.590 1684.400 1960.910 1684.460 ;
        RECT 1967.950 1684.400 1968.270 1684.460 ;
        RECT 1967.950 1642.100 1968.270 1642.160 ;
        RECT 1968.410 1642.100 1968.730 1642.160 ;
        RECT 1967.950 1641.960 1968.730 1642.100 ;
        RECT 1967.950 1641.900 1968.270 1641.960 ;
        RECT 1968.410 1641.900 1968.730 1641.960 ;
        RECT 1967.950 1587.020 1968.270 1587.080 ;
        RECT 1967.755 1586.880 1968.270 1587.020 ;
        RECT 1967.950 1586.820 1968.270 1586.880 ;
        RECT 1967.950 1539.080 1968.270 1539.140 ;
        RECT 1967.755 1538.940 1968.270 1539.080 ;
        RECT 1967.950 1538.880 1968.270 1538.940 ;
        RECT 1967.950 1490.460 1968.270 1490.520 ;
        RECT 1967.755 1490.320 1968.270 1490.460 ;
        RECT 1967.950 1490.260 1968.270 1490.320 ;
        RECT 1967.950 1401.040 1968.270 1401.100 ;
        RECT 1967.755 1400.900 1968.270 1401.040 ;
        RECT 1967.950 1400.840 1968.270 1400.900 ;
        RECT 1967.950 1393.560 1968.270 1393.620 ;
        RECT 1967.755 1393.420 1968.270 1393.560 ;
        RECT 1967.950 1393.360 1968.270 1393.420 ;
        RECT 1967.950 1304.480 1968.270 1304.540 ;
        RECT 1967.755 1304.340 1968.270 1304.480 ;
        RECT 1967.950 1304.280 1968.270 1304.340 ;
        RECT 1967.950 1249.060 1968.270 1249.120 ;
        RECT 1968.870 1249.060 1969.190 1249.120 ;
        RECT 1967.950 1248.920 1969.190 1249.060 ;
        RECT 1967.950 1248.860 1968.270 1248.920 ;
        RECT 1968.870 1248.860 1969.190 1248.920 ;
        RECT 1966.570 1193.640 1966.890 1193.700 ;
        RECT 1967.490 1193.640 1967.810 1193.700 ;
        RECT 1966.570 1193.500 1967.810 1193.640 ;
        RECT 1966.570 1193.440 1966.890 1193.500 ;
        RECT 1967.490 1193.440 1967.810 1193.500 ;
        RECT 1966.570 1121.220 1966.890 1121.280 ;
        RECT 1967.490 1121.220 1967.810 1121.280 ;
        RECT 1966.570 1121.080 1967.810 1121.220 ;
        RECT 1966.570 1121.020 1966.890 1121.080 ;
        RECT 1967.490 1121.020 1967.810 1121.080 ;
        RECT 1967.490 1024.660 1967.810 1024.720 ;
        RECT 1967.295 1024.520 1967.810 1024.660 ;
        RECT 1967.490 1024.460 1967.810 1024.520 ;
        RECT 1967.490 965.500 1967.810 965.560 ;
        RECT 1967.295 965.360 1967.810 965.500 ;
        RECT 1967.490 965.300 1967.810 965.360 ;
        RECT 1967.490 959.040 1967.810 959.100 ;
        RECT 1967.295 958.900 1967.810 959.040 ;
        RECT 1967.490 958.840 1967.810 958.900 ;
        RECT 1967.490 917.560 1967.810 917.620 ;
        RECT 1967.295 917.420 1967.810 917.560 ;
        RECT 1967.490 917.360 1967.810 917.420 ;
        RECT 1966.570 910.760 1966.890 910.820 ;
        RECT 1967.490 910.760 1967.810 910.820 ;
        RECT 1966.570 910.620 1967.810 910.760 ;
        RECT 1966.570 910.560 1966.890 910.620 ;
        RECT 1967.490 910.560 1967.810 910.620 ;
        RECT 1967.965 814.200 1968.255 814.245 ;
        RECT 1968.410 814.200 1968.730 814.260 ;
        RECT 1967.965 814.060 1968.730 814.200 ;
        RECT 1967.965 814.015 1968.255 814.060 ;
        RECT 1968.410 814.000 1968.730 814.060 ;
        RECT 1967.950 766.260 1968.270 766.320 ;
        RECT 1967.755 766.120 1968.270 766.260 ;
        RECT 1967.950 766.060 1968.270 766.120 ;
        RECT 1967.950 742.460 1968.270 742.520 ;
        RECT 1967.755 742.320 1968.270 742.460 ;
        RECT 1967.950 742.260 1968.270 742.320 ;
        RECT 1967.965 710.840 1968.255 710.885 ;
        RECT 1968.410 710.840 1968.730 710.900 ;
        RECT 1967.965 710.700 1968.730 710.840 ;
        RECT 1967.965 710.655 1968.255 710.700 ;
        RECT 1968.410 710.640 1968.730 710.700 ;
        RECT 1967.950 655.420 1968.270 655.480 ;
        RECT 1968.870 655.420 1969.190 655.480 ;
        RECT 1967.950 655.280 1969.190 655.420 ;
        RECT 1967.950 655.220 1968.270 655.280 ;
        RECT 1968.870 655.220 1969.190 655.280 ;
        RECT 1967.950 600.340 1968.270 600.400 ;
        RECT 1967.755 600.200 1968.270 600.340 ;
        RECT 1967.950 600.140 1968.270 600.200 ;
        RECT 1967.950 552.400 1968.270 552.460 ;
        RECT 1967.755 552.260 1968.270 552.400 ;
        RECT 1967.950 552.200 1968.270 552.260 ;
        RECT 1967.950 524.320 1968.270 524.580 ;
        RECT 1968.040 523.840 1968.180 524.320 ;
        RECT 1968.410 523.840 1968.730 523.900 ;
        RECT 1968.040 523.700 1968.730 523.840 ;
        RECT 1968.410 523.640 1968.730 523.700 ;
        RECT 1967.965 503.440 1968.255 503.485 ;
        RECT 1968.410 503.440 1968.730 503.500 ;
        RECT 1967.965 503.300 1968.730 503.440 ;
        RECT 1967.965 503.255 1968.255 503.300 ;
        RECT 1968.410 503.240 1968.730 503.300 ;
        RECT 1967.950 434.420 1968.270 434.480 ;
        RECT 1967.755 434.280 1968.270 434.420 ;
        RECT 1967.950 434.220 1968.270 434.280 ;
        RECT 1968.410 372.540 1968.730 372.600 ;
        RECT 1968.215 372.400 1968.730 372.540 ;
        RECT 1968.410 372.340 1968.730 372.400 ;
        RECT 1968.425 324.600 1968.715 324.645 ;
        RECT 1968.870 324.600 1969.190 324.660 ;
        RECT 1968.425 324.460 1969.190 324.600 ;
        RECT 1968.425 324.415 1968.715 324.460 ;
        RECT 1968.870 324.400 1969.190 324.460 ;
        RECT 1967.490 276.320 1967.810 276.380 ;
        RECT 1968.870 276.320 1969.190 276.380 ;
        RECT 1967.490 276.180 1969.190 276.320 ;
        RECT 1967.490 276.120 1967.810 276.180 ;
        RECT 1968.870 276.120 1969.190 276.180 ;
        RECT 1967.030 228.040 1967.350 228.100 ;
        RECT 1968.410 228.040 1968.730 228.100 ;
        RECT 1967.030 227.900 1968.730 228.040 ;
        RECT 1967.030 227.840 1967.350 227.900 ;
        RECT 1968.410 227.840 1968.730 227.900 ;
        RECT 1967.950 186.220 1968.270 186.280 ;
        RECT 1967.755 186.080 1968.270 186.220 ;
        RECT 1967.950 186.020 1968.270 186.080 ;
        RECT 1967.965 138.280 1968.255 138.325 ;
        RECT 1968.410 138.280 1968.730 138.340 ;
        RECT 1967.965 138.140 1968.730 138.280 ;
        RECT 1967.965 138.095 1968.255 138.140 ;
        RECT 1968.410 138.080 1968.730 138.140 ;
        RECT 1968.410 90.140 1968.730 90.400 ;
        RECT 1968.500 89.720 1968.640 90.140 ;
        RECT 1968.410 89.460 1968.730 89.720 ;
        RECT 1968.410 34.580 1968.730 34.640 ;
        RECT 1970.710 34.580 1971.030 34.640 ;
        RECT 1968.410 34.440 1971.030 34.580 ;
        RECT 1968.410 34.380 1968.730 34.440 ;
        RECT 1970.710 34.380 1971.030 34.440 ;
        RECT 1970.710 5.340 1971.030 5.400 ;
        RECT 1971.185 5.340 1971.475 5.385 ;
        RECT 1970.710 5.200 1971.475 5.340 ;
        RECT 1970.710 5.140 1971.030 5.200 ;
        RECT 1971.185 5.155 1971.475 5.200 ;
        RECT 1971.170 2.960 1971.490 3.020 ;
        RECT 1970.975 2.820 1971.490 2.960 ;
        RECT 1971.170 2.760 1971.490 2.820 ;
      LAYER via ;
        RECT 1960.620 1684.400 1960.880 1684.660 ;
        RECT 1967.980 1684.400 1968.240 1684.660 ;
        RECT 1967.980 1641.900 1968.240 1642.160 ;
        RECT 1968.440 1641.900 1968.700 1642.160 ;
        RECT 1967.980 1586.820 1968.240 1587.080 ;
        RECT 1967.980 1538.880 1968.240 1539.140 ;
        RECT 1967.980 1490.260 1968.240 1490.520 ;
        RECT 1967.980 1400.840 1968.240 1401.100 ;
        RECT 1967.980 1393.360 1968.240 1393.620 ;
        RECT 1967.980 1304.280 1968.240 1304.540 ;
        RECT 1967.980 1248.860 1968.240 1249.120 ;
        RECT 1968.900 1248.860 1969.160 1249.120 ;
        RECT 1966.600 1193.440 1966.860 1193.700 ;
        RECT 1967.520 1193.440 1967.780 1193.700 ;
        RECT 1966.600 1121.020 1966.860 1121.280 ;
        RECT 1967.520 1121.020 1967.780 1121.280 ;
        RECT 1967.520 1024.460 1967.780 1024.720 ;
        RECT 1967.520 965.300 1967.780 965.560 ;
        RECT 1967.520 958.840 1967.780 959.100 ;
        RECT 1967.520 917.360 1967.780 917.620 ;
        RECT 1966.600 910.560 1966.860 910.820 ;
        RECT 1967.520 910.560 1967.780 910.820 ;
        RECT 1968.440 814.000 1968.700 814.260 ;
        RECT 1967.980 766.060 1968.240 766.320 ;
        RECT 1967.980 742.260 1968.240 742.520 ;
        RECT 1968.440 710.640 1968.700 710.900 ;
        RECT 1967.980 655.220 1968.240 655.480 ;
        RECT 1968.900 655.220 1969.160 655.480 ;
        RECT 1967.980 600.140 1968.240 600.400 ;
        RECT 1967.980 552.200 1968.240 552.460 ;
        RECT 1967.980 524.320 1968.240 524.580 ;
        RECT 1968.440 523.640 1968.700 523.900 ;
        RECT 1968.440 503.240 1968.700 503.500 ;
        RECT 1967.980 434.220 1968.240 434.480 ;
        RECT 1968.440 372.340 1968.700 372.600 ;
        RECT 1968.900 324.400 1969.160 324.660 ;
        RECT 1967.520 276.120 1967.780 276.380 ;
        RECT 1968.900 276.120 1969.160 276.380 ;
        RECT 1967.060 227.840 1967.320 228.100 ;
        RECT 1968.440 227.840 1968.700 228.100 ;
        RECT 1967.980 186.020 1968.240 186.280 ;
        RECT 1968.440 138.080 1968.700 138.340 ;
        RECT 1968.440 90.140 1968.700 90.400 ;
        RECT 1968.440 89.460 1968.700 89.720 ;
        RECT 1968.440 34.380 1968.700 34.640 ;
        RECT 1970.740 34.380 1971.000 34.640 ;
        RECT 1970.740 5.140 1971.000 5.400 ;
        RECT 1971.200 2.760 1971.460 3.020 ;
      LAYER met2 ;
        RECT 1960.545 1700.000 1960.825 1704.000 ;
        RECT 1960.680 1684.690 1960.820 1700.000 ;
        RECT 1960.620 1684.370 1960.880 1684.690 ;
        RECT 1967.980 1684.370 1968.240 1684.690 ;
        RECT 1968.040 1642.190 1968.180 1684.370 ;
        RECT 1967.980 1641.870 1968.240 1642.190 ;
        RECT 1968.440 1641.870 1968.700 1642.190 ;
        RECT 1968.500 1594.330 1968.640 1641.870 ;
        RECT 1968.040 1594.190 1968.640 1594.330 ;
        RECT 1968.040 1587.110 1968.180 1594.190 ;
        RECT 1967.980 1586.790 1968.240 1587.110 ;
        RECT 1967.980 1538.850 1968.240 1539.170 ;
        RECT 1968.040 1490.550 1968.180 1538.850 ;
        RECT 1967.980 1490.230 1968.240 1490.550 ;
        RECT 1967.980 1400.810 1968.240 1401.130 ;
        RECT 1968.040 1393.650 1968.180 1400.810 ;
        RECT 1967.980 1393.330 1968.240 1393.650 ;
        RECT 1967.980 1304.250 1968.240 1304.570 ;
        RECT 1968.040 1297.285 1968.180 1304.250 ;
        RECT 1967.970 1296.915 1968.250 1297.285 ;
        RECT 1968.890 1296.915 1969.170 1297.285 ;
        RECT 1968.960 1249.150 1969.100 1296.915 ;
        RECT 1967.980 1248.830 1968.240 1249.150 ;
        RECT 1968.900 1248.830 1969.160 1249.150 ;
        RECT 1968.040 1200.610 1968.180 1248.830 ;
        RECT 1967.580 1200.470 1968.180 1200.610 ;
        RECT 1967.580 1193.730 1967.720 1200.470 ;
        RECT 1966.600 1193.410 1966.860 1193.730 ;
        RECT 1967.520 1193.410 1967.780 1193.730 ;
        RECT 1966.660 1145.645 1966.800 1193.410 ;
        RECT 1966.590 1145.275 1966.870 1145.645 ;
        RECT 1967.510 1145.275 1967.790 1145.645 ;
        RECT 1967.580 1121.310 1967.720 1145.275 ;
        RECT 1966.600 1120.990 1966.860 1121.310 ;
        RECT 1967.520 1120.990 1967.780 1121.310 ;
        RECT 1966.660 1097.365 1966.800 1120.990 ;
        RECT 1966.590 1096.995 1966.870 1097.365 ;
        RECT 1967.510 1096.995 1967.790 1097.365 ;
        RECT 1967.580 1024.750 1967.720 1096.995 ;
        RECT 1967.520 1024.430 1967.780 1024.750 ;
        RECT 1967.520 965.270 1967.780 965.590 ;
        RECT 1967.580 959.130 1967.720 965.270 ;
        RECT 1967.520 958.810 1967.780 959.130 ;
        RECT 1967.520 917.330 1967.780 917.650 ;
        RECT 1967.580 910.850 1967.720 917.330 ;
        RECT 1966.600 910.530 1966.860 910.850 ;
        RECT 1967.520 910.530 1967.780 910.850 ;
        RECT 1966.660 862.765 1966.800 910.530 ;
        RECT 1966.590 862.395 1966.870 862.765 ;
        RECT 1967.970 862.395 1968.250 862.765 ;
        RECT 1968.040 815.165 1968.180 862.395 ;
        RECT 1967.970 814.795 1968.250 815.165 ;
        RECT 1968.430 814.115 1968.710 814.485 ;
        RECT 1968.440 813.970 1968.700 814.115 ;
        RECT 1967.980 766.030 1968.240 766.350 ;
        RECT 1968.040 742.550 1968.180 766.030 ;
        RECT 1967.980 742.230 1968.240 742.550 ;
        RECT 1968.440 710.610 1968.700 710.930 ;
        RECT 1968.500 669.530 1968.640 710.610 ;
        RECT 1968.500 669.390 1969.100 669.530 ;
        RECT 1968.960 655.510 1969.100 669.390 ;
        RECT 1967.980 655.190 1968.240 655.510 ;
        RECT 1968.900 655.190 1969.160 655.510 ;
        RECT 1968.040 608.445 1968.180 655.190 ;
        RECT 1967.970 608.075 1968.250 608.445 ;
        RECT 1967.970 607.395 1968.250 607.765 ;
        RECT 1968.040 600.430 1968.180 607.395 ;
        RECT 1967.980 600.110 1968.240 600.430 ;
        RECT 1967.980 552.170 1968.240 552.490 ;
        RECT 1968.040 524.610 1968.180 552.170 ;
        RECT 1967.980 524.290 1968.240 524.610 ;
        RECT 1968.440 523.610 1968.700 523.930 ;
        RECT 1968.500 503.530 1968.640 523.610 ;
        RECT 1968.440 503.210 1968.700 503.530 ;
        RECT 1967.980 434.190 1968.240 434.510 ;
        RECT 1968.040 379.170 1968.180 434.190 ;
        RECT 1968.040 379.030 1968.640 379.170 ;
        RECT 1968.500 372.630 1968.640 379.030 ;
        RECT 1968.440 372.310 1968.700 372.630 ;
        RECT 1968.900 324.370 1969.160 324.690 ;
        RECT 1968.960 276.410 1969.100 324.370 ;
        RECT 1967.520 276.090 1967.780 276.410 ;
        RECT 1968.900 276.090 1969.160 276.410 ;
        RECT 1967.580 275.925 1967.720 276.090 ;
        RECT 1967.510 275.555 1967.790 275.925 ;
        RECT 1968.430 275.555 1968.710 275.925 ;
        RECT 1968.500 228.130 1968.640 275.555 ;
        RECT 1967.060 227.810 1967.320 228.130 ;
        RECT 1968.440 227.810 1968.700 228.130 ;
        RECT 1967.120 186.845 1967.260 227.810 ;
        RECT 1967.050 186.475 1967.330 186.845 ;
        RECT 1967.970 186.475 1968.250 186.845 ;
        RECT 1968.040 186.310 1968.180 186.475 ;
        RECT 1967.980 185.990 1968.240 186.310 ;
        RECT 1968.440 138.050 1968.700 138.370 ;
        RECT 1968.500 90.430 1968.640 138.050 ;
        RECT 1968.440 90.110 1968.700 90.430 ;
        RECT 1968.440 89.430 1968.700 89.750 ;
        RECT 1968.500 34.670 1968.640 89.430 ;
        RECT 1968.440 34.350 1968.700 34.670 ;
        RECT 1970.740 34.350 1971.000 34.670 ;
        RECT 1970.800 5.430 1970.940 34.350 ;
        RECT 1970.740 5.110 1971.000 5.430 ;
        RECT 1971.200 2.730 1971.460 3.050 ;
        RECT 1971.260 2.400 1971.400 2.730 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
      LAYER via2 ;
        RECT 1967.970 1296.960 1968.250 1297.240 ;
        RECT 1968.890 1296.960 1969.170 1297.240 ;
        RECT 1966.590 1145.320 1966.870 1145.600 ;
        RECT 1967.510 1145.320 1967.790 1145.600 ;
        RECT 1966.590 1097.040 1966.870 1097.320 ;
        RECT 1967.510 1097.040 1967.790 1097.320 ;
        RECT 1966.590 862.440 1966.870 862.720 ;
        RECT 1967.970 862.440 1968.250 862.720 ;
        RECT 1967.970 814.840 1968.250 815.120 ;
        RECT 1968.430 814.160 1968.710 814.440 ;
        RECT 1967.970 608.120 1968.250 608.400 ;
        RECT 1967.970 607.440 1968.250 607.720 ;
        RECT 1967.510 275.600 1967.790 275.880 ;
        RECT 1968.430 275.600 1968.710 275.880 ;
        RECT 1967.050 186.520 1967.330 186.800 ;
        RECT 1967.970 186.520 1968.250 186.800 ;
      LAYER met3 ;
        RECT 1967.945 1297.250 1968.275 1297.265 ;
        RECT 1968.865 1297.250 1969.195 1297.265 ;
        RECT 1967.945 1296.950 1969.195 1297.250 ;
        RECT 1967.945 1296.935 1968.275 1296.950 ;
        RECT 1968.865 1296.935 1969.195 1296.950 ;
        RECT 1966.565 1145.610 1966.895 1145.625 ;
        RECT 1967.485 1145.610 1967.815 1145.625 ;
        RECT 1966.565 1145.310 1967.815 1145.610 ;
        RECT 1966.565 1145.295 1966.895 1145.310 ;
        RECT 1967.485 1145.295 1967.815 1145.310 ;
        RECT 1966.565 1097.330 1966.895 1097.345 ;
        RECT 1967.485 1097.330 1967.815 1097.345 ;
        RECT 1966.565 1097.030 1967.815 1097.330 ;
        RECT 1966.565 1097.015 1966.895 1097.030 ;
        RECT 1967.485 1097.015 1967.815 1097.030 ;
        RECT 1966.565 862.730 1966.895 862.745 ;
        RECT 1967.945 862.730 1968.275 862.745 ;
        RECT 1966.565 862.430 1968.275 862.730 ;
        RECT 1966.565 862.415 1966.895 862.430 ;
        RECT 1967.945 862.415 1968.275 862.430 ;
        RECT 1967.945 815.130 1968.275 815.145 ;
        RECT 1967.945 814.815 1968.490 815.130 ;
        RECT 1968.190 814.465 1968.490 814.815 ;
        RECT 1968.190 814.150 1968.735 814.465 ;
        RECT 1968.405 814.135 1968.735 814.150 ;
        RECT 1967.945 608.095 1968.275 608.425 ;
        RECT 1967.960 607.745 1968.260 608.095 ;
        RECT 1967.945 607.415 1968.275 607.745 ;
        RECT 1967.485 275.890 1967.815 275.905 ;
        RECT 1968.405 275.890 1968.735 275.905 ;
        RECT 1967.485 275.590 1968.735 275.890 ;
        RECT 1967.485 275.575 1967.815 275.590 ;
        RECT 1968.405 275.575 1968.735 275.590 ;
        RECT 1967.025 186.810 1967.355 186.825 ;
        RECT 1967.945 186.810 1968.275 186.825 ;
        RECT 1967.025 186.510 1968.275 186.810 ;
        RECT 1967.025 186.495 1967.355 186.510 ;
        RECT 1967.945 186.495 1968.275 186.510 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1967.950 1685.280 1968.270 1685.340 ;
        RECT 1987.270 1685.280 1987.590 1685.340 ;
        RECT 1967.950 1685.140 1987.590 1685.280 ;
        RECT 1967.950 1685.080 1968.270 1685.140 ;
        RECT 1987.270 1685.080 1987.590 1685.140 ;
      LAYER via ;
        RECT 1967.980 1685.080 1968.240 1685.340 ;
        RECT 1987.300 1685.080 1987.560 1685.340 ;
      LAYER met2 ;
        RECT 1967.905 1700.000 1968.185 1704.000 ;
        RECT 1968.040 1685.370 1968.180 1700.000 ;
        RECT 1967.980 1685.050 1968.240 1685.370 ;
        RECT 1987.300 1685.050 1987.560 1685.370 ;
        RECT 1987.360 7.210 1987.500 1685.050 ;
        RECT 1987.360 7.070 1989.340 7.210 ;
        RECT 1989.200 2.400 1989.340 7.070 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1975.310 1683.920 1975.630 1683.980 ;
        RECT 1979.450 1683.920 1979.770 1683.980 ;
        RECT 1975.310 1683.780 1979.770 1683.920 ;
        RECT 1975.310 1683.720 1975.630 1683.780 ;
        RECT 1979.450 1683.720 1979.770 1683.780 ;
        RECT 1979.450 15.200 1979.770 15.260 ;
        RECT 2006.590 15.200 2006.910 15.260 ;
        RECT 1979.450 15.060 2006.910 15.200 ;
        RECT 1979.450 15.000 1979.770 15.060 ;
        RECT 2006.590 15.000 2006.910 15.060 ;
      LAYER via ;
        RECT 1975.340 1683.720 1975.600 1683.980 ;
        RECT 1979.480 1683.720 1979.740 1683.980 ;
        RECT 1979.480 15.000 1979.740 15.260 ;
        RECT 2006.620 15.000 2006.880 15.260 ;
      LAYER met2 ;
        RECT 1975.265 1700.000 1975.545 1704.000 ;
        RECT 1975.400 1684.010 1975.540 1700.000 ;
        RECT 1975.340 1683.690 1975.600 1684.010 ;
        RECT 1979.480 1683.690 1979.740 1684.010 ;
        RECT 1979.540 15.290 1979.680 1683.690 ;
        RECT 1979.480 14.970 1979.740 15.290 ;
        RECT 2006.620 14.970 2006.880 15.290 ;
        RECT 2006.680 2.400 2006.820 14.970 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1982.670 1683.920 1982.990 1683.980 ;
        RECT 1990.950 1683.920 1991.270 1683.980 ;
        RECT 1982.670 1683.780 1991.270 1683.920 ;
        RECT 1982.670 1683.720 1982.990 1683.780 ;
        RECT 1990.950 1683.720 1991.270 1683.780 ;
        RECT 1990.950 15.540 1991.270 15.600 ;
        RECT 1990.950 15.400 2007.280 15.540 ;
        RECT 1990.950 15.340 1991.270 15.400 ;
        RECT 2007.140 15.200 2007.280 15.400 ;
        RECT 2024.530 15.200 2024.850 15.260 ;
        RECT 2007.140 15.060 2024.850 15.200 ;
        RECT 2024.530 15.000 2024.850 15.060 ;
      LAYER via ;
        RECT 1982.700 1683.720 1982.960 1683.980 ;
        RECT 1990.980 1683.720 1991.240 1683.980 ;
        RECT 1990.980 15.340 1991.240 15.600 ;
        RECT 2024.560 15.000 2024.820 15.260 ;
      LAYER met2 ;
        RECT 1982.625 1700.000 1982.905 1704.000 ;
        RECT 1982.760 1684.010 1982.900 1700.000 ;
        RECT 1982.700 1683.690 1982.960 1684.010 ;
        RECT 1990.980 1683.690 1991.240 1684.010 ;
        RECT 1991.040 15.630 1991.180 1683.690 ;
        RECT 1990.980 15.310 1991.240 15.630 ;
        RECT 2024.560 14.970 2024.820 15.290 ;
        RECT 2024.620 2.400 2024.760 14.970 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1990.030 1689.020 1990.350 1689.080 ;
        RECT 1997.850 1689.020 1998.170 1689.080 ;
        RECT 1990.030 1688.880 1998.170 1689.020 ;
        RECT 1990.030 1688.820 1990.350 1688.880 ;
        RECT 1997.850 1688.820 1998.170 1688.880 ;
        RECT 1997.850 18.940 1998.170 19.000 ;
        RECT 2042.470 18.940 2042.790 19.000 ;
        RECT 1997.850 18.800 2042.790 18.940 ;
        RECT 1997.850 18.740 1998.170 18.800 ;
        RECT 2042.470 18.740 2042.790 18.800 ;
      LAYER via ;
        RECT 1990.060 1688.820 1990.320 1689.080 ;
        RECT 1997.880 1688.820 1998.140 1689.080 ;
        RECT 1997.880 18.740 1998.140 19.000 ;
        RECT 2042.500 18.740 2042.760 19.000 ;
      LAYER met2 ;
        RECT 1989.985 1700.000 1990.265 1704.000 ;
        RECT 1990.120 1689.110 1990.260 1700.000 ;
        RECT 1990.060 1688.790 1990.320 1689.110 ;
        RECT 1997.880 1688.790 1998.140 1689.110 ;
        RECT 1997.940 19.030 1998.080 1688.790 ;
        RECT 1997.880 18.710 1998.140 19.030 ;
        RECT 2042.500 18.710 2042.760 19.030 ;
        RECT 2042.560 2.400 2042.700 18.710 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1457.885 1482.485 1458.055 1518.015 ;
        RECT 1456.965 1373.345 1457.135 1462.595 ;
        RECT 1458.345 1021.445 1458.515 1097.095 ;
        RECT 1458.345 868.445 1458.515 910.775 ;
        RECT 1456.965 648.125 1457.135 649.655 ;
        RECT 1457.425 552.245 1457.595 600.355 ;
        RECT 1457.425 179.605 1457.595 234.515 ;
        RECT 1457.885 83.045 1458.055 131.155 ;
      LAYER mcon ;
        RECT 1457.885 1517.845 1458.055 1518.015 ;
        RECT 1456.965 1462.425 1457.135 1462.595 ;
        RECT 1458.345 1096.925 1458.515 1097.095 ;
        RECT 1458.345 910.605 1458.515 910.775 ;
        RECT 1456.965 649.485 1457.135 649.655 ;
        RECT 1457.425 600.185 1457.595 600.355 ;
        RECT 1457.425 234.345 1457.595 234.515 ;
        RECT 1457.885 130.985 1458.055 131.155 ;
      LAYER met1 ;
        RECT 1457.810 1587.020 1458.130 1587.080 ;
        RECT 1458.270 1587.020 1458.590 1587.080 ;
        RECT 1457.810 1586.880 1458.590 1587.020 ;
        RECT 1457.810 1586.820 1458.130 1586.880 ;
        RECT 1458.270 1586.820 1458.590 1586.880 ;
        RECT 1458.730 1524.800 1459.050 1524.860 ;
        RECT 1459.190 1524.800 1459.510 1524.860 ;
        RECT 1458.730 1524.660 1459.510 1524.800 ;
        RECT 1458.730 1524.600 1459.050 1524.660 ;
        RECT 1459.190 1524.600 1459.510 1524.660 ;
        RECT 1457.825 1518.000 1458.115 1518.045 ;
        RECT 1458.730 1518.000 1459.050 1518.060 ;
        RECT 1457.825 1517.860 1459.050 1518.000 ;
        RECT 1457.825 1517.815 1458.115 1517.860 ;
        RECT 1458.730 1517.800 1459.050 1517.860 ;
        RECT 1457.810 1482.640 1458.130 1482.700 ;
        RECT 1457.615 1482.500 1458.130 1482.640 ;
        RECT 1457.810 1482.440 1458.130 1482.500 ;
        RECT 1456.905 1462.580 1457.195 1462.625 ;
        RECT 1457.810 1462.580 1458.130 1462.640 ;
        RECT 1456.905 1462.440 1458.130 1462.580 ;
        RECT 1456.905 1462.395 1457.195 1462.440 ;
        RECT 1457.810 1462.380 1458.130 1462.440 ;
        RECT 1456.890 1373.500 1457.210 1373.560 ;
        RECT 1456.695 1373.360 1457.210 1373.500 ;
        RECT 1456.890 1373.300 1457.210 1373.360 ;
        RECT 1457.350 1290.200 1457.670 1290.260 ;
        RECT 1457.810 1290.200 1458.130 1290.260 ;
        RECT 1457.350 1290.060 1458.130 1290.200 ;
        RECT 1457.350 1290.000 1457.670 1290.060 ;
        RECT 1457.810 1290.000 1458.130 1290.060 ;
        RECT 1457.350 1207.580 1457.670 1207.640 ;
        RECT 1458.270 1207.580 1458.590 1207.640 ;
        RECT 1457.350 1207.440 1458.590 1207.580 ;
        RECT 1457.350 1207.380 1457.670 1207.440 ;
        RECT 1458.270 1207.380 1458.590 1207.440 ;
        RECT 1459.190 1104.900 1459.510 1104.960 ;
        RECT 1458.360 1104.760 1459.510 1104.900 ;
        RECT 1458.360 1104.280 1458.500 1104.760 ;
        RECT 1459.190 1104.700 1459.510 1104.760 ;
        RECT 1458.270 1104.020 1458.590 1104.280 ;
        RECT 1458.270 1097.080 1458.590 1097.140 ;
        RECT 1458.075 1096.940 1458.590 1097.080 ;
        RECT 1458.270 1096.880 1458.590 1096.940 ;
        RECT 1458.270 1021.600 1458.590 1021.660 ;
        RECT 1458.075 1021.460 1458.590 1021.600 ;
        RECT 1458.270 1021.400 1458.590 1021.460 ;
        RECT 1457.810 917.900 1458.130 917.960 ;
        RECT 1458.270 917.900 1458.590 917.960 ;
        RECT 1457.810 917.760 1458.590 917.900 ;
        RECT 1457.810 917.700 1458.130 917.760 ;
        RECT 1458.270 917.700 1458.590 917.760 ;
        RECT 1458.270 910.760 1458.590 910.820 ;
        RECT 1458.075 910.620 1458.590 910.760 ;
        RECT 1458.270 910.560 1458.590 910.620 ;
        RECT 1458.270 868.600 1458.590 868.660 ;
        RECT 1458.075 868.460 1458.590 868.600 ;
        RECT 1458.270 868.400 1458.590 868.460 ;
        RECT 1457.350 765.920 1457.670 765.980 ;
        RECT 1457.810 765.920 1458.130 765.980 ;
        RECT 1457.350 765.780 1458.130 765.920 ;
        RECT 1457.350 765.720 1457.670 765.780 ;
        RECT 1457.810 765.720 1458.130 765.780 ;
        RECT 1456.905 649.640 1457.195 649.685 ;
        RECT 1457.810 649.640 1458.130 649.700 ;
        RECT 1456.905 649.500 1458.130 649.640 ;
        RECT 1456.905 649.455 1457.195 649.500 ;
        RECT 1457.810 649.440 1458.130 649.500 ;
        RECT 1456.905 648.280 1457.195 648.325 ;
        RECT 1457.350 648.280 1457.670 648.340 ;
        RECT 1456.905 648.140 1457.670 648.280 ;
        RECT 1456.905 648.095 1457.195 648.140 ;
        RECT 1457.350 648.080 1457.670 648.140 ;
        RECT 1457.350 600.340 1457.670 600.400 ;
        RECT 1457.155 600.200 1457.670 600.340 ;
        RECT 1457.350 600.140 1457.670 600.200 ;
        RECT 1457.350 552.400 1457.670 552.460 ;
        RECT 1457.155 552.260 1457.670 552.400 ;
        RECT 1457.350 552.200 1457.670 552.260 ;
        RECT 1457.350 517.520 1457.670 517.780 ;
        RECT 1457.440 517.380 1457.580 517.520 ;
        RECT 1458.270 517.380 1458.590 517.440 ;
        RECT 1457.440 517.240 1458.590 517.380 ;
        RECT 1458.270 517.180 1458.590 517.240 ;
        RECT 1457.810 427.960 1458.130 428.020 ;
        RECT 1458.270 427.960 1458.590 428.020 ;
        RECT 1457.810 427.820 1458.590 427.960 ;
        RECT 1457.810 427.760 1458.130 427.820 ;
        RECT 1458.270 427.760 1458.590 427.820 ;
        RECT 1456.890 372.880 1457.210 372.940 ;
        RECT 1457.810 372.880 1458.130 372.940 ;
        RECT 1456.890 372.740 1458.130 372.880 ;
        RECT 1456.890 372.680 1457.210 372.740 ;
        RECT 1457.810 372.680 1458.130 372.740 ;
        RECT 1456.890 338.200 1457.210 338.260 ;
        RECT 1457.350 338.200 1457.670 338.260 ;
        RECT 1456.890 338.060 1457.670 338.200 ;
        RECT 1456.890 338.000 1457.210 338.060 ;
        RECT 1457.350 338.000 1457.670 338.060 ;
        RECT 1457.350 290.260 1457.670 290.320 ;
        RECT 1456.980 290.120 1457.670 290.260 ;
        RECT 1456.980 289.640 1457.120 290.120 ;
        RECT 1457.350 290.060 1457.670 290.120 ;
        RECT 1456.890 289.380 1457.210 289.640 ;
        RECT 1456.890 241.640 1457.210 241.700 ;
        RECT 1457.350 241.640 1457.670 241.700 ;
        RECT 1456.890 241.500 1457.670 241.640 ;
        RECT 1456.890 241.440 1457.210 241.500 ;
        RECT 1457.350 241.440 1457.670 241.500 ;
        RECT 1457.350 234.500 1457.670 234.560 ;
        RECT 1457.155 234.360 1457.670 234.500 ;
        RECT 1457.350 234.300 1457.670 234.360 ;
        RECT 1457.365 179.760 1457.655 179.805 ;
        RECT 1457.810 179.760 1458.130 179.820 ;
        RECT 1457.365 179.620 1458.130 179.760 ;
        RECT 1457.365 179.575 1457.655 179.620 ;
        RECT 1457.810 179.560 1458.130 179.620 ;
        RECT 1457.810 138.280 1458.130 138.340 ;
        RECT 1458.270 138.280 1458.590 138.340 ;
        RECT 1457.810 138.140 1458.590 138.280 ;
        RECT 1457.810 138.080 1458.130 138.140 ;
        RECT 1458.270 138.080 1458.590 138.140 ;
        RECT 1457.825 131.140 1458.115 131.185 ;
        RECT 1458.270 131.140 1458.590 131.200 ;
        RECT 1457.825 131.000 1458.590 131.140 ;
        RECT 1457.825 130.955 1458.115 131.000 ;
        RECT 1458.270 130.940 1458.590 131.000 ;
        RECT 1457.810 83.200 1458.130 83.260 ;
        RECT 1457.615 83.060 1458.130 83.200 ;
        RECT 1457.810 83.000 1458.130 83.060 ;
        RECT 758.610 60.760 758.930 60.820 ;
        RECT 1457.810 60.760 1458.130 60.820 ;
        RECT 758.610 60.620 1458.130 60.760 ;
        RECT 758.610 60.560 758.930 60.620 ;
        RECT 1457.810 60.560 1458.130 60.620 ;
      LAYER via ;
        RECT 1457.840 1586.820 1458.100 1587.080 ;
        RECT 1458.300 1586.820 1458.560 1587.080 ;
        RECT 1458.760 1524.600 1459.020 1524.860 ;
        RECT 1459.220 1524.600 1459.480 1524.860 ;
        RECT 1458.760 1517.800 1459.020 1518.060 ;
        RECT 1457.840 1482.440 1458.100 1482.700 ;
        RECT 1457.840 1462.380 1458.100 1462.640 ;
        RECT 1456.920 1373.300 1457.180 1373.560 ;
        RECT 1457.380 1290.000 1457.640 1290.260 ;
        RECT 1457.840 1290.000 1458.100 1290.260 ;
        RECT 1457.380 1207.380 1457.640 1207.640 ;
        RECT 1458.300 1207.380 1458.560 1207.640 ;
        RECT 1459.220 1104.700 1459.480 1104.960 ;
        RECT 1458.300 1104.020 1458.560 1104.280 ;
        RECT 1458.300 1096.880 1458.560 1097.140 ;
        RECT 1458.300 1021.400 1458.560 1021.660 ;
        RECT 1457.840 917.700 1458.100 917.960 ;
        RECT 1458.300 917.700 1458.560 917.960 ;
        RECT 1458.300 910.560 1458.560 910.820 ;
        RECT 1458.300 868.400 1458.560 868.660 ;
        RECT 1457.380 765.720 1457.640 765.980 ;
        RECT 1457.840 765.720 1458.100 765.980 ;
        RECT 1457.840 649.440 1458.100 649.700 ;
        RECT 1457.380 648.080 1457.640 648.340 ;
        RECT 1457.380 600.140 1457.640 600.400 ;
        RECT 1457.380 552.200 1457.640 552.460 ;
        RECT 1457.380 517.520 1457.640 517.780 ;
        RECT 1458.300 517.180 1458.560 517.440 ;
        RECT 1457.840 427.760 1458.100 428.020 ;
        RECT 1458.300 427.760 1458.560 428.020 ;
        RECT 1456.920 372.680 1457.180 372.940 ;
        RECT 1457.840 372.680 1458.100 372.940 ;
        RECT 1456.920 338.000 1457.180 338.260 ;
        RECT 1457.380 338.000 1457.640 338.260 ;
        RECT 1457.380 290.060 1457.640 290.320 ;
        RECT 1456.920 289.380 1457.180 289.640 ;
        RECT 1456.920 241.440 1457.180 241.700 ;
        RECT 1457.380 241.440 1457.640 241.700 ;
        RECT 1457.380 234.300 1457.640 234.560 ;
        RECT 1457.840 179.560 1458.100 179.820 ;
        RECT 1457.840 138.080 1458.100 138.340 ;
        RECT 1458.300 138.080 1458.560 138.340 ;
        RECT 1458.300 130.940 1458.560 131.200 ;
        RECT 1457.840 83.000 1458.100 83.260 ;
        RECT 758.640 60.560 758.900 60.820 ;
        RECT 1457.840 60.560 1458.100 60.820 ;
      LAYER met2 ;
        RECT 1460.985 1701.090 1461.265 1704.000 ;
        RECT 1458.820 1700.950 1461.265 1701.090 ;
        RECT 1458.820 1677.970 1458.960 1700.950 ;
        RECT 1460.985 1700.000 1461.265 1700.950 ;
        RECT 1457.900 1677.830 1458.960 1677.970 ;
        RECT 1457.900 1597.050 1458.040 1677.830 ;
        RECT 1457.440 1596.910 1458.040 1597.050 ;
        RECT 1457.440 1595.690 1457.580 1596.910 ;
        RECT 1457.440 1595.550 1458.040 1595.690 ;
        RECT 1457.900 1587.110 1458.040 1595.550 ;
        RECT 1457.840 1586.790 1458.100 1587.110 ;
        RECT 1458.300 1586.790 1458.560 1587.110 ;
        RECT 1458.360 1531.885 1458.500 1586.790 ;
        RECT 1458.290 1531.515 1458.570 1531.885 ;
        RECT 1459.210 1531.515 1459.490 1531.885 ;
        RECT 1459.280 1524.890 1459.420 1531.515 ;
        RECT 1458.760 1524.570 1459.020 1524.890 ;
        RECT 1459.220 1524.570 1459.480 1524.890 ;
        RECT 1458.820 1518.090 1458.960 1524.570 ;
        RECT 1458.760 1517.770 1459.020 1518.090 ;
        RECT 1457.840 1482.410 1458.100 1482.730 ;
        RECT 1457.900 1462.670 1458.040 1482.410 ;
        RECT 1457.840 1462.350 1458.100 1462.670 ;
        RECT 1456.920 1373.270 1457.180 1373.590 ;
        RECT 1456.980 1290.485 1457.120 1373.270 ;
        RECT 1456.910 1290.115 1457.190 1290.485 ;
        RECT 1457.380 1289.970 1457.640 1290.290 ;
        RECT 1457.830 1290.115 1458.110 1290.485 ;
        RECT 1457.840 1289.970 1458.100 1290.115 ;
        RECT 1457.440 1207.670 1457.580 1289.970 ;
        RECT 1457.380 1207.350 1457.640 1207.670 ;
        RECT 1458.300 1207.350 1458.560 1207.670 ;
        RECT 1458.360 1176.810 1458.500 1207.350 ;
        RECT 1458.360 1176.670 1459.420 1176.810 ;
        RECT 1459.280 1104.990 1459.420 1176.670 ;
        RECT 1459.220 1104.670 1459.480 1104.990 ;
        RECT 1458.300 1103.990 1458.560 1104.310 ;
        RECT 1458.360 1097.170 1458.500 1103.990 ;
        RECT 1458.300 1096.850 1458.560 1097.170 ;
        RECT 1458.300 1021.370 1458.560 1021.690 ;
        RECT 1458.360 966.010 1458.500 1021.370 ;
        RECT 1457.900 965.870 1458.500 966.010 ;
        RECT 1457.900 917.990 1458.040 965.870 ;
        RECT 1457.840 917.670 1458.100 917.990 ;
        RECT 1458.300 917.670 1458.560 917.990 ;
        RECT 1458.360 910.850 1458.500 917.670 ;
        RECT 1458.300 910.530 1458.560 910.850 ;
        RECT 1458.300 868.370 1458.560 868.690 ;
        RECT 1458.360 821.285 1458.500 868.370 ;
        RECT 1457.370 820.915 1457.650 821.285 ;
        RECT 1458.290 820.915 1458.570 821.285 ;
        RECT 1457.440 766.010 1457.580 820.915 ;
        RECT 1457.380 765.690 1457.640 766.010 ;
        RECT 1457.840 765.690 1458.100 766.010 ;
        RECT 1457.900 649.730 1458.040 765.690 ;
        RECT 1457.840 649.410 1458.100 649.730 ;
        RECT 1457.380 648.050 1457.640 648.370 ;
        RECT 1457.440 600.430 1457.580 648.050 ;
        RECT 1457.380 600.110 1457.640 600.430 ;
        RECT 1457.380 552.170 1457.640 552.490 ;
        RECT 1457.440 517.810 1457.580 552.170 ;
        RECT 1457.380 517.490 1457.640 517.810 ;
        RECT 1458.300 517.150 1458.560 517.470 ;
        RECT 1458.360 428.050 1458.500 517.150 ;
        RECT 1457.840 427.730 1458.100 428.050 ;
        RECT 1458.300 427.730 1458.560 428.050 ;
        RECT 1457.900 372.970 1458.040 427.730 ;
        RECT 1456.920 372.650 1457.180 372.970 ;
        RECT 1457.840 372.650 1458.100 372.970 ;
        RECT 1456.980 338.290 1457.120 372.650 ;
        RECT 1456.920 337.970 1457.180 338.290 ;
        RECT 1457.380 337.970 1457.640 338.290 ;
        RECT 1457.440 290.350 1457.580 337.970 ;
        RECT 1457.380 290.030 1457.640 290.350 ;
        RECT 1456.920 289.350 1457.180 289.670 ;
        RECT 1456.980 241.730 1457.120 289.350 ;
        RECT 1456.920 241.410 1457.180 241.730 ;
        RECT 1457.380 241.410 1457.640 241.730 ;
        RECT 1457.440 234.590 1457.580 241.410 ;
        RECT 1457.380 234.270 1457.640 234.590 ;
        RECT 1457.840 179.530 1458.100 179.850 ;
        RECT 1457.900 138.370 1458.040 179.530 ;
        RECT 1457.840 138.050 1458.100 138.370 ;
        RECT 1458.300 138.050 1458.560 138.370 ;
        RECT 1458.360 131.230 1458.500 138.050 ;
        RECT 1458.300 130.910 1458.560 131.230 ;
        RECT 1457.840 82.970 1458.100 83.290 ;
        RECT 1457.900 60.850 1458.040 82.970 ;
        RECT 758.640 60.530 758.900 60.850 ;
        RECT 1457.840 60.530 1458.100 60.850 ;
        RECT 758.700 17.410 758.840 60.530 ;
        RECT 757.780 17.270 758.840 17.410 ;
        RECT 757.780 2.400 757.920 17.270 ;
        RECT 757.570 -4.800 758.130 2.400 ;
      LAYER via2 ;
        RECT 1458.290 1531.560 1458.570 1531.840 ;
        RECT 1459.210 1531.560 1459.490 1531.840 ;
        RECT 1456.910 1290.160 1457.190 1290.440 ;
        RECT 1457.830 1290.160 1458.110 1290.440 ;
        RECT 1457.370 820.960 1457.650 821.240 ;
        RECT 1458.290 820.960 1458.570 821.240 ;
      LAYER met3 ;
        RECT 1458.265 1531.850 1458.595 1531.865 ;
        RECT 1459.185 1531.850 1459.515 1531.865 ;
        RECT 1458.265 1531.550 1459.515 1531.850 ;
        RECT 1458.265 1531.535 1458.595 1531.550 ;
        RECT 1459.185 1531.535 1459.515 1531.550 ;
        RECT 1456.885 1290.450 1457.215 1290.465 ;
        RECT 1457.805 1290.450 1458.135 1290.465 ;
        RECT 1456.885 1290.150 1458.135 1290.450 ;
        RECT 1456.885 1290.135 1457.215 1290.150 ;
        RECT 1457.805 1290.135 1458.135 1290.150 ;
        RECT 1457.345 821.250 1457.675 821.265 ;
        RECT 1458.265 821.250 1458.595 821.265 ;
        RECT 1457.345 820.950 1458.595 821.250 ;
        RECT 1457.345 820.935 1457.675 820.950 ;
        RECT 1458.265 820.935 1458.595 820.950 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1997.390 1690.040 1997.710 1690.100 ;
        RECT 2000.610 1690.040 2000.930 1690.100 ;
        RECT 1997.390 1689.900 2000.930 1690.040 ;
        RECT 1997.390 1689.840 1997.710 1689.900 ;
        RECT 2000.610 1689.840 2000.930 1689.900 ;
        RECT 2000.610 18.260 2000.930 18.320 ;
        RECT 2060.410 18.260 2060.730 18.320 ;
        RECT 2000.610 18.120 2060.730 18.260 ;
        RECT 2000.610 18.060 2000.930 18.120 ;
        RECT 2060.410 18.060 2060.730 18.120 ;
      LAYER via ;
        RECT 1997.420 1689.840 1997.680 1690.100 ;
        RECT 2000.640 1689.840 2000.900 1690.100 ;
        RECT 2000.640 18.060 2000.900 18.320 ;
        RECT 2060.440 18.060 2060.700 18.320 ;
      LAYER met2 ;
        RECT 1997.345 1700.000 1997.625 1704.000 ;
        RECT 1997.480 1690.130 1997.620 1700.000 ;
        RECT 1997.420 1689.810 1997.680 1690.130 ;
        RECT 2000.640 1689.810 2000.900 1690.130 ;
        RECT 2000.700 18.350 2000.840 1689.810 ;
        RECT 2000.640 18.030 2000.900 18.350 ;
        RECT 2060.440 18.030 2060.700 18.350 ;
        RECT 2060.500 2.400 2060.640 18.030 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2004.750 1686.980 2005.070 1687.040 ;
        RECT 2011.190 1686.980 2011.510 1687.040 ;
        RECT 2004.750 1686.840 2011.510 1686.980 ;
        RECT 2004.750 1686.780 2005.070 1686.840 ;
        RECT 2011.190 1686.780 2011.510 1686.840 ;
        RECT 2011.190 17.580 2011.510 17.640 ;
        RECT 2078.350 17.580 2078.670 17.640 ;
        RECT 2011.190 17.440 2078.670 17.580 ;
        RECT 2011.190 17.380 2011.510 17.440 ;
        RECT 2078.350 17.380 2078.670 17.440 ;
      LAYER via ;
        RECT 2004.780 1686.780 2005.040 1687.040 ;
        RECT 2011.220 1686.780 2011.480 1687.040 ;
        RECT 2011.220 17.380 2011.480 17.640 ;
        RECT 2078.380 17.380 2078.640 17.640 ;
      LAYER met2 ;
        RECT 2004.705 1700.000 2004.985 1704.000 ;
        RECT 2004.840 1687.070 2004.980 1700.000 ;
        RECT 2004.780 1686.750 2005.040 1687.070 ;
        RECT 2011.220 1686.750 2011.480 1687.070 ;
        RECT 2011.280 17.670 2011.420 1686.750 ;
        RECT 2011.220 17.350 2011.480 17.670 ;
        RECT 2078.380 17.350 2078.640 17.670 ;
        RECT 2078.440 2.400 2078.580 17.350 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2013.950 18.600 2014.270 18.660 ;
        RECT 2095.830 18.600 2096.150 18.660 ;
        RECT 2013.950 18.460 2096.150 18.600 ;
        RECT 2013.950 18.400 2014.270 18.460 ;
        RECT 2095.830 18.400 2096.150 18.460 ;
      LAYER via ;
        RECT 2013.980 18.400 2014.240 18.660 ;
        RECT 2095.860 18.400 2096.120 18.660 ;
      LAYER met2 ;
        RECT 2012.065 1700.410 2012.345 1704.000 ;
        RECT 2012.065 1700.270 2014.180 1700.410 ;
        RECT 2012.065 1700.000 2012.345 1700.270 ;
        RECT 2014.040 18.690 2014.180 1700.270 ;
        RECT 2013.980 18.370 2014.240 18.690 ;
        RECT 2095.860 18.370 2096.120 18.690 ;
        RECT 2095.920 2.400 2096.060 18.370 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2021.310 17.240 2021.630 17.300 ;
        RECT 2113.770 17.240 2114.090 17.300 ;
        RECT 2021.310 17.100 2114.090 17.240 ;
        RECT 2021.310 17.040 2021.630 17.100 ;
        RECT 2113.770 17.040 2114.090 17.100 ;
      LAYER via ;
        RECT 2021.340 17.040 2021.600 17.300 ;
        RECT 2113.800 17.040 2114.060 17.300 ;
      LAYER met2 ;
        RECT 2019.425 1700.410 2019.705 1704.000 ;
        RECT 2019.425 1700.270 2021.540 1700.410 ;
        RECT 2019.425 1700.000 2019.705 1700.270 ;
        RECT 2021.400 17.330 2021.540 1700.270 ;
        RECT 2021.340 17.010 2021.600 17.330 ;
        RECT 2113.800 17.010 2114.060 17.330 ;
        RECT 2113.860 2.400 2114.000 17.010 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2028.210 15.880 2028.530 15.940 ;
        RECT 2131.710 15.880 2132.030 15.940 ;
        RECT 2028.210 15.740 2132.030 15.880 ;
        RECT 2028.210 15.680 2028.530 15.740 ;
        RECT 2131.710 15.680 2132.030 15.740 ;
      LAYER via ;
        RECT 2028.240 15.680 2028.500 15.940 ;
        RECT 2131.740 15.680 2132.000 15.940 ;
      LAYER met2 ;
        RECT 2026.785 1700.410 2027.065 1704.000 ;
        RECT 2026.785 1700.270 2028.440 1700.410 ;
        RECT 2026.785 1700.000 2027.065 1700.270 ;
        RECT 2028.300 15.970 2028.440 1700.270 ;
        RECT 2028.240 15.650 2028.500 15.970 ;
        RECT 2131.740 15.650 2132.000 15.970 ;
        RECT 2131.800 2.400 2131.940 15.650 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2135.005 16.065 2136.095 16.235 ;
      LAYER mcon ;
        RECT 2135.925 16.065 2136.095 16.235 ;
      LAYER met1 ;
        RECT 2035.110 16.220 2035.430 16.280 ;
        RECT 2134.945 16.220 2135.235 16.265 ;
        RECT 2035.110 16.080 2135.235 16.220 ;
        RECT 2035.110 16.020 2035.430 16.080 ;
        RECT 2134.945 16.035 2135.235 16.080 ;
        RECT 2135.865 16.220 2136.155 16.265 ;
        RECT 2149.650 16.220 2149.970 16.280 ;
        RECT 2135.865 16.080 2149.970 16.220 ;
        RECT 2135.865 16.035 2136.155 16.080 ;
        RECT 2149.650 16.020 2149.970 16.080 ;
      LAYER via ;
        RECT 2035.140 16.020 2035.400 16.280 ;
        RECT 2149.680 16.020 2149.940 16.280 ;
      LAYER met2 ;
        RECT 2034.145 1700.410 2034.425 1704.000 ;
        RECT 2034.145 1700.270 2035.340 1700.410 ;
        RECT 2034.145 1700.000 2034.425 1700.270 ;
        RECT 2035.200 16.310 2035.340 1700.270 ;
        RECT 2035.140 15.990 2035.400 16.310 ;
        RECT 2149.680 15.990 2149.940 16.310 ;
        RECT 2149.740 2.400 2149.880 15.990 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2042.010 27.100 2042.330 27.160 ;
        RECT 2167.590 27.100 2167.910 27.160 ;
        RECT 2042.010 26.960 2167.910 27.100 ;
        RECT 2042.010 26.900 2042.330 26.960 ;
        RECT 2167.590 26.900 2167.910 26.960 ;
      LAYER via ;
        RECT 2042.040 26.900 2042.300 27.160 ;
        RECT 2167.620 26.900 2167.880 27.160 ;
      LAYER met2 ;
        RECT 2041.505 1700.410 2041.785 1704.000 ;
        RECT 2041.505 1700.270 2042.240 1700.410 ;
        RECT 2041.505 1700.000 2041.785 1700.270 ;
        RECT 2042.100 27.190 2042.240 1700.270 ;
        RECT 2042.040 26.870 2042.300 27.190 ;
        RECT 2167.620 26.870 2167.880 27.190 ;
        RECT 2167.680 2.400 2167.820 26.870 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2048.450 20.640 2048.770 20.700 ;
        RECT 2185.070 20.640 2185.390 20.700 ;
        RECT 2048.450 20.500 2185.390 20.640 ;
        RECT 2048.450 20.440 2048.770 20.500 ;
        RECT 2185.070 20.440 2185.390 20.500 ;
      LAYER via ;
        RECT 2048.480 20.440 2048.740 20.700 ;
        RECT 2185.100 20.440 2185.360 20.700 ;
      LAYER met2 ;
        RECT 2048.865 1700.410 2049.145 1704.000 ;
        RECT 2048.540 1700.270 2049.145 1700.410 ;
        RECT 2048.540 20.730 2048.680 1700.270 ;
        RECT 2048.865 1700.000 2049.145 1700.270 ;
        RECT 2048.480 20.410 2048.740 20.730 ;
        RECT 2185.100 20.410 2185.360 20.730 ;
        RECT 2185.160 2.400 2185.300 20.410 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2056.270 1690.380 2056.590 1690.440 ;
        RECT 2062.250 1690.380 2062.570 1690.440 ;
        RECT 2056.270 1690.240 2062.570 1690.380 ;
        RECT 2056.270 1690.180 2056.590 1690.240 ;
        RECT 2062.250 1690.180 2062.570 1690.240 ;
        RECT 2062.250 26.760 2062.570 26.820 ;
        RECT 2203.010 26.760 2203.330 26.820 ;
        RECT 2062.250 26.620 2203.330 26.760 ;
        RECT 2062.250 26.560 2062.570 26.620 ;
        RECT 2203.010 26.560 2203.330 26.620 ;
      LAYER via ;
        RECT 2056.300 1690.180 2056.560 1690.440 ;
        RECT 2062.280 1690.180 2062.540 1690.440 ;
        RECT 2062.280 26.560 2062.540 26.820 ;
        RECT 2203.040 26.560 2203.300 26.820 ;
      LAYER met2 ;
        RECT 2056.225 1700.000 2056.505 1704.000 ;
        RECT 2056.360 1690.470 2056.500 1700.000 ;
        RECT 2056.300 1690.150 2056.560 1690.470 ;
        RECT 2062.280 1690.150 2062.540 1690.470 ;
        RECT 2062.340 26.850 2062.480 1690.150 ;
        RECT 2062.280 26.530 2062.540 26.850 ;
        RECT 2203.040 26.530 2203.300 26.850 ;
        RECT 2203.100 2.400 2203.240 26.530 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2063.630 1686.640 2063.950 1686.700 ;
        RECT 2069.150 1686.640 2069.470 1686.700 ;
        RECT 2063.630 1686.500 2069.470 1686.640 ;
        RECT 2063.630 1686.440 2063.950 1686.500 ;
        RECT 2069.150 1686.440 2069.470 1686.500 ;
        RECT 2069.150 26.420 2069.470 26.480 ;
        RECT 2220.950 26.420 2221.270 26.480 ;
        RECT 2069.150 26.280 2221.270 26.420 ;
        RECT 2069.150 26.220 2069.470 26.280 ;
        RECT 2220.950 26.220 2221.270 26.280 ;
      LAYER via ;
        RECT 2063.660 1686.440 2063.920 1686.700 ;
        RECT 2069.180 1686.440 2069.440 1686.700 ;
        RECT 2069.180 26.220 2069.440 26.480 ;
        RECT 2220.980 26.220 2221.240 26.480 ;
      LAYER met2 ;
        RECT 2063.585 1700.000 2063.865 1704.000 ;
        RECT 2063.720 1686.730 2063.860 1700.000 ;
        RECT 2063.660 1686.410 2063.920 1686.730 ;
        RECT 2069.180 1686.410 2069.440 1686.730 ;
        RECT 2069.240 26.510 2069.380 1686.410 ;
        RECT 2069.180 26.190 2069.440 26.510 ;
        RECT 2220.980 26.190 2221.240 26.510 ;
        RECT 2221.040 2.400 2221.180 26.190 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1463.790 1678.140 1464.110 1678.200 ;
        RECT 1466.550 1678.140 1466.870 1678.200 ;
        RECT 1463.790 1678.000 1466.870 1678.140 ;
        RECT 1463.790 1677.940 1464.110 1678.000 ;
        RECT 1466.550 1677.940 1466.870 1678.000 ;
        RECT 779.310 66.200 779.630 66.260 ;
        RECT 1463.790 66.200 1464.110 66.260 ;
        RECT 779.310 66.060 1464.110 66.200 ;
        RECT 779.310 66.000 779.630 66.060 ;
        RECT 1463.790 66.000 1464.110 66.060 ;
      LAYER via ;
        RECT 1463.820 1677.940 1464.080 1678.200 ;
        RECT 1466.580 1677.940 1466.840 1678.200 ;
        RECT 779.340 66.000 779.600 66.260 ;
        RECT 1463.820 66.000 1464.080 66.260 ;
      LAYER met2 ;
        RECT 1468.345 1700.410 1468.625 1704.000 ;
        RECT 1466.640 1700.270 1468.625 1700.410 ;
        RECT 1466.640 1678.230 1466.780 1700.270 ;
        RECT 1468.345 1700.000 1468.625 1700.270 ;
        RECT 1463.820 1677.910 1464.080 1678.230 ;
        RECT 1466.580 1677.910 1466.840 1678.230 ;
        RECT 1463.880 66.290 1464.020 1677.910 ;
        RECT 779.340 65.970 779.600 66.290 ;
        RECT 1463.820 65.970 1464.080 66.290 ;
        RECT 779.400 17.410 779.540 65.970 ;
        RECT 775.720 17.270 779.540 17.410 ;
        RECT 775.720 2.400 775.860 17.270 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2070.990 1686.300 2071.310 1686.360 ;
        RECT 2076.510 1686.300 2076.830 1686.360 ;
        RECT 2070.990 1686.160 2076.830 1686.300 ;
        RECT 2070.990 1686.100 2071.310 1686.160 ;
        RECT 2076.510 1686.100 2076.830 1686.160 ;
        RECT 2076.510 26.080 2076.830 26.140 ;
        RECT 2238.890 26.080 2239.210 26.140 ;
        RECT 2076.510 25.940 2239.210 26.080 ;
        RECT 2076.510 25.880 2076.830 25.940 ;
        RECT 2238.890 25.880 2239.210 25.940 ;
      LAYER via ;
        RECT 2071.020 1686.100 2071.280 1686.360 ;
        RECT 2076.540 1686.100 2076.800 1686.360 ;
        RECT 2076.540 25.880 2076.800 26.140 ;
        RECT 2238.920 25.880 2239.180 26.140 ;
      LAYER met2 ;
        RECT 2070.945 1700.000 2071.225 1704.000 ;
        RECT 2071.080 1686.390 2071.220 1700.000 ;
        RECT 2071.020 1686.070 2071.280 1686.390 ;
        RECT 2076.540 1686.070 2076.800 1686.390 ;
        RECT 2076.600 26.170 2076.740 1686.070 ;
        RECT 2076.540 25.850 2076.800 26.170 ;
        RECT 2238.920 25.850 2239.180 26.170 ;
        RECT 2238.980 2.400 2239.120 25.850 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2077.890 1688.000 2078.210 1688.060 ;
        RECT 2082.950 1688.000 2083.270 1688.060 ;
        RECT 2077.890 1687.860 2083.270 1688.000 ;
        RECT 2077.890 1687.800 2078.210 1687.860 ;
        RECT 2082.950 1687.800 2083.270 1687.860 ;
        RECT 2082.950 25.740 2083.270 25.800 ;
        RECT 2256.370 25.740 2256.690 25.800 ;
        RECT 2082.950 25.600 2256.690 25.740 ;
        RECT 2082.950 25.540 2083.270 25.600 ;
        RECT 2256.370 25.540 2256.690 25.600 ;
      LAYER via ;
        RECT 2077.920 1687.800 2078.180 1688.060 ;
        RECT 2082.980 1687.800 2083.240 1688.060 ;
        RECT 2082.980 25.540 2083.240 25.800 ;
        RECT 2256.400 25.540 2256.660 25.800 ;
      LAYER met2 ;
        RECT 2077.845 1700.000 2078.125 1704.000 ;
        RECT 2077.980 1688.090 2078.120 1700.000 ;
        RECT 2077.920 1687.770 2078.180 1688.090 ;
        RECT 2082.980 1687.770 2083.240 1688.090 ;
        RECT 2083.040 25.830 2083.180 1687.770 ;
        RECT 2082.980 25.510 2083.240 25.830 ;
        RECT 2256.400 25.510 2256.660 25.830 ;
        RECT 2256.460 2.400 2256.600 25.510 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2085.250 1685.620 2085.570 1685.680 ;
        RECT 2089.850 1685.620 2090.170 1685.680 ;
        RECT 2085.250 1685.480 2090.170 1685.620 ;
        RECT 2085.250 1685.420 2085.570 1685.480 ;
        RECT 2089.850 1685.420 2090.170 1685.480 ;
        RECT 2089.850 25.400 2090.170 25.460 ;
        RECT 2274.310 25.400 2274.630 25.460 ;
        RECT 2089.850 25.260 2274.630 25.400 ;
        RECT 2089.850 25.200 2090.170 25.260 ;
        RECT 2274.310 25.200 2274.630 25.260 ;
      LAYER via ;
        RECT 2085.280 1685.420 2085.540 1685.680 ;
        RECT 2089.880 1685.420 2090.140 1685.680 ;
        RECT 2089.880 25.200 2090.140 25.460 ;
        RECT 2274.340 25.200 2274.600 25.460 ;
      LAYER met2 ;
        RECT 2085.205 1700.000 2085.485 1704.000 ;
        RECT 2085.340 1685.710 2085.480 1700.000 ;
        RECT 2085.280 1685.390 2085.540 1685.710 ;
        RECT 2089.880 1685.390 2090.140 1685.710 ;
        RECT 2089.940 25.490 2090.080 1685.390 ;
        RECT 2089.880 25.170 2090.140 25.490 ;
        RECT 2274.340 25.170 2274.600 25.490 ;
        RECT 2274.400 2.400 2274.540 25.170 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2092.610 1686.640 2092.930 1686.700 ;
        RECT 2097.210 1686.640 2097.530 1686.700 ;
        RECT 2092.610 1686.500 2097.530 1686.640 ;
        RECT 2092.610 1686.440 2092.930 1686.500 ;
        RECT 2097.210 1686.440 2097.530 1686.500 ;
        RECT 2097.210 25.060 2097.530 25.120 ;
        RECT 2292.250 25.060 2292.570 25.120 ;
        RECT 2097.210 24.920 2292.570 25.060 ;
        RECT 2097.210 24.860 2097.530 24.920 ;
        RECT 2292.250 24.860 2292.570 24.920 ;
      LAYER via ;
        RECT 2092.640 1686.440 2092.900 1686.700 ;
        RECT 2097.240 1686.440 2097.500 1686.700 ;
        RECT 2097.240 24.860 2097.500 25.120 ;
        RECT 2292.280 24.860 2292.540 25.120 ;
      LAYER met2 ;
        RECT 2092.565 1700.000 2092.845 1704.000 ;
        RECT 2092.700 1686.730 2092.840 1700.000 ;
        RECT 2092.640 1686.410 2092.900 1686.730 ;
        RECT 2097.240 1686.410 2097.500 1686.730 ;
        RECT 2097.300 25.150 2097.440 1686.410 ;
        RECT 2097.240 24.830 2097.500 25.150 ;
        RECT 2292.280 24.830 2292.540 25.150 ;
        RECT 2292.340 2.400 2292.480 24.830 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2273.465 13.685 2273.635 24.735 ;
      LAYER mcon ;
        RECT 2273.465 24.565 2273.635 24.735 ;
      LAYER met1 ;
        RECT 2099.970 1689.020 2100.290 1689.080 ;
        RECT 2103.650 1689.020 2103.970 1689.080 ;
        RECT 2099.970 1688.880 2103.970 1689.020 ;
        RECT 2099.970 1688.820 2100.290 1688.880 ;
        RECT 2103.650 1688.820 2103.970 1688.880 ;
        RECT 2103.650 24.720 2103.970 24.780 ;
        RECT 2273.405 24.720 2273.695 24.765 ;
        RECT 2103.650 24.580 2273.695 24.720 ;
        RECT 2103.650 24.520 2103.970 24.580 ;
        RECT 2273.405 24.535 2273.695 24.580 ;
        RECT 2273.405 13.840 2273.695 13.885 ;
        RECT 2310.190 13.840 2310.510 13.900 ;
        RECT 2273.405 13.700 2310.510 13.840 ;
        RECT 2273.405 13.655 2273.695 13.700 ;
        RECT 2310.190 13.640 2310.510 13.700 ;
      LAYER via ;
        RECT 2100.000 1688.820 2100.260 1689.080 ;
        RECT 2103.680 1688.820 2103.940 1689.080 ;
        RECT 2103.680 24.520 2103.940 24.780 ;
        RECT 2310.220 13.640 2310.480 13.900 ;
      LAYER met2 ;
        RECT 2099.925 1700.000 2100.205 1704.000 ;
        RECT 2100.060 1689.110 2100.200 1700.000 ;
        RECT 2100.000 1688.790 2100.260 1689.110 ;
        RECT 2103.680 1688.790 2103.940 1689.110 ;
        RECT 2103.740 24.810 2103.880 1688.790 ;
        RECT 2103.680 24.490 2103.940 24.810 ;
        RECT 2310.220 13.610 2310.480 13.930 ;
        RECT 2310.280 2.400 2310.420 13.610 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2306.125 24.225 2306.295 25.755 ;
      LAYER mcon ;
        RECT 2306.125 25.585 2306.295 25.755 ;
      LAYER met1 ;
        RECT 2107.330 1688.680 2107.650 1688.740 ;
        RECT 2111.010 1688.680 2111.330 1688.740 ;
        RECT 2107.330 1688.540 2111.330 1688.680 ;
        RECT 2107.330 1688.480 2107.650 1688.540 ;
        RECT 2111.010 1688.480 2111.330 1688.540 ;
        RECT 2306.065 25.740 2306.355 25.785 ;
        RECT 2306.065 25.600 2311.340 25.740 ;
        RECT 2306.065 25.555 2306.355 25.600 ;
        RECT 2311.200 25.060 2311.340 25.600 ;
        RECT 2328.130 25.060 2328.450 25.120 ;
        RECT 2311.200 24.920 2328.450 25.060 ;
        RECT 2328.130 24.860 2328.450 24.920 ;
        RECT 2111.010 24.380 2111.330 24.440 ;
        RECT 2306.065 24.380 2306.355 24.425 ;
        RECT 2111.010 24.240 2306.355 24.380 ;
        RECT 2111.010 24.180 2111.330 24.240 ;
        RECT 2306.065 24.195 2306.355 24.240 ;
      LAYER via ;
        RECT 2107.360 1688.480 2107.620 1688.740 ;
        RECT 2111.040 1688.480 2111.300 1688.740 ;
        RECT 2328.160 24.860 2328.420 25.120 ;
        RECT 2111.040 24.180 2111.300 24.440 ;
      LAYER met2 ;
        RECT 2107.285 1700.000 2107.565 1704.000 ;
        RECT 2107.420 1688.770 2107.560 1700.000 ;
        RECT 2107.360 1688.450 2107.620 1688.770 ;
        RECT 2111.040 1688.450 2111.300 1688.770 ;
        RECT 2111.100 24.470 2111.240 1688.450 ;
        RECT 2328.160 24.830 2328.420 25.150 ;
        RECT 2111.040 24.150 2111.300 24.470 ;
        RECT 2328.220 2.400 2328.360 24.830 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2345.610 24.380 2345.930 24.440 ;
        RECT 2307.980 24.240 2345.930 24.380 ;
        RECT 2117.910 24.040 2118.230 24.100 ;
        RECT 2307.980 24.040 2308.120 24.240 ;
        RECT 2345.610 24.180 2345.930 24.240 ;
        RECT 2117.910 23.900 2308.120 24.040 ;
        RECT 2117.910 23.840 2118.230 23.900 ;
      LAYER via ;
        RECT 2117.940 23.840 2118.200 24.100 ;
        RECT 2345.640 24.180 2345.900 24.440 ;
      LAYER met2 ;
        RECT 2114.645 1701.090 2114.925 1704.000 ;
        RECT 2114.645 1700.950 2117.220 1701.090 ;
        RECT 2114.645 1700.000 2114.925 1700.950 ;
        RECT 2117.080 1685.450 2117.220 1700.950 ;
        RECT 2117.080 1685.310 2118.140 1685.450 ;
        RECT 2118.000 24.130 2118.140 1685.310 ;
        RECT 2345.640 24.150 2345.900 24.470 ;
        RECT 2117.940 23.810 2118.200 24.130 ;
        RECT 2345.700 2.400 2345.840 24.150 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2124.810 20.980 2125.130 21.040 ;
        RECT 2363.550 20.980 2363.870 21.040 ;
        RECT 2124.810 20.840 2363.870 20.980 ;
        RECT 2124.810 20.780 2125.130 20.840 ;
        RECT 2363.550 20.780 2363.870 20.840 ;
      LAYER via ;
        RECT 2124.840 20.780 2125.100 21.040 ;
        RECT 2363.580 20.780 2363.840 21.040 ;
      LAYER met2 ;
        RECT 2122.005 1701.090 2122.285 1704.000 ;
        RECT 2122.005 1700.950 2124.580 1701.090 ;
        RECT 2122.005 1700.000 2122.285 1700.950 ;
        RECT 2124.440 1688.170 2124.580 1700.950 ;
        RECT 2124.440 1688.030 2125.040 1688.170 ;
        RECT 2124.900 21.070 2125.040 1688.030 ;
        RECT 2124.840 20.750 2125.100 21.070 ;
        RECT 2363.580 20.750 2363.840 21.070 ;
        RECT 2363.640 2.400 2363.780 20.750 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2131.710 28.800 2132.030 28.860 ;
        RECT 2381.490 28.800 2381.810 28.860 ;
        RECT 2131.710 28.660 2381.810 28.800 ;
        RECT 2131.710 28.600 2132.030 28.660 ;
        RECT 2381.490 28.600 2381.810 28.660 ;
      LAYER via ;
        RECT 2131.740 28.600 2132.000 28.860 ;
        RECT 2381.520 28.600 2381.780 28.860 ;
      LAYER met2 ;
        RECT 2129.365 1700.410 2129.645 1704.000 ;
        RECT 2129.365 1700.270 2131.940 1700.410 ;
        RECT 2129.365 1700.000 2129.645 1700.270 ;
        RECT 2131.800 28.890 2131.940 1700.270 ;
        RECT 2131.740 28.570 2132.000 28.890 ;
        RECT 2381.520 28.570 2381.780 28.890 ;
        RECT 2381.580 2.400 2381.720 28.570 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2138.610 29.140 2138.930 29.200 ;
        RECT 2399.430 29.140 2399.750 29.200 ;
        RECT 2138.610 29.000 2399.750 29.140 ;
        RECT 2138.610 28.940 2138.930 29.000 ;
        RECT 2399.430 28.940 2399.750 29.000 ;
      LAYER via ;
        RECT 2138.640 28.940 2138.900 29.200 ;
        RECT 2399.460 28.940 2399.720 29.200 ;
      LAYER met2 ;
        RECT 2136.725 1700.410 2137.005 1704.000 ;
        RECT 2136.725 1700.270 2138.840 1700.410 ;
        RECT 2136.725 1700.000 2137.005 1700.270 ;
        RECT 2138.700 29.230 2138.840 1700.270 ;
        RECT 2138.640 28.910 2138.900 29.230 ;
        RECT 2399.460 28.910 2399.720 29.230 ;
        RECT 2399.520 2.400 2399.660 28.910 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1471.225 1193.825 1471.395 1259.275 ;
        RECT 1472.145 565.845 1472.315 613.955 ;
        RECT 1471.225 324.445 1471.395 372.555 ;
      LAYER mcon ;
        RECT 1471.225 1259.105 1471.395 1259.275 ;
        RECT 1472.145 613.785 1472.315 613.955 ;
        RECT 1471.225 372.385 1471.395 372.555 ;
      LAYER met1 ;
        RECT 1471.150 1642.100 1471.470 1642.160 ;
        RECT 1472.070 1642.100 1472.390 1642.160 ;
        RECT 1471.150 1641.960 1472.390 1642.100 ;
        RECT 1471.150 1641.900 1471.470 1641.960 ;
        RECT 1472.070 1641.900 1472.390 1641.960 ;
        RECT 1471.150 1521.400 1471.470 1521.460 ;
        RECT 1472.070 1521.400 1472.390 1521.460 ;
        RECT 1471.150 1521.260 1472.390 1521.400 ;
        RECT 1471.150 1521.200 1471.470 1521.260 ;
        RECT 1472.070 1521.200 1472.390 1521.260 ;
        RECT 1471.150 1401.040 1471.470 1401.100 ;
        RECT 1471.610 1401.040 1471.930 1401.100 ;
        RECT 1471.150 1400.900 1471.930 1401.040 ;
        RECT 1471.150 1400.840 1471.470 1400.900 ;
        RECT 1471.610 1400.840 1471.930 1400.900 ;
        RECT 1471.150 1379.960 1471.470 1380.020 ;
        RECT 1471.610 1379.960 1471.930 1380.020 ;
        RECT 1471.150 1379.820 1471.930 1379.960 ;
        RECT 1471.150 1379.760 1471.470 1379.820 ;
        RECT 1471.610 1379.760 1471.930 1379.820 ;
        RECT 1471.610 1331.680 1471.930 1331.740 ;
        RECT 1472.070 1331.680 1472.390 1331.740 ;
        RECT 1471.610 1331.540 1472.390 1331.680 ;
        RECT 1471.610 1331.480 1471.930 1331.540 ;
        RECT 1472.070 1331.480 1472.390 1331.540 ;
        RECT 1471.165 1259.260 1471.455 1259.305 ;
        RECT 1472.070 1259.260 1472.390 1259.320 ;
        RECT 1471.165 1259.120 1472.390 1259.260 ;
        RECT 1471.165 1259.075 1471.455 1259.120 ;
        RECT 1472.070 1259.060 1472.390 1259.120 ;
        RECT 1471.165 1193.980 1471.455 1194.025 ;
        RECT 1472.070 1193.980 1472.390 1194.040 ;
        RECT 1471.165 1193.840 1472.390 1193.980 ;
        RECT 1471.165 1193.795 1471.455 1193.840 ;
        RECT 1472.070 1193.780 1472.390 1193.840 ;
        RECT 1471.610 1111.020 1471.930 1111.080 ;
        RECT 1472.070 1111.020 1472.390 1111.080 ;
        RECT 1471.610 1110.880 1472.390 1111.020 ;
        RECT 1471.610 1110.820 1471.930 1110.880 ;
        RECT 1472.070 1110.820 1472.390 1110.880 ;
        RECT 1471.150 1014.460 1471.470 1014.520 ;
        RECT 1471.610 1014.460 1471.930 1014.520 ;
        RECT 1471.150 1014.320 1471.930 1014.460 ;
        RECT 1471.150 1014.260 1471.470 1014.320 ;
        RECT 1471.610 1014.260 1471.930 1014.320 ;
        RECT 1471.150 893.760 1471.470 893.820 ;
        RECT 1472.070 893.760 1472.390 893.820 ;
        RECT 1471.150 893.620 1472.390 893.760 ;
        RECT 1471.150 893.560 1471.470 893.620 ;
        RECT 1472.070 893.560 1472.390 893.620 ;
        RECT 1471.610 807.400 1471.930 807.460 ;
        RECT 1472.070 807.400 1472.390 807.460 ;
        RECT 1471.610 807.260 1472.390 807.400 ;
        RECT 1471.610 807.200 1471.930 807.260 ;
        RECT 1472.070 807.200 1472.390 807.260 ;
        RECT 1471.150 765.920 1471.470 765.980 ;
        RECT 1471.610 765.920 1471.930 765.980 ;
        RECT 1471.150 765.780 1471.930 765.920 ;
        RECT 1471.150 765.720 1471.470 765.780 ;
        RECT 1471.610 765.720 1471.930 765.780 ;
        RECT 1472.070 613.940 1472.390 614.000 ;
        RECT 1471.875 613.800 1472.390 613.940 ;
        RECT 1472.070 613.740 1472.390 613.800 ;
        RECT 1472.070 566.000 1472.390 566.060 ;
        RECT 1471.875 565.860 1472.390 566.000 ;
        RECT 1472.070 565.800 1472.390 565.860 ;
        RECT 1472.070 517.520 1472.390 517.780 ;
        RECT 1472.160 517.380 1472.300 517.520 ;
        RECT 1472.990 517.380 1473.310 517.440 ;
        RECT 1472.160 517.240 1473.310 517.380 ;
        RECT 1472.990 517.180 1473.310 517.240 ;
        RECT 1472.070 427.960 1472.390 428.020 ;
        RECT 1472.990 427.960 1473.310 428.020 ;
        RECT 1472.070 427.820 1473.310 427.960 ;
        RECT 1472.070 427.760 1472.390 427.820 ;
        RECT 1472.990 427.760 1473.310 427.820 ;
        RECT 1471.165 372.540 1471.455 372.585 ;
        RECT 1472.070 372.540 1472.390 372.600 ;
        RECT 1471.165 372.400 1472.390 372.540 ;
        RECT 1471.165 372.355 1471.455 372.400 ;
        RECT 1472.070 372.340 1472.390 372.400 ;
        RECT 1471.150 324.600 1471.470 324.660 ;
        RECT 1470.955 324.460 1471.470 324.600 ;
        RECT 1471.150 324.400 1471.470 324.460 ;
        RECT 1470.690 179.420 1471.010 179.480 ;
        RECT 1472.530 179.420 1472.850 179.480 ;
        RECT 1470.690 179.280 1472.850 179.420 ;
        RECT 1470.690 179.220 1471.010 179.280 ;
        RECT 1472.530 179.220 1472.850 179.280 ;
        RECT 800.010 66.540 800.330 66.600 ;
        RECT 1472.070 66.540 1472.390 66.600 ;
        RECT 800.010 66.400 1472.390 66.540 ;
        RECT 800.010 66.340 800.330 66.400 ;
        RECT 1472.070 66.340 1472.390 66.400 ;
        RECT 793.570 20.980 793.890 21.040 ;
        RECT 800.010 20.980 800.330 21.040 ;
        RECT 793.570 20.840 800.330 20.980 ;
        RECT 793.570 20.780 793.890 20.840 ;
        RECT 800.010 20.780 800.330 20.840 ;
      LAYER via ;
        RECT 1471.180 1641.900 1471.440 1642.160 ;
        RECT 1472.100 1641.900 1472.360 1642.160 ;
        RECT 1471.180 1521.200 1471.440 1521.460 ;
        RECT 1472.100 1521.200 1472.360 1521.460 ;
        RECT 1471.180 1400.840 1471.440 1401.100 ;
        RECT 1471.640 1400.840 1471.900 1401.100 ;
        RECT 1471.180 1379.760 1471.440 1380.020 ;
        RECT 1471.640 1379.760 1471.900 1380.020 ;
        RECT 1471.640 1331.480 1471.900 1331.740 ;
        RECT 1472.100 1331.480 1472.360 1331.740 ;
        RECT 1472.100 1259.060 1472.360 1259.320 ;
        RECT 1472.100 1193.780 1472.360 1194.040 ;
        RECT 1471.640 1110.820 1471.900 1111.080 ;
        RECT 1472.100 1110.820 1472.360 1111.080 ;
        RECT 1471.180 1014.260 1471.440 1014.520 ;
        RECT 1471.640 1014.260 1471.900 1014.520 ;
        RECT 1471.180 893.560 1471.440 893.820 ;
        RECT 1472.100 893.560 1472.360 893.820 ;
        RECT 1471.640 807.200 1471.900 807.460 ;
        RECT 1472.100 807.200 1472.360 807.460 ;
        RECT 1471.180 765.720 1471.440 765.980 ;
        RECT 1471.640 765.720 1471.900 765.980 ;
        RECT 1472.100 613.740 1472.360 614.000 ;
        RECT 1472.100 565.800 1472.360 566.060 ;
        RECT 1472.100 517.520 1472.360 517.780 ;
        RECT 1473.020 517.180 1473.280 517.440 ;
        RECT 1472.100 427.760 1472.360 428.020 ;
        RECT 1473.020 427.760 1473.280 428.020 ;
        RECT 1472.100 372.340 1472.360 372.600 ;
        RECT 1471.180 324.400 1471.440 324.660 ;
        RECT 1470.720 179.220 1470.980 179.480 ;
        RECT 1472.560 179.220 1472.820 179.480 ;
        RECT 800.040 66.340 800.300 66.600 ;
        RECT 1472.100 66.340 1472.360 66.600 ;
        RECT 793.600 20.780 793.860 21.040 ;
        RECT 800.040 20.780 800.300 21.040 ;
      LAYER met2 ;
        RECT 1475.705 1701.090 1475.985 1704.000 ;
        RECT 1473.540 1700.950 1475.985 1701.090 ;
        RECT 1473.540 1677.970 1473.680 1700.950 ;
        RECT 1475.705 1700.000 1475.985 1700.950 ;
        RECT 1471.240 1677.830 1473.680 1677.970 ;
        RECT 1471.240 1642.190 1471.380 1677.830 ;
        RECT 1471.180 1641.870 1471.440 1642.190 ;
        RECT 1472.100 1641.870 1472.360 1642.190 ;
        RECT 1472.160 1617.450 1472.300 1641.870 ;
        RECT 1471.700 1617.310 1472.300 1617.450 ;
        RECT 1471.700 1563.050 1471.840 1617.310 ;
        RECT 1471.700 1562.910 1472.300 1563.050 ;
        RECT 1472.160 1521.490 1472.300 1562.910 ;
        RECT 1471.180 1521.170 1471.440 1521.490 ;
        RECT 1472.100 1521.170 1472.360 1521.490 ;
        RECT 1471.240 1466.490 1471.380 1521.170 ;
        RECT 1471.240 1466.350 1472.300 1466.490 ;
        RECT 1472.160 1448.980 1472.300 1466.350 ;
        RECT 1471.700 1448.840 1472.300 1448.980 ;
        RECT 1471.700 1401.130 1471.840 1448.840 ;
        RECT 1471.180 1400.810 1471.440 1401.130 ;
        RECT 1471.640 1400.810 1471.900 1401.130 ;
        RECT 1471.240 1380.050 1471.380 1400.810 ;
        RECT 1471.180 1379.730 1471.440 1380.050 ;
        RECT 1471.640 1379.730 1471.900 1380.050 ;
        RECT 1471.700 1331.770 1471.840 1379.730 ;
        RECT 1471.640 1331.450 1471.900 1331.770 ;
        RECT 1472.100 1331.450 1472.360 1331.770 ;
        RECT 1472.160 1259.350 1472.300 1331.450 ;
        RECT 1472.100 1259.030 1472.360 1259.350 ;
        RECT 1472.100 1193.750 1472.360 1194.070 ;
        RECT 1472.160 1111.110 1472.300 1193.750 ;
        RECT 1471.640 1110.790 1471.900 1111.110 ;
        RECT 1472.100 1110.790 1472.360 1111.110 ;
        RECT 1471.240 1014.550 1471.380 1014.705 ;
        RECT 1471.700 1014.550 1471.840 1110.790 ;
        RECT 1471.180 1014.290 1471.440 1014.550 ;
        RECT 1471.640 1014.290 1471.900 1014.550 ;
        RECT 1471.180 1014.230 1471.900 1014.290 ;
        RECT 1471.240 1014.150 1471.840 1014.230 ;
        RECT 1471.700 942.210 1471.840 1014.150 ;
        RECT 1471.240 942.070 1471.840 942.210 ;
        RECT 1471.240 893.850 1471.380 942.070 ;
        RECT 1471.180 893.530 1471.440 893.850 ;
        RECT 1472.100 893.530 1472.360 893.850 ;
        RECT 1472.160 807.490 1472.300 893.530 ;
        RECT 1471.640 807.170 1471.900 807.490 ;
        RECT 1472.100 807.170 1472.360 807.490 ;
        RECT 1471.700 766.010 1471.840 807.170 ;
        RECT 1471.180 765.690 1471.440 766.010 ;
        RECT 1471.640 765.690 1471.900 766.010 ;
        RECT 1471.240 686.530 1471.380 765.690 ;
        RECT 1471.240 686.390 1472.300 686.530 ;
        RECT 1472.160 614.030 1472.300 686.390 ;
        RECT 1472.100 613.710 1472.360 614.030 ;
        RECT 1472.100 565.770 1472.360 566.090 ;
        RECT 1472.160 517.810 1472.300 565.770 ;
        RECT 1472.100 517.490 1472.360 517.810 ;
        RECT 1473.020 517.150 1473.280 517.470 ;
        RECT 1473.080 428.050 1473.220 517.150 ;
        RECT 1472.100 427.730 1472.360 428.050 ;
        RECT 1473.020 427.730 1473.280 428.050 ;
        RECT 1472.160 372.630 1472.300 427.730 ;
        RECT 1472.100 372.310 1472.360 372.630 ;
        RECT 1471.180 324.370 1471.440 324.690 ;
        RECT 1471.240 227.645 1471.380 324.370 ;
        RECT 1471.170 227.275 1471.450 227.645 ;
        RECT 1470.710 179.675 1470.990 180.045 ;
        RECT 1470.780 179.510 1470.920 179.675 ;
        RECT 1470.720 179.190 1470.980 179.510 ;
        RECT 1472.560 179.190 1472.820 179.510 ;
        RECT 1472.620 96.460 1472.760 179.190 ;
        RECT 1472.160 96.320 1472.760 96.460 ;
        RECT 1472.160 66.630 1472.300 96.320 ;
        RECT 800.040 66.310 800.300 66.630 ;
        RECT 1472.100 66.310 1472.360 66.630 ;
        RECT 800.100 21.070 800.240 66.310 ;
        RECT 793.600 20.750 793.860 21.070 ;
        RECT 800.040 20.750 800.300 21.070 ;
        RECT 793.660 2.400 793.800 20.750 ;
        RECT 793.450 -4.800 794.010 2.400 ;
      LAYER via2 ;
        RECT 1471.170 227.320 1471.450 227.600 ;
        RECT 1470.710 179.720 1470.990 180.000 ;
      LAYER met3 ;
        RECT 1470.430 227.610 1470.810 227.620 ;
        RECT 1471.145 227.610 1471.475 227.625 ;
        RECT 1470.430 227.310 1471.475 227.610 ;
        RECT 1470.430 227.300 1470.810 227.310 ;
        RECT 1471.145 227.295 1471.475 227.310 ;
        RECT 1470.685 180.020 1471.015 180.025 ;
        RECT 1470.430 180.010 1471.015 180.020 ;
        RECT 1470.430 179.710 1471.240 180.010 ;
        RECT 1470.430 179.700 1471.015 179.710 ;
        RECT 1470.685 179.695 1471.015 179.700 ;
      LAYER via3 ;
        RECT 1470.460 227.300 1470.780 227.620 ;
        RECT 1470.460 179.700 1470.780 180.020 ;
      LAYER met4 ;
        RECT 1470.455 227.295 1470.785 227.625 ;
        RECT 1470.470 180.025 1470.770 227.295 ;
        RECT 1470.455 179.695 1470.785 180.025 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1408.665 1580.065 1408.835 1608.115 ;
        RECT 1409.125 1297.185 1409.295 1304.495 ;
        RECT 1409.125 1207.425 1409.295 1255.875 ;
        RECT 1408.665 717.825 1408.835 741.795 ;
        RECT 1409.125 379.525 1409.295 444.975 ;
        RECT 1408.665 241.485 1408.835 307.275 ;
        RECT 1408.665 144.925 1408.835 193.035 ;
      LAYER mcon ;
        RECT 1408.665 1607.945 1408.835 1608.115 ;
        RECT 1409.125 1304.325 1409.295 1304.495 ;
        RECT 1409.125 1255.705 1409.295 1255.875 ;
        RECT 1408.665 741.625 1408.835 741.795 ;
        RECT 1409.125 444.805 1409.295 444.975 ;
        RECT 1408.665 307.105 1408.835 307.275 ;
        RECT 1408.665 192.865 1408.835 193.035 ;
      LAYER met1 ;
        RECT 1408.605 1608.100 1408.895 1608.145 ;
        RECT 1409.050 1608.100 1409.370 1608.160 ;
        RECT 1408.605 1607.960 1409.370 1608.100 ;
        RECT 1408.605 1607.915 1408.895 1607.960 ;
        RECT 1409.050 1607.900 1409.370 1607.960 ;
        RECT 1408.590 1580.220 1408.910 1580.280 ;
        RECT 1408.395 1580.080 1408.910 1580.220 ;
        RECT 1408.590 1580.020 1408.910 1580.080 ;
        RECT 1408.590 1497.260 1408.910 1497.320 ;
        RECT 1409.050 1497.260 1409.370 1497.320 ;
        RECT 1408.590 1497.120 1409.370 1497.260 ;
        RECT 1408.590 1497.060 1408.910 1497.120 ;
        RECT 1409.050 1497.060 1409.370 1497.120 ;
        RECT 1408.590 1490.460 1408.910 1490.520 ;
        RECT 1409.050 1490.460 1409.370 1490.520 ;
        RECT 1408.590 1490.320 1409.370 1490.460 ;
        RECT 1408.590 1490.260 1408.910 1490.320 ;
        RECT 1409.050 1490.260 1409.370 1490.320 ;
        RECT 1408.590 1400.700 1408.910 1400.760 ;
        RECT 1409.050 1400.700 1409.370 1400.760 ;
        RECT 1408.590 1400.560 1409.370 1400.700 ;
        RECT 1408.590 1400.500 1408.910 1400.560 ;
        RECT 1409.050 1400.500 1409.370 1400.560 ;
        RECT 1409.050 1304.480 1409.370 1304.540 ;
        RECT 1408.855 1304.340 1409.370 1304.480 ;
        RECT 1409.050 1304.280 1409.370 1304.340 ;
        RECT 1409.050 1297.340 1409.370 1297.400 ;
        RECT 1408.855 1297.200 1409.370 1297.340 ;
        RECT 1409.050 1297.140 1409.370 1297.200 ;
        RECT 1409.050 1255.860 1409.370 1255.920 ;
        RECT 1408.855 1255.720 1409.370 1255.860 ;
        RECT 1409.050 1255.660 1409.370 1255.720 ;
        RECT 1409.050 1207.580 1409.370 1207.640 ;
        RECT 1408.855 1207.440 1409.370 1207.580 ;
        RECT 1409.050 1207.380 1409.370 1207.440 ;
        RECT 1409.050 1173.380 1409.370 1173.640 ;
        RECT 1409.140 1172.960 1409.280 1173.380 ;
        RECT 1409.050 1172.700 1409.370 1172.960 ;
        RECT 1408.590 1062.740 1408.910 1062.800 ;
        RECT 1409.510 1062.740 1409.830 1062.800 ;
        RECT 1408.590 1062.600 1409.830 1062.740 ;
        RECT 1408.590 1062.540 1408.910 1062.600 ;
        RECT 1409.510 1062.540 1409.830 1062.600 ;
        RECT 1408.590 1028.200 1408.910 1028.460 ;
        RECT 1408.680 1027.720 1408.820 1028.200 ;
        RECT 1409.050 1027.720 1409.370 1027.780 ;
        RECT 1408.680 1027.580 1409.370 1027.720 ;
        RECT 1409.050 1027.520 1409.370 1027.580 ;
        RECT 1408.590 966.180 1408.910 966.240 ;
        RECT 1409.510 966.180 1409.830 966.240 ;
        RECT 1408.590 966.040 1409.830 966.180 ;
        RECT 1408.590 965.980 1408.910 966.040 ;
        RECT 1409.510 965.980 1409.830 966.040 ;
        RECT 1408.590 869.620 1408.910 869.680 ;
        RECT 1409.510 869.620 1409.830 869.680 ;
        RECT 1408.590 869.480 1409.830 869.620 ;
        RECT 1408.590 869.420 1408.910 869.480 ;
        RECT 1409.510 869.420 1409.830 869.480 ;
        RECT 1408.590 741.780 1408.910 741.840 ;
        RECT 1408.395 741.640 1408.910 741.780 ;
        RECT 1408.590 741.580 1408.910 741.640 ;
        RECT 1408.590 717.980 1408.910 718.040 ;
        RECT 1408.395 717.840 1408.910 717.980 ;
        RECT 1408.590 717.780 1408.910 717.840 ;
        RECT 1408.590 444.960 1408.910 445.020 ;
        RECT 1409.065 444.960 1409.355 445.005 ;
        RECT 1408.590 444.820 1409.355 444.960 ;
        RECT 1408.590 444.760 1408.910 444.820 ;
        RECT 1409.065 444.775 1409.355 444.820 ;
        RECT 1409.050 379.680 1409.370 379.740 ;
        RECT 1408.855 379.540 1409.370 379.680 ;
        RECT 1409.050 379.480 1409.370 379.540 ;
        RECT 1408.590 338.200 1408.910 338.260 ;
        RECT 1409.050 338.200 1409.370 338.260 ;
        RECT 1408.590 338.060 1409.370 338.200 ;
        RECT 1408.590 338.000 1408.910 338.060 ;
        RECT 1409.050 338.000 1409.370 338.060 ;
        RECT 1408.590 307.260 1408.910 307.320 ;
        RECT 1408.395 307.120 1408.910 307.260 ;
        RECT 1408.590 307.060 1408.910 307.120 ;
        RECT 1408.590 241.640 1408.910 241.700 ;
        RECT 1408.395 241.500 1408.910 241.640 ;
        RECT 1408.590 241.440 1408.910 241.500 ;
        RECT 1408.590 193.020 1408.910 193.080 ;
        RECT 1408.395 192.880 1408.910 193.020 ;
        RECT 1408.590 192.820 1408.910 192.880 ;
        RECT 1408.590 145.080 1408.910 145.140 ;
        RECT 1408.395 144.940 1408.910 145.080 ;
        RECT 1408.590 144.880 1408.910 144.940 ;
        RECT 1408.590 97.140 1408.910 97.200 ;
        RECT 1408.220 97.000 1408.910 97.140 ;
        RECT 1408.220 96.860 1408.360 97.000 ;
        RECT 1408.590 96.940 1408.910 97.000 ;
        RECT 1408.130 96.600 1408.450 96.860 ;
        RECT 641.310 59.400 641.630 59.460 ;
        RECT 1408.130 59.400 1408.450 59.460 ;
        RECT 641.310 59.260 1408.450 59.400 ;
        RECT 641.310 59.200 641.630 59.260 ;
        RECT 1408.130 59.200 1408.450 59.260 ;
      LAYER via ;
        RECT 1409.080 1607.900 1409.340 1608.160 ;
        RECT 1408.620 1580.020 1408.880 1580.280 ;
        RECT 1408.620 1497.060 1408.880 1497.320 ;
        RECT 1409.080 1497.060 1409.340 1497.320 ;
        RECT 1408.620 1490.260 1408.880 1490.520 ;
        RECT 1409.080 1490.260 1409.340 1490.520 ;
        RECT 1408.620 1400.500 1408.880 1400.760 ;
        RECT 1409.080 1400.500 1409.340 1400.760 ;
        RECT 1409.080 1304.280 1409.340 1304.540 ;
        RECT 1409.080 1297.140 1409.340 1297.400 ;
        RECT 1409.080 1255.660 1409.340 1255.920 ;
        RECT 1409.080 1207.380 1409.340 1207.640 ;
        RECT 1409.080 1173.380 1409.340 1173.640 ;
        RECT 1409.080 1172.700 1409.340 1172.960 ;
        RECT 1408.620 1062.540 1408.880 1062.800 ;
        RECT 1409.540 1062.540 1409.800 1062.800 ;
        RECT 1408.620 1028.200 1408.880 1028.460 ;
        RECT 1409.080 1027.520 1409.340 1027.780 ;
        RECT 1408.620 965.980 1408.880 966.240 ;
        RECT 1409.540 965.980 1409.800 966.240 ;
        RECT 1408.620 869.420 1408.880 869.680 ;
        RECT 1409.540 869.420 1409.800 869.680 ;
        RECT 1408.620 741.580 1408.880 741.840 ;
        RECT 1408.620 717.780 1408.880 718.040 ;
        RECT 1408.620 444.760 1408.880 445.020 ;
        RECT 1409.080 379.480 1409.340 379.740 ;
        RECT 1408.620 338.000 1408.880 338.260 ;
        RECT 1409.080 338.000 1409.340 338.260 ;
        RECT 1408.620 307.060 1408.880 307.320 ;
        RECT 1408.620 241.440 1408.880 241.700 ;
        RECT 1408.620 192.820 1408.880 193.080 ;
        RECT 1408.620 144.880 1408.880 145.140 ;
        RECT 1408.620 96.940 1408.880 97.200 ;
        RECT 1408.160 96.600 1408.420 96.860 ;
        RECT 641.340 59.200 641.600 59.460 ;
        RECT 1408.160 59.200 1408.420 59.460 ;
      LAYER met2 ;
        RECT 1411.765 1701.090 1412.045 1704.000 ;
        RECT 1410.060 1700.950 1412.045 1701.090 ;
        RECT 1410.060 1678.140 1410.200 1700.950 ;
        RECT 1411.765 1700.000 1412.045 1700.950 ;
        RECT 1409.140 1678.000 1410.200 1678.140 ;
        RECT 1409.140 1608.190 1409.280 1678.000 ;
        RECT 1409.080 1607.870 1409.340 1608.190 ;
        RECT 1408.620 1579.990 1408.880 1580.310 ;
        RECT 1408.680 1556.250 1408.820 1579.990 ;
        RECT 1408.680 1556.110 1409.280 1556.250 ;
        RECT 1409.140 1497.350 1409.280 1556.110 ;
        RECT 1408.620 1497.030 1408.880 1497.350 ;
        RECT 1409.080 1497.030 1409.340 1497.350 ;
        RECT 1408.680 1490.550 1408.820 1497.030 ;
        RECT 1408.620 1490.230 1408.880 1490.550 ;
        RECT 1409.080 1490.230 1409.340 1490.550 ;
        RECT 1409.140 1400.790 1409.280 1490.230 ;
        RECT 1408.620 1400.470 1408.880 1400.790 ;
        RECT 1409.080 1400.470 1409.340 1400.790 ;
        RECT 1408.680 1393.845 1408.820 1400.470 ;
        RECT 1408.610 1393.475 1408.890 1393.845 ;
        RECT 1409.070 1392.795 1409.350 1393.165 ;
        RECT 1409.140 1304.570 1409.280 1392.795 ;
        RECT 1409.080 1304.250 1409.340 1304.570 ;
        RECT 1409.080 1297.110 1409.340 1297.430 ;
        RECT 1409.140 1255.950 1409.280 1297.110 ;
        RECT 1409.080 1255.630 1409.340 1255.950 ;
        RECT 1409.080 1207.350 1409.340 1207.670 ;
        RECT 1409.140 1173.670 1409.280 1207.350 ;
        RECT 1409.080 1173.350 1409.340 1173.670 ;
        RECT 1409.080 1172.670 1409.340 1172.990 ;
        RECT 1409.140 1087.050 1409.280 1172.670 ;
        RECT 1409.140 1086.910 1409.740 1087.050 ;
        RECT 1409.600 1062.830 1409.740 1086.910 ;
        RECT 1408.620 1062.510 1408.880 1062.830 ;
        RECT 1409.540 1062.510 1409.800 1062.830 ;
        RECT 1408.680 1028.490 1408.820 1062.510 ;
        RECT 1408.620 1028.170 1408.880 1028.490 ;
        RECT 1409.080 1027.490 1409.340 1027.810 ;
        RECT 1409.140 990.490 1409.280 1027.490 ;
        RECT 1409.140 990.350 1409.740 990.490 ;
        RECT 1409.600 966.270 1409.740 990.350 ;
        RECT 1408.620 966.125 1408.880 966.270 ;
        RECT 1409.540 966.125 1409.800 966.270 ;
        RECT 1408.610 965.755 1408.890 966.125 ;
        RECT 1409.530 965.755 1409.810 966.125 ;
        RECT 1409.600 931.330 1409.740 965.755 ;
        RECT 1409.140 931.190 1409.740 931.330 ;
        RECT 1409.140 893.930 1409.280 931.190 ;
        RECT 1409.140 893.790 1409.740 893.930 ;
        RECT 1409.600 869.710 1409.740 893.790 ;
        RECT 1408.620 869.565 1408.880 869.710 ;
        RECT 1409.540 869.565 1409.800 869.710 ;
        RECT 1408.610 869.195 1408.890 869.565 ;
        RECT 1409.530 869.195 1409.810 869.565 ;
        RECT 1409.600 834.090 1409.740 869.195 ;
        RECT 1409.140 833.950 1409.740 834.090 ;
        RECT 1409.140 787.170 1409.280 833.950 ;
        RECT 1408.680 787.030 1409.280 787.170 ;
        RECT 1408.680 741.870 1408.820 787.030 ;
        RECT 1408.620 741.550 1408.880 741.870 ;
        RECT 1408.620 717.750 1408.880 718.070 ;
        RECT 1408.680 628.845 1408.820 717.750 ;
        RECT 1408.610 628.475 1408.890 628.845 ;
        RECT 1408.610 627.795 1408.890 628.165 ;
        RECT 1408.680 610.370 1408.820 627.795 ;
        RECT 1408.680 610.230 1409.740 610.370 ;
        RECT 1409.600 592.690 1409.740 610.230 ;
        RECT 1409.140 592.550 1409.740 592.690 ;
        RECT 1409.140 502.930 1409.280 592.550 ;
        RECT 1408.680 502.790 1409.280 502.930 ;
        RECT 1408.680 445.050 1408.820 502.790 ;
        RECT 1408.620 444.730 1408.880 445.050 ;
        RECT 1409.080 379.450 1409.340 379.770 ;
        RECT 1409.140 338.290 1409.280 379.450 ;
        RECT 1408.620 337.970 1408.880 338.290 ;
        RECT 1409.080 337.970 1409.340 338.290 ;
        RECT 1408.680 307.350 1408.820 337.970 ;
        RECT 1408.620 307.030 1408.880 307.350 ;
        RECT 1408.620 241.410 1408.880 241.730 ;
        RECT 1408.680 193.110 1408.820 241.410 ;
        RECT 1408.620 192.790 1408.880 193.110 ;
        RECT 1408.620 144.850 1408.880 145.170 ;
        RECT 1408.680 97.230 1408.820 144.850 ;
        RECT 1408.620 96.910 1408.880 97.230 ;
        RECT 1408.160 96.570 1408.420 96.890 ;
        RECT 1408.220 59.490 1408.360 96.570 ;
        RECT 641.340 59.170 641.600 59.490 ;
        RECT 1408.160 59.170 1408.420 59.490 ;
        RECT 641.400 17.410 641.540 59.170 ;
        RECT 639.100 17.270 641.540 17.410 ;
        RECT 639.100 2.400 639.240 17.270 ;
        RECT 638.890 -4.800 639.450 2.400 ;
      LAYER via2 ;
        RECT 1408.610 1393.520 1408.890 1393.800 ;
        RECT 1409.070 1392.840 1409.350 1393.120 ;
        RECT 1408.610 965.800 1408.890 966.080 ;
        RECT 1409.530 965.800 1409.810 966.080 ;
        RECT 1408.610 869.240 1408.890 869.520 ;
        RECT 1409.530 869.240 1409.810 869.520 ;
        RECT 1408.610 628.520 1408.890 628.800 ;
        RECT 1408.610 627.840 1408.890 628.120 ;
      LAYER met3 ;
        RECT 1408.585 1393.810 1408.915 1393.825 ;
        RECT 1407.910 1393.510 1408.915 1393.810 ;
        RECT 1407.910 1393.130 1408.210 1393.510 ;
        RECT 1408.585 1393.495 1408.915 1393.510 ;
        RECT 1409.045 1393.130 1409.375 1393.145 ;
        RECT 1407.910 1392.830 1409.375 1393.130 ;
        RECT 1409.045 1392.815 1409.375 1392.830 ;
        RECT 1408.585 966.090 1408.915 966.105 ;
        RECT 1409.505 966.090 1409.835 966.105 ;
        RECT 1408.585 965.790 1409.835 966.090 ;
        RECT 1408.585 965.775 1408.915 965.790 ;
        RECT 1409.505 965.775 1409.835 965.790 ;
        RECT 1408.585 869.530 1408.915 869.545 ;
        RECT 1409.505 869.530 1409.835 869.545 ;
        RECT 1408.585 869.230 1409.835 869.530 ;
        RECT 1408.585 869.215 1408.915 869.230 ;
        RECT 1409.505 869.215 1409.835 869.230 ;
        RECT 1408.585 628.810 1408.915 628.825 ;
        RECT 1408.585 628.495 1409.130 628.810 ;
        RECT 1408.830 628.145 1409.130 628.495 ;
        RECT 1408.585 627.830 1409.130 628.145 ;
        RECT 1408.585 627.815 1408.915 627.830 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2146.890 1683.920 2147.210 1683.980 ;
        RECT 2151.950 1683.920 2152.270 1683.980 ;
        RECT 2146.890 1683.780 2152.270 1683.920 ;
        RECT 2146.890 1683.720 2147.210 1683.780 ;
        RECT 2151.950 1683.720 2152.270 1683.780 ;
        RECT 2151.950 29.820 2152.270 29.880 ;
        RECT 2422.890 29.820 2423.210 29.880 ;
        RECT 2151.950 29.680 2423.210 29.820 ;
        RECT 2151.950 29.620 2152.270 29.680 ;
        RECT 2422.890 29.620 2423.210 29.680 ;
      LAYER via ;
        RECT 2146.920 1683.720 2147.180 1683.980 ;
        RECT 2151.980 1683.720 2152.240 1683.980 ;
        RECT 2151.980 29.620 2152.240 29.880 ;
        RECT 2422.920 29.620 2423.180 29.880 ;
      LAYER met2 ;
        RECT 2146.845 1700.000 2147.125 1704.000 ;
        RECT 2146.980 1684.010 2147.120 1700.000 ;
        RECT 2146.920 1683.690 2147.180 1684.010 ;
        RECT 2151.980 1683.690 2152.240 1684.010 ;
        RECT 2152.040 29.910 2152.180 1683.690 ;
        RECT 2151.980 29.590 2152.240 29.910 ;
        RECT 2422.920 29.590 2423.180 29.910 ;
        RECT 2422.980 2.400 2423.120 29.590 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2154.250 1683.920 2154.570 1683.980 ;
        RECT 2158.850 1683.920 2159.170 1683.980 ;
        RECT 2154.250 1683.780 2159.170 1683.920 ;
        RECT 2154.250 1683.720 2154.570 1683.780 ;
        RECT 2158.850 1683.720 2159.170 1683.780 ;
        RECT 2158.850 30.500 2159.170 30.560 ;
        RECT 2440.830 30.500 2441.150 30.560 ;
        RECT 2158.850 30.360 2441.150 30.500 ;
        RECT 2158.850 30.300 2159.170 30.360 ;
        RECT 2440.830 30.300 2441.150 30.360 ;
      LAYER via ;
        RECT 2154.280 1683.720 2154.540 1683.980 ;
        RECT 2158.880 1683.720 2159.140 1683.980 ;
        RECT 2158.880 30.300 2159.140 30.560 ;
        RECT 2440.860 30.300 2441.120 30.560 ;
      LAYER met2 ;
        RECT 2154.205 1700.000 2154.485 1704.000 ;
        RECT 2154.340 1684.010 2154.480 1700.000 ;
        RECT 2154.280 1683.690 2154.540 1684.010 ;
        RECT 2158.880 1683.690 2159.140 1684.010 ;
        RECT 2158.940 30.590 2159.080 1683.690 ;
        RECT 2158.880 30.270 2159.140 30.590 ;
        RECT 2440.860 30.270 2441.120 30.590 ;
        RECT 2440.920 2.400 2441.060 30.270 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2161.610 1683.920 2161.930 1683.980 ;
        RECT 2165.750 1683.920 2166.070 1683.980 ;
        RECT 2161.610 1683.780 2166.070 1683.920 ;
        RECT 2161.610 1683.720 2161.930 1683.780 ;
        RECT 2165.750 1683.720 2166.070 1683.780 ;
        RECT 2165.750 33.900 2166.070 33.960 ;
        RECT 2458.770 33.900 2459.090 33.960 ;
        RECT 2165.750 33.760 2459.090 33.900 ;
        RECT 2165.750 33.700 2166.070 33.760 ;
        RECT 2458.770 33.700 2459.090 33.760 ;
      LAYER via ;
        RECT 2161.640 1683.720 2161.900 1683.980 ;
        RECT 2165.780 1683.720 2166.040 1683.980 ;
        RECT 2165.780 33.700 2166.040 33.960 ;
        RECT 2458.800 33.700 2459.060 33.960 ;
      LAYER met2 ;
        RECT 2161.565 1700.000 2161.845 1704.000 ;
        RECT 2161.700 1684.010 2161.840 1700.000 ;
        RECT 2161.640 1683.690 2161.900 1684.010 ;
        RECT 2165.780 1683.690 2166.040 1684.010 ;
        RECT 2165.840 33.990 2165.980 1683.690 ;
        RECT 2165.780 33.670 2166.040 33.990 ;
        RECT 2458.800 33.670 2459.060 33.990 ;
        RECT 2458.860 2.400 2459.000 33.670 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2168.510 1683.920 2168.830 1683.980 ;
        RECT 2173.110 1683.920 2173.430 1683.980 ;
        RECT 2168.510 1683.780 2173.430 1683.920 ;
        RECT 2168.510 1683.720 2168.830 1683.780 ;
        RECT 2173.110 1683.720 2173.430 1683.780 ;
        RECT 2173.110 33.560 2173.430 33.620 ;
        RECT 2476.710 33.560 2477.030 33.620 ;
        RECT 2173.110 33.420 2477.030 33.560 ;
        RECT 2173.110 33.360 2173.430 33.420 ;
        RECT 2476.710 33.360 2477.030 33.420 ;
      LAYER via ;
        RECT 2168.540 1683.720 2168.800 1683.980 ;
        RECT 2173.140 1683.720 2173.400 1683.980 ;
        RECT 2173.140 33.360 2173.400 33.620 ;
        RECT 2476.740 33.360 2477.000 33.620 ;
      LAYER met2 ;
        RECT 2168.465 1700.000 2168.745 1704.000 ;
        RECT 2168.600 1684.010 2168.740 1700.000 ;
        RECT 2168.540 1683.690 2168.800 1684.010 ;
        RECT 2173.140 1683.690 2173.400 1684.010 ;
        RECT 2173.200 33.650 2173.340 1683.690 ;
        RECT 2173.140 33.330 2173.400 33.650 ;
        RECT 2476.740 33.330 2477.000 33.650 ;
        RECT 2476.800 2.400 2476.940 33.330 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2175.870 1683.920 2176.190 1683.980 ;
        RECT 2180.010 1683.920 2180.330 1683.980 ;
        RECT 2175.870 1683.780 2180.330 1683.920 ;
        RECT 2175.870 1683.720 2176.190 1683.780 ;
        RECT 2180.010 1683.720 2180.330 1683.780 ;
        RECT 2180.010 32.540 2180.330 32.600 ;
        RECT 2494.650 32.540 2494.970 32.600 ;
        RECT 2180.010 32.400 2494.970 32.540 ;
        RECT 2180.010 32.340 2180.330 32.400 ;
        RECT 2494.650 32.340 2494.970 32.400 ;
      LAYER via ;
        RECT 2175.900 1683.720 2176.160 1683.980 ;
        RECT 2180.040 1683.720 2180.300 1683.980 ;
        RECT 2180.040 32.340 2180.300 32.600 ;
        RECT 2494.680 32.340 2494.940 32.600 ;
      LAYER met2 ;
        RECT 2175.825 1700.000 2176.105 1704.000 ;
        RECT 2175.960 1684.010 2176.100 1700.000 ;
        RECT 2175.900 1683.690 2176.160 1684.010 ;
        RECT 2180.040 1683.690 2180.300 1684.010 ;
        RECT 2180.100 32.630 2180.240 1683.690 ;
        RECT 2180.040 32.310 2180.300 32.630 ;
        RECT 2494.680 32.310 2494.940 32.630 ;
        RECT 2494.740 2.400 2494.880 32.310 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2183.230 1688.000 2183.550 1688.060 ;
        RECT 2186.450 1688.000 2186.770 1688.060 ;
        RECT 2183.230 1687.860 2186.770 1688.000 ;
        RECT 2183.230 1687.800 2183.550 1687.860 ;
        RECT 2186.450 1687.800 2186.770 1687.860 ;
        RECT 2186.450 31.860 2186.770 31.920 ;
        RECT 2512.130 31.860 2512.450 31.920 ;
        RECT 2186.450 31.720 2512.450 31.860 ;
        RECT 2186.450 31.660 2186.770 31.720 ;
        RECT 2512.130 31.660 2512.450 31.720 ;
      LAYER via ;
        RECT 2183.260 1687.800 2183.520 1688.060 ;
        RECT 2186.480 1687.800 2186.740 1688.060 ;
        RECT 2186.480 31.660 2186.740 31.920 ;
        RECT 2512.160 31.660 2512.420 31.920 ;
      LAYER met2 ;
        RECT 2183.185 1700.000 2183.465 1704.000 ;
        RECT 2183.320 1688.090 2183.460 1700.000 ;
        RECT 2183.260 1687.770 2183.520 1688.090 ;
        RECT 2186.480 1687.770 2186.740 1688.090 ;
        RECT 2186.540 31.950 2186.680 1687.770 ;
        RECT 2186.480 31.630 2186.740 31.950 ;
        RECT 2512.160 31.630 2512.420 31.950 ;
        RECT 2512.220 2.400 2512.360 31.630 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2193.810 31.180 2194.130 31.240 ;
        RECT 2530.070 31.180 2530.390 31.240 ;
        RECT 2193.810 31.040 2530.390 31.180 ;
        RECT 2193.810 30.980 2194.130 31.040 ;
        RECT 2530.070 30.980 2530.390 31.040 ;
      LAYER via ;
        RECT 2193.840 30.980 2194.100 31.240 ;
        RECT 2530.100 30.980 2530.360 31.240 ;
      LAYER met2 ;
        RECT 2190.545 1700.410 2190.825 1704.000 ;
        RECT 2190.545 1700.270 2193.120 1700.410 ;
        RECT 2190.545 1700.000 2190.825 1700.270 ;
        RECT 2192.980 1688.680 2193.120 1700.270 ;
        RECT 2192.980 1688.540 2194.040 1688.680 ;
        RECT 2193.900 31.270 2194.040 1688.540 ;
        RECT 2193.840 30.950 2194.100 31.270 ;
        RECT 2530.100 30.950 2530.360 31.270 ;
        RECT 2530.160 2.400 2530.300 30.950 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2200.250 36.620 2200.570 36.680 ;
        RECT 2548.010 36.620 2548.330 36.680 ;
        RECT 2200.250 36.480 2548.330 36.620 ;
        RECT 2200.250 36.420 2200.570 36.480 ;
        RECT 2548.010 36.420 2548.330 36.480 ;
      LAYER via ;
        RECT 2200.280 36.420 2200.540 36.680 ;
        RECT 2548.040 36.420 2548.300 36.680 ;
      LAYER met2 ;
        RECT 2197.905 1700.410 2198.185 1704.000 ;
        RECT 2197.905 1700.270 2200.480 1700.410 ;
        RECT 2197.905 1700.000 2198.185 1700.270 ;
        RECT 2200.340 36.710 2200.480 1700.270 ;
        RECT 2200.280 36.390 2200.540 36.710 ;
        RECT 2548.040 36.390 2548.300 36.710 ;
        RECT 2548.100 2.400 2548.240 36.390 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2207.150 36.960 2207.470 37.020 ;
        RECT 2565.950 36.960 2566.270 37.020 ;
        RECT 2207.150 36.820 2566.270 36.960 ;
        RECT 2207.150 36.760 2207.470 36.820 ;
        RECT 2565.950 36.760 2566.270 36.820 ;
      LAYER via ;
        RECT 2207.180 36.760 2207.440 37.020 ;
        RECT 2565.980 36.760 2566.240 37.020 ;
      LAYER met2 ;
        RECT 2205.265 1700.410 2205.545 1704.000 ;
        RECT 2205.265 1700.270 2207.380 1700.410 ;
        RECT 2205.265 1700.000 2205.545 1700.270 ;
        RECT 2207.240 37.050 2207.380 1700.270 ;
        RECT 2207.180 36.730 2207.440 37.050 ;
        RECT 2565.980 36.730 2566.240 37.050 ;
        RECT 2566.040 2.400 2566.180 36.730 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2214.050 37.300 2214.370 37.360 ;
        RECT 2583.890 37.300 2584.210 37.360 ;
        RECT 2214.050 37.160 2584.210 37.300 ;
        RECT 2214.050 37.100 2214.370 37.160 ;
        RECT 2583.890 37.100 2584.210 37.160 ;
      LAYER via ;
        RECT 2214.080 37.100 2214.340 37.360 ;
        RECT 2583.920 37.100 2584.180 37.360 ;
      LAYER met2 ;
        RECT 2212.625 1700.410 2212.905 1704.000 ;
        RECT 2212.625 1700.270 2214.280 1700.410 ;
        RECT 2212.625 1700.000 2212.905 1700.270 ;
        RECT 2214.140 37.390 2214.280 1700.270 ;
        RECT 2214.080 37.070 2214.340 37.390 ;
        RECT 2583.920 37.070 2584.180 37.390 ;
        RECT 2583.980 2.400 2584.120 37.070 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 817.490 33.560 817.810 33.620 ;
        RECT 1483.570 33.560 1483.890 33.620 ;
        RECT 817.490 33.420 1483.890 33.560 ;
        RECT 817.490 33.360 817.810 33.420 ;
        RECT 1483.570 33.360 1483.890 33.420 ;
      LAYER via ;
        RECT 817.520 33.360 817.780 33.620 ;
        RECT 1483.600 33.360 1483.860 33.620 ;
      LAYER met2 ;
        RECT 1485.365 1700.410 1485.645 1704.000 ;
        RECT 1483.660 1700.270 1485.645 1700.410 ;
        RECT 1483.660 33.650 1483.800 1700.270 ;
        RECT 1485.365 1700.000 1485.645 1700.270 ;
        RECT 817.520 33.330 817.780 33.650 ;
        RECT 1483.600 33.330 1483.860 33.650 ;
        RECT 817.580 2.400 817.720 33.330 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2220.950 37.640 2221.270 37.700 ;
        RECT 2601.370 37.640 2601.690 37.700 ;
        RECT 2220.950 37.500 2601.690 37.640 ;
        RECT 2220.950 37.440 2221.270 37.500 ;
        RECT 2601.370 37.440 2601.690 37.500 ;
      LAYER via ;
        RECT 2220.980 37.440 2221.240 37.700 ;
        RECT 2601.400 37.440 2601.660 37.700 ;
      LAYER met2 ;
        RECT 2219.985 1700.410 2220.265 1704.000 ;
        RECT 2219.985 1700.270 2221.180 1700.410 ;
        RECT 2219.985 1700.000 2220.265 1700.270 ;
        RECT 2221.040 37.730 2221.180 1700.270 ;
        RECT 2220.980 37.410 2221.240 37.730 ;
        RECT 2601.400 37.410 2601.660 37.730 ;
        RECT 2601.460 2.400 2601.600 37.410 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2227.390 41.380 2227.710 41.440 ;
        RECT 2619.310 41.380 2619.630 41.440 ;
        RECT 2227.390 41.240 2619.630 41.380 ;
        RECT 2227.390 41.180 2227.710 41.240 ;
        RECT 2619.310 41.180 2619.630 41.240 ;
      LAYER via ;
        RECT 2227.420 41.180 2227.680 41.440 ;
        RECT 2619.340 41.180 2619.600 41.440 ;
      LAYER met2 ;
        RECT 2227.345 1700.000 2227.625 1704.000 ;
        RECT 2227.480 41.470 2227.620 1700.000 ;
        RECT 2227.420 41.150 2227.680 41.470 ;
        RECT 2619.340 41.150 2619.600 41.470 ;
        RECT 2619.400 2.400 2619.540 41.150 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2234.750 41.040 2235.070 41.100 ;
        RECT 2637.250 41.040 2637.570 41.100 ;
        RECT 2234.750 40.900 2637.570 41.040 ;
        RECT 2234.750 40.840 2235.070 40.900 ;
        RECT 2637.250 40.840 2637.570 40.900 ;
      LAYER via ;
        RECT 2234.780 40.840 2235.040 41.100 ;
        RECT 2637.280 40.840 2637.540 41.100 ;
      LAYER met2 ;
        RECT 2234.705 1700.000 2234.985 1704.000 ;
        RECT 2234.840 41.130 2234.980 1700.000 ;
        RECT 2234.780 40.810 2235.040 41.130 ;
        RECT 2637.280 40.810 2637.540 41.130 ;
        RECT 2637.340 2.400 2637.480 40.810 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2241.190 1688.340 2241.510 1688.400 ;
        RECT 2242.110 1688.340 2242.430 1688.400 ;
        RECT 2241.190 1688.200 2242.430 1688.340 ;
        RECT 2241.190 1688.140 2241.510 1688.200 ;
        RECT 2242.110 1688.140 2242.430 1688.200 ;
        RECT 2241.190 40.700 2241.510 40.760 ;
        RECT 2655.190 40.700 2655.510 40.760 ;
        RECT 2241.190 40.560 2655.510 40.700 ;
        RECT 2241.190 40.500 2241.510 40.560 ;
        RECT 2655.190 40.500 2655.510 40.560 ;
      LAYER via ;
        RECT 2241.220 1688.140 2241.480 1688.400 ;
        RECT 2242.140 1688.140 2242.400 1688.400 ;
        RECT 2241.220 40.500 2241.480 40.760 ;
        RECT 2655.220 40.500 2655.480 40.760 ;
      LAYER met2 ;
        RECT 2242.065 1700.000 2242.345 1704.000 ;
        RECT 2242.200 1688.430 2242.340 1700.000 ;
        RECT 2241.220 1688.110 2241.480 1688.430 ;
        RECT 2242.140 1688.110 2242.400 1688.430 ;
        RECT 2241.280 40.790 2241.420 1688.110 ;
        RECT 2241.220 40.470 2241.480 40.790 ;
        RECT 2655.220 40.470 2655.480 40.790 ;
        RECT 2655.280 2.400 2655.420 40.470 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2249.470 1688.340 2249.790 1688.400 ;
        RECT 2254.990 1688.340 2255.310 1688.400 ;
        RECT 2249.470 1688.200 2255.310 1688.340 ;
        RECT 2249.470 1688.140 2249.790 1688.200 ;
        RECT 2254.990 1688.140 2255.310 1688.200 ;
        RECT 2254.990 40.360 2255.310 40.420 ;
        RECT 2672.670 40.360 2672.990 40.420 ;
        RECT 2254.990 40.220 2672.990 40.360 ;
        RECT 2254.990 40.160 2255.310 40.220 ;
        RECT 2672.670 40.160 2672.990 40.220 ;
      LAYER via ;
        RECT 2249.500 1688.140 2249.760 1688.400 ;
        RECT 2255.020 1688.140 2255.280 1688.400 ;
        RECT 2255.020 40.160 2255.280 40.420 ;
        RECT 2672.700 40.160 2672.960 40.420 ;
      LAYER met2 ;
        RECT 2249.425 1700.000 2249.705 1704.000 ;
        RECT 2249.560 1688.430 2249.700 1700.000 ;
        RECT 2249.500 1688.110 2249.760 1688.430 ;
        RECT 2255.020 1688.110 2255.280 1688.430 ;
        RECT 2255.080 40.450 2255.220 1688.110 ;
        RECT 2255.020 40.130 2255.280 40.450 ;
        RECT 2672.700 40.130 2672.960 40.450 ;
        RECT 2672.760 2.400 2672.900 40.130 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2256.830 1688.340 2257.150 1688.400 ;
        RECT 2262.350 1688.340 2262.670 1688.400 ;
        RECT 2256.830 1688.200 2262.670 1688.340 ;
        RECT 2256.830 1688.140 2257.150 1688.200 ;
        RECT 2262.350 1688.140 2262.670 1688.200 ;
        RECT 2262.350 40.020 2262.670 40.080 ;
        RECT 2690.610 40.020 2690.930 40.080 ;
        RECT 2262.350 39.880 2690.930 40.020 ;
        RECT 2262.350 39.820 2262.670 39.880 ;
        RECT 2690.610 39.820 2690.930 39.880 ;
      LAYER via ;
        RECT 2256.860 1688.140 2257.120 1688.400 ;
        RECT 2262.380 1688.140 2262.640 1688.400 ;
        RECT 2262.380 39.820 2262.640 40.080 ;
        RECT 2690.640 39.820 2690.900 40.080 ;
      LAYER met2 ;
        RECT 2256.785 1700.000 2257.065 1704.000 ;
        RECT 2256.920 1688.430 2257.060 1700.000 ;
        RECT 2256.860 1688.110 2257.120 1688.430 ;
        RECT 2262.380 1688.110 2262.640 1688.430 ;
        RECT 2262.440 40.110 2262.580 1688.110 ;
        RECT 2262.380 39.790 2262.640 40.110 ;
        RECT 2690.640 39.790 2690.900 40.110 ;
        RECT 2690.700 2.400 2690.840 39.790 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2264.190 1688.340 2264.510 1688.400 ;
        RECT 2268.790 1688.340 2269.110 1688.400 ;
        RECT 2264.190 1688.200 2269.110 1688.340 ;
        RECT 2264.190 1688.140 2264.510 1688.200 ;
        RECT 2268.790 1688.140 2269.110 1688.200 ;
        RECT 2268.790 39.680 2269.110 39.740 ;
        RECT 2708.550 39.680 2708.870 39.740 ;
        RECT 2268.790 39.540 2708.870 39.680 ;
        RECT 2268.790 39.480 2269.110 39.540 ;
        RECT 2708.550 39.480 2708.870 39.540 ;
      LAYER via ;
        RECT 2264.220 1688.140 2264.480 1688.400 ;
        RECT 2268.820 1688.140 2269.080 1688.400 ;
        RECT 2268.820 39.480 2269.080 39.740 ;
        RECT 2708.580 39.480 2708.840 39.740 ;
      LAYER met2 ;
        RECT 2264.145 1700.000 2264.425 1704.000 ;
        RECT 2264.280 1688.430 2264.420 1700.000 ;
        RECT 2264.220 1688.110 2264.480 1688.430 ;
        RECT 2268.820 1688.110 2269.080 1688.430 ;
        RECT 2268.880 39.770 2269.020 1688.110 ;
        RECT 2268.820 39.450 2269.080 39.770 ;
        RECT 2708.580 39.450 2708.840 39.770 ;
        RECT 2708.640 2.400 2708.780 39.450 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2271.550 1688.340 2271.870 1688.400 ;
        RECT 2276.150 1688.340 2276.470 1688.400 ;
        RECT 2271.550 1688.200 2276.470 1688.340 ;
        RECT 2271.550 1688.140 2271.870 1688.200 ;
        RECT 2276.150 1688.140 2276.470 1688.200 ;
        RECT 2276.150 39.340 2276.470 39.400 ;
        RECT 2726.490 39.340 2726.810 39.400 ;
        RECT 2276.150 39.200 2726.810 39.340 ;
        RECT 2276.150 39.140 2276.470 39.200 ;
        RECT 2726.490 39.140 2726.810 39.200 ;
      LAYER via ;
        RECT 2271.580 1688.140 2271.840 1688.400 ;
        RECT 2276.180 1688.140 2276.440 1688.400 ;
        RECT 2276.180 39.140 2276.440 39.400 ;
        RECT 2726.520 39.140 2726.780 39.400 ;
      LAYER met2 ;
        RECT 2271.505 1700.000 2271.785 1704.000 ;
        RECT 2271.640 1688.430 2271.780 1700.000 ;
        RECT 2271.580 1688.110 2271.840 1688.430 ;
        RECT 2276.180 1688.110 2276.440 1688.430 ;
        RECT 2276.240 39.430 2276.380 1688.110 ;
        RECT 2276.180 39.110 2276.440 39.430 ;
        RECT 2726.520 39.110 2726.780 39.430 ;
        RECT 2726.580 2.400 2726.720 39.110 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2278.910 1688.340 2279.230 1688.400 ;
        RECT 2283.050 1688.340 2283.370 1688.400 ;
        RECT 2278.910 1688.200 2283.370 1688.340 ;
        RECT 2278.910 1688.140 2279.230 1688.200 ;
        RECT 2283.050 1688.140 2283.370 1688.200 ;
        RECT 2283.050 39.000 2283.370 39.060 ;
        RECT 2744.430 39.000 2744.750 39.060 ;
        RECT 2283.050 38.860 2744.750 39.000 ;
        RECT 2283.050 38.800 2283.370 38.860 ;
        RECT 2744.430 38.800 2744.750 38.860 ;
      LAYER via ;
        RECT 2278.940 1688.140 2279.200 1688.400 ;
        RECT 2283.080 1688.140 2283.340 1688.400 ;
        RECT 2283.080 38.800 2283.340 39.060 ;
        RECT 2744.460 38.800 2744.720 39.060 ;
      LAYER met2 ;
        RECT 2278.865 1700.000 2279.145 1704.000 ;
        RECT 2279.000 1688.430 2279.140 1700.000 ;
        RECT 2278.940 1688.110 2279.200 1688.430 ;
        RECT 2283.080 1688.110 2283.340 1688.430 ;
        RECT 2283.140 39.090 2283.280 1688.110 ;
        RECT 2283.080 38.770 2283.340 39.090 ;
        RECT 2744.460 38.770 2744.720 39.090 ;
        RECT 2744.520 2.400 2744.660 38.770 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2286.270 1683.920 2286.590 1683.980 ;
        RECT 2289.950 1683.920 2290.270 1683.980 ;
        RECT 2286.270 1683.780 2290.270 1683.920 ;
        RECT 2286.270 1683.720 2286.590 1683.780 ;
        RECT 2289.950 1683.720 2290.270 1683.780 ;
        RECT 2289.950 38.660 2290.270 38.720 ;
        RECT 2761.910 38.660 2762.230 38.720 ;
        RECT 2289.950 38.520 2762.230 38.660 ;
        RECT 2289.950 38.460 2290.270 38.520 ;
        RECT 2761.910 38.460 2762.230 38.520 ;
      LAYER via ;
        RECT 2286.300 1683.720 2286.560 1683.980 ;
        RECT 2289.980 1683.720 2290.240 1683.980 ;
        RECT 2289.980 38.460 2290.240 38.720 ;
        RECT 2761.940 38.460 2762.200 38.720 ;
      LAYER met2 ;
        RECT 2286.225 1700.000 2286.505 1704.000 ;
        RECT 2286.360 1684.010 2286.500 1700.000 ;
        RECT 2286.300 1683.690 2286.560 1684.010 ;
        RECT 2289.980 1683.690 2290.240 1684.010 ;
        RECT 2290.040 38.750 2290.180 1683.690 ;
        RECT 2289.980 38.430 2290.240 38.750 ;
        RECT 2761.940 38.430 2762.200 38.750 ;
        RECT 2762.000 2.400 2762.140 38.430 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 835.430 33.900 835.750 33.960 ;
        RECT 1491.850 33.900 1492.170 33.960 ;
        RECT 835.430 33.760 1492.170 33.900 ;
        RECT 835.430 33.700 835.750 33.760 ;
        RECT 1491.850 33.700 1492.170 33.760 ;
      LAYER via ;
        RECT 835.460 33.700 835.720 33.960 ;
        RECT 1491.880 33.700 1492.140 33.960 ;
      LAYER met2 ;
        RECT 1492.725 1700.410 1493.005 1704.000 ;
        RECT 1491.940 1700.270 1493.005 1700.410 ;
        RECT 1491.940 33.990 1492.080 1700.270 ;
        RECT 1492.725 1700.000 1493.005 1700.270 ;
        RECT 835.460 33.670 835.720 33.990 ;
        RECT 1491.880 33.670 1492.140 33.990 ;
        RECT 835.520 2.400 835.660 33.670 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2293.630 1689.360 2293.950 1689.420 ;
        RECT 2296.850 1689.360 2297.170 1689.420 ;
        RECT 2293.630 1689.220 2297.170 1689.360 ;
        RECT 2293.630 1689.160 2293.950 1689.220 ;
        RECT 2296.850 1689.160 2297.170 1689.220 ;
        RECT 2296.850 38.320 2297.170 38.380 ;
        RECT 2779.850 38.320 2780.170 38.380 ;
        RECT 2296.850 38.180 2780.170 38.320 ;
        RECT 2296.850 38.120 2297.170 38.180 ;
        RECT 2779.850 38.120 2780.170 38.180 ;
      LAYER via ;
        RECT 2293.660 1689.160 2293.920 1689.420 ;
        RECT 2296.880 1689.160 2297.140 1689.420 ;
        RECT 2296.880 38.120 2297.140 38.380 ;
        RECT 2779.880 38.120 2780.140 38.380 ;
      LAYER met2 ;
        RECT 2293.585 1700.000 2293.865 1704.000 ;
        RECT 2293.720 1689.450 2293.860 1700.000 ;
        RECT 2293.660 1689.130 2293.920 1689.450 ;
        RECT 2296.880 1689.130 2297.140 1689.450 ;
        RECT 2296.940 38.410 2297.080 1689.130 ;
        RECT 2296.880 38.090 2297.140 38.410 ;
        RECT 2779.880 38.090 2780.140 38.410 ;
        RECT 2779.940 2.400 2780.080 38.090 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2300.990 1684.260 2301.310 1684.320 ;
        RECT 2303.750 1684.260 2304.070 1684.320 ;
        RECT 2300.990 1684.120 2304.070 1684.260 ;
        RECT 2300.990 1684.060 2301.310 1684.120 ;
        RECT 2303.750 1684.060 2304.070 1684.120 ;
        RECT 2303.750 37.980 2304.070 38.040 ;
        RECT 2797.790 37.980 2798.110 38.040 ;
        RECT 2303.750 37.840 2798.110 37.980 ;
        RECT 2303.750 37.780 2304.070 37.840 ;
        RECT 2797.790 37.780 2798.110 37.840 ;
      LAYER via ;
        RECT 2301.020 1684.060 2301.280 1684.320 ;
        RECT 2303.780 1684.060 2304.040 1684.320 ;
        RECT 2303.780 37.780 2304.040 38.040 ;
        RECT 2797.820 37.780 2798.080 38.040 ;
      LAYER met2 ;
        RECT 2300.945 1700.000 2301.225 1704.000 ;
        RECT 2301.080 1684.350 2301.220 1700.000 ;
        RECT 2301.020 1684.030 2301.280 1684.350 ;
        RECT 2303.780 1684.030 2304.040 1684.350 ;
        RECT 2303.840 38.070 2303.980 1684.030 ;
        RECT 2303.780 37.750 2304.040 38.070 ;
        RECT 2797.820 37.750 2798.080 38.070 ;
        RECT 2797.880 2.400 2798.020 37.750 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2324.985 1684.445 2326.075 1684.615 ;
        RECT 2325.905 1683.425 2326.075 1684.445 ;
      LAYER met1 ;
        RECT 2308.350 1684.600 2308.670 1684.660 ;
        RECT 2324.925 1684.600 2325.215 1684.645 ;
        RECT 2308.350 1684.460 2325.215 1684.600 ;
        RECT 2308.350 1684.400 2308.670 1684.460 ;
        RECT 2324.925 1684.415 2325.215 1684.460 ;
        RECT 2528.690 1683.920 2529.010 1683.980 ;
        RECT 2347.080 1683.780 2529.010 1683.920 ;
        RECT 2325.845 1683.580 2326.135 1683.625 ;
        RECT 2347.080 1683.580 2347.220 1683.780 ;
        RECT 2528.690 1683.720 2529.010 1683.780 ;
        RECT 2325.845 1683.440 2347.220 1683.580 ;
        RECT 2325.845 1683.395 2326.135 1683.440 ;
        RECT 2528.690 15.880 2529.010 15.940 ;
        RECT 2815.730 15.880 2816.050 15.940 ;
        RECT 2528.690 15.740 2816.050 15.880 ;
        RECT 2528.690 15.680 2529.010 15.740 ;
        RECT 2815.730 15.680 2816.050 15.740 ;
      LAYER via ;
        RECT 2308.380 1684.400 2308.640 1684.660 ;
        RECT 2528.720 1683.720 2528.980 1683.980 ;
        RECT 2528.720 15.680 2528.980 15.940 ;
        RECT 2815.760 15.680 2816.020 15.940 ;
      LAYER met2 ;
        RECT 2308.305 1700.000 2308.585 1704.000 ;
        RECT 2308.440 1684.690 2308.580 1700.000 ;
        RECT 2308.380 1684.370 2308.640 1684.690 ;
        RECT 2528.720 1683.690 2528.980 1684.010 ;
        RECT 2528.780 15.970 2528.920 1683.690 ;
        RECT 2528.720 15.650 2528.980 15.970 ;
        RECT 2815.760 15.650 2816.020 15.970 ;
        RECT 2815.820 2.400 2815.960 15.650 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2318.010 18.260 2318.330 18.320 ;
        RECT 2833.670 18.260 2833.990 18.320 ;
        RECT 2318.010 18.120 2833.990 18.260 ;
        RECT 2318.010 18.060 2318.330 18.120 ;
        RECT 2833.670 18.060 2833.990 18.120 ;
      LAYER via ;
        RECT 2318.040 18.060 2318.300 18.320 ;
        RECT 2833.700 18.060 2833.960 18.320 ;
      LAYER met2 ;
        RECT 2315.665 1700.410 2315.945 1704.000 ;
        RECT 2315.665 1700.270 2317.320 1700.410 ;
        RECT 2315.665 1700.000 2315.945 1700.270 ;
        RECT 2317.180 1684.600 2317.320 1700.270 ;
        RECT 2317.180 1684.460 2318.240 1684.600 ;
        RECT 2318.100 18.350 2318.240 1684.460 ;
        RECT 2318.040 18.030 2318.300 18.350 ;
        RECT 2833.700 18.030 2833.960 18.350 ;
        RECT 2833.760 2.400 2833.900 18.030 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2590.865 15.045 2591.035 16.235 ;
      LAYER mcon ;
        RECT 2590.865 16.065 2591.035 16.235 ;
      LAYER met1 ;
        RECT 2549.390 1684.260 2549.710 1684.320 ;
        RECT 2346.620 1684.120 2549.710 1684.260 ;
        RECT 2346.620 1683.920 2346.760 1684.120 ;
        RECT 2549.390 1684.060 2549.710 1684.120 ;
        RECT 2325.460 1683.780 2346.760 1683.920 ;
        RECT 2324.450 1683.580 2324.770 1683.640 ;
        RECT 2325.460 1683.580 2325.600 1683.780 ;
        RECT 2324.450 1683.440 2325.600 1683.580 ;
        RECT 2324.450 1683.380 2324.770 1683.440 ;
        RECT 2590.805 16.220 2591.095 16.265 ;
        RECT 2851.150 16.220 2851.470 16.280 ;
        RECT 2590.805 16.080 2851.470 16.220 ;
        RECT 2590.805 16.035 2591.095 16.080 ;
        RECT 2851.150 16.020 2851.470 16.080 ;
        RECT 2549.390 15.200 2549.710 15.260 ;
        RECT 2590.805 15.200 2591.095 15.245 ;
        RECT 2549.390 15.060 2591.095 15.200 ;
        RECT 2549.390 15.000 2549.710 15.060 ;
        RECT 2590.805 15.015 2591.095 15.060 ;
      LAYER via ;
        RECT 2549.420 1684.060 2549.680 1684.320 ;
        RECT 2324.480 1683.380 2324.740 1683.640 ;
        RECT 2851.180 16.020 2851.440 16.280 ;
        RECT 2549.420 15.000 2549.680 15.260 ;
      LAYER met2 ;
        RECT 2323.025 1700.410 2323.305 1704.000 ;
        RECT 2323.025 1700.270 2324.680 1700.410 ;
        RECT 2323.025 1700.000 2323.305 1700.270 ;
        RECT 2324.540 1683.670 2324.680 1700.270 ;
        RECT 2549.420 1684.030 2549.680 1684.350 ;
        RECT 2324.480 1683.350 2324.740 1683.670 ;
        RECT 2549.480 15.290 2549.620 1684.030 ;
        RECT 2851.180 15.990 2851.440 16.310 ;
        RECT 2549.420 14.970 2549.680 15.290 ;
        RECT 2851.240 2.400 2851.380 15.990 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2331.350 17.580 2331.670 17.640 ;
        RECT 2869.090 17.580 2869.410 17.640 ;
        RECT 2331.350 17.440 2869.410 17.580 ;
        RECT 2331.350 17.380 2331.670 17.440 ;
        RECT 2869.090 17.380 2869.410 17.440 ;
      LAYER via ;
        RECT 2331.380 17.380 2331.640 17.640 ;
        RECT 2869.120 17.380 2869.380 17.640 ;
      LAYER met2 ;
        RECT 2330.385 1700.410 2330.665 1704.000 ;
        RECT 2330.385 1700.270 2331.580 1700.410 ;
        RECT 2330.385 1700.000 2330.665 1700.270 ;
        RECT 2331.440 17.670 2331.580 1700.270 ;
        RECT 2331.380 17.350 2331.640 17.670 ;
        RECT 2869.120 17.350 2869.380 17.670 ;
        RECT 2869.180 2.400 2869.320 17.350 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2887.030 16.560 2887.350 16.620 ;
        RECT 2590.420 16.420 2887.350 16.560 ;
        RECT 2563.190 16.220 2563.510 16.280 ;
        RECT 2590.420 16.220 2590.560 16.420 ;
        RECT 2887.030 16.360 2887.350 16.420 ;
        RECT 2563.190 16.080 2590.560 16.220 ;
        RECT 2563.190 16.020 2563.510 16.080 ;
      LAYER via ;
        RECT 2563.220 16.020 2563.480 16.280 ;
        RECT 2887.060 16.360 2887.320 16.620 ;
      LAYER met2 ;
        RECT 2337.745 1700.000 2338.025 1704.000 ;
        RECT 2337.880 1686.925 2338.020 1700.000 ;
        RECT 2337.810 1686.555 2338.090 1686.925 ;
        RECT 2563.210 1686.555 2563.490 1686.925 ;
        RECT 2563.280 16.310 2563.420 1686.555 ;
        RECT 2887.060 16.330 2887.320 16.650 ;
        RECT 2563.220 15.990 2563.480 16.310 ;
        RECT 2887.120 2.400 2887.260 16.330 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
      LAYER via2 ;
        RECT 2337.810 1686.600 2338.090 1686.880 ;
        RECT 2563.210 1686.600 2563.490 1686.880 ;
      LAYER met3 ;
        RECT 2337.785 1686.890 2338.115 1686.905 ;
        RECT 2563.185 1686.890 2563.515 1686.905 ;
        RECT 2337.785 1686.590 2563.515 1686.890 ;
        RECT 2337.785 1686.575 2338.115 1686.590 ;
        RECT 2563.185 1686.575 2563.515 1686.590 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2344.230 58.720 2344.550 58.780 ;
        RECT 2345.610 58.720 2345.930 58.780 ;
        RECT 2344.230 58.580 2345.930 58.720 ;
        RECT 2344.230 58.520 2344.550 58.580 ;
        RECT 2345.610 58.520 2345.930 58.580 ;
      LAYER via ;
        RECT 2344.260 58.520 2344.520 58.780 ;
        RECT 2345.640 58.520 2345.900 58.780 ;
      LAYER met2 ;
        RECT 2345.105 1700.410 2345.385 1704.000 ;
        RECT 2345.105 1700.270 2345.840 1700.410 ;
        RECT 2345.105 1700.000 2345.385 1700.270 ;
        RECT 2345.700 58.810 2345.840 1700.270 ;
        RECT 2344.260 58.490 2344.520 58.810 ;
        RECT 2345.640 58.490 2345.900 58.810 ;
        RECT 2344.320 16.845 2344.460 58.490 ;
        RECT 2344.250 16.475 2344.530 16.845 ;
        RECT 2904.990 16.475 2905.270 16.845 ;
        RECT 2905.060 2.400 2905.200 16.475 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
      LAYER via2 ;
        RECT 2344.250 16.520 2344.530 16.800 ;
        RECT 2904.990 16.520 2905.270 16.800 ;
      LAYER met3 ;
        RECT 2344.225 16.810 2344.555 16.825 ;
        RECT 2904.965 16.810 2905.295 16.825 ;
        RECT 2344.225 16.510 2905.295 16.810 ;
        RECT 2344.225 16.495 2344.555 16.510 ;
        RECT 2904.965 16.495 2905.295 16.510 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1497.445 1159.145 1497.615 1207.255 ;
      LAYER mcon ;
        RECT 1497.445 1207.085 1497.615 1207.255 ;
      LAYER met1 ;
        RECT 1497.370 1655.360 1497.690 1655.420 ;
        RECT 1498.290 1655.360 1498.610 1655.420 ;
        RECT 1497.370 1655.220 1498.610 1655.360 ;
        RECT 1497.370 1655.160 1497.690 1655.220 ;
        RECT 1498.290 1655.160 1498.610 1655.220 ;
        RECT 1497.370 1207.240 1497.690 1207.300 ;
        RECT 1497.370 1207.100 1497.885 1207.240 ;
        RECT 1497.370 1207.040 1497.690 1207.100 ;
        RECT 1497.370 1159.300 1497.690 1159.360 ;
        RECT 1497.370 1159.160 1497.885 1159.300 ;
        RECT 1497.370 1159.100 1497.690 1159.160 ;
        RECT 852.910 34.240 853.230 34.300 ;
        RECT 1497.370 34.240 1497.690 34.300 ;
        RECT 852.910 34.100 1497.690 34.240 ;
        RECT 852.910 34.040 853.230 34.100 ;
        RECT 1497.370 34.040 1497.690 34.100 ;
      LAYER via ;
        RECT 1497.400 1655.160 1497.660 1655.420 ;
        RECT 1498.320 1655.160 1498.580 1655.420 ;
        RECT 1497.400 1207.040 1497.660 1207.300 ;
        RECT 1497.400 1159.100 1497.660 1159.360 ;
        RECT 852.940 34.040 853.200 34.300 ;
        RECT 1497.400 34.040 1497.660 34.300 ;
      LAYER met2 ;
        RECT 1500.085 1700.410 1500.365 1704.000 ;
        RECT 1498.840 1700.270 1500.365 1700.410 ;
        RECT 1498.840 1656.210 1498.980 1700.270 ;
        RECT 1500.085 1700.000 1500.365 1700.270 ;
        RECT 1498.380 1656.070 1498.980 1656.210 ;
        RECT 1498.380 1655.450 1498.520 1656.070 ;
        RECT 1497.400 1655.130 1497.660 1655.450 ;
        RECT 1498.320 1655.130 1498.580 1655.450 ;
        RECT 1497.460 1207.330 1497.600 1655.130 ;
        RECT 1497.400 1207.010 1497.660 1207.330 ;
        RECT 1497.400 1159.070 1497.660 1159.390 ;
        RECT 1497.460 34.330 1497.600 1159.070 ;
        RECT 852.940 34.010 853.200 34.330 ;
        RECT 1497.400 34.010 1497.660 34.330 ;
        RECT 853.000 2.400 853.140 34.010 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1504.270 1678.140 1504.590 1678.200 ;
        RECT 1506.110 1678.140 1506.430 1678.200 ;
        RECT 1504.270 1678.000 1506.430 1678.140 ;
        RECT 1504.270 1677.940 1504.590 1678.000 ;
        RECT 1506.110 1677.940 1506.430 1678.000 ;
        RECT 870.850 30.500 871.170 30.560 ;
        RECT 1504.270 30.500 1504.590 30.560 ;
        RECT 870.850 30.360 1504.590 30.500 ;
        RECT 870.850 30.300 871.170 30.360 ;
        RECT 1504.270 30.300 1504.590 30.360 ;
      LAYER via ;
        RECT 1504.300 1677.940 1504.560 1678.200 ;
        RECT 1506.140 1677.940 1506.400 1678.200 ;
        RECT 870.880 30.300 871.140 30.560 ;
        RECT 1504.300 30.300 1504.560 30.560 ;
      LAYER met2 ;
        RECT 1507.445 1700.410 1507.725 1704.000 ;
        RECT 1506.200 1700.270 1507.725 1700.410 ;
        RECT 1506.200 1678.230 1506.340 1700.270 ;
        RECT 1507.445 1700.000 1507.725 1700.270 ;
        RECT 1504.300 1677.910 1504.560 1678.230 ;
        RECT 1506.140 1677.910 1506.400 1678.230 ;
        RECT 1504.360 30.590 1504.500 1677.910 ;
        RECT 870.880 30.270 871.140 30.590 ;
        RECT 1504.300 30.270 1504.560 30.590 ;
        RECT 870.940 2.400 871.080 30.270 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1511.170 1678.480 1511.490 1678.540 ;
        RECT 1513.470 1678.480 1513.790 1678.540 ;
        RECT 1511.170 1678.340 1513.790 1678.480 ;
        RECT 1511.170 1678.280 1511.490 1678.340 ;
        RECT 1513.470 1678.280 1513.790 1678.340 ;
        RECT 888.790 30.160 889.110 30.220 ;
        RECT 1511.170 30.160 1511.490 30.220 ;
        RECT 888.790 30.020 1511.490 30.160 ;
        RECT 888.790 29.960 889.110 30.020 ;
        RECT 1511.170 29.960 1511.490 30.020 ;
      LAYER via ;
        RECT 1511.200 1678.280 1511.460 1678.540 ;
        RECT 1513.500 1678.280 1513.760 1678.540 ;
        RECT 888.820 29.960 889.080 30.220 ;
        RECT 1511.200 29.960 1511.460 30.220 ;
      LAYER met2 ;
        RECT 1514.805 1700.410 1515.085 1704.000 ;
        RECT 1513.560 1700.270 1515.085 1700.410 ;
        RECT 1513.560 1678.570 1513.700 1700.270 ;
        RECT 1514.805 1700.000 1515.085 1700.270 ;
        RECT 1511.200 1678.250 1511.460 1678.570 ;
        RECT 1513.500 1678.250 1513.760 1678.570 ;
        RECT 1511.260 30.250 1511.400 1678.250 ;
        RECT 888.820 29.930 889.080 30.250 ;
        RECT 1511.200 29.930 1511.460 30.250 ;
        RECT 888.880 2.400 889.020 29.930 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1518.070 1678.140 1518.390 1678.200 ;
        RECT 1520.830 1678.140 1521.150 1678.200 ;
        RECT 1518.070 1678.000 1521.150 1678.140 ;
        RECT 1518.070 1677.940 1518.390 1678.000 ;
        RECT 1520.830 1677.940 1521.150 1678.000 ;
        RECT 906.730 29.820 907.050 29.880 ;
        RECT 1518.070 29.820 1518.390 29.880 ;
        RECT 906.730 29.680 1518.390 29.820 ;
        RECT 906.730 29.620 907.050 29.680 ;
        RECT 1518.070 29.620 1518.390 29.680 ;
      LAYER via ;
        RECT 1518.100 1677.940 1518.360 1678.200 ;
        RECT 1520.860 1677.940 1521.120 1678.200 ;
        RECT 906.760 29.620 907.020 29.880 ;
        RECT 1518.100 29.620 1518.360 29.880 ;
      LAYER met2 ;
        RECT 1522.165 1700.410 1522.445 1704.000 ;
        RECT 1520.920 1700.270 1522.445 1700.410 ;
        RECT 1520.920 1678.230 1521.060 1700.270 ;
        RECT 1522.165 1700.000 1522.445 1700.270 ;
        RECT 1518.100 1677.910 1518.360 1678.230 ;
        RECT 1520.860 1677.910 1521.120 1678.230 ;
        RECT 1518.160 29.910 1518.300 1677.910 ;
        RECT 906.760 29.590 907.020 29.910 ;
        RECT 1518.100 29.590 1518.360 29.910 ;
        RECT 906.820 2.400 906.960 29.590 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1524.970 1678.140 1525.290 1678.200 ;
        RECT 1528.190 1678.140 1528.510 1678.200 ;
        RECT 1524.970 1678.000 1528.510 1678.140 ;
        RECT 1524.970 1677.940 1525.290 1678.000 ;
        RECT 1528.190 1677.940 1528.510 1678.000 ;
        RECT 924.210 29.480 924.530 29.540 ;
        RECT 1524.970 29.480 1525.290 29.540 ;
        RECT 924.210 29.340 1525.290 29.480 ;
        RECT 924.210 29.280 924.530 29.340 ;
        RECT 1524.970 29.280 1525.290 29.340 ;
      LAYER via ;
        RECT 1525.000 1677.940 1525.260 1678.200 ;
        RECT 1528.220 1677.940 1528.480 1678.200 ;
        RECT 924.240 29.280 924.500 29.540 ;
        RECT 1525.000 29.280 1525.260 29.540 ;
      LAYER met2 ;
        RECT 1529.525 1700.410 1529.805 1704.000 ;
        RECT 1528.280 1700.270 1529.805 1700.410 ;
        RECT 1528.280 1678.230 1528.420 1700.270 ;
        RECT 1529.525 1700.000 1529.805 1700.270 ;
        RECT 1525.000 1677.910 1525.260 1678.230 ;
        RECT 1528.220 1677.910 1528.480 1678.230 ;
        RECT 1525.060 29.570 1525.200 1677.910 ;
        RECT 924.240 29.250 924.500 29.570 ;
        RECT 1525.000 29.250 1525.260 29.570 ;
        RECT 924.300 2.400 924.440 29.250 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1534.245 1497.445 1534.415 1587.035 ;
        RECT 1533.785 1200.285 1533.955 1241.935 ;
        RECT 1534.245 855.525 1534.415 903.975 ;
        RECT 1534.705 179.605 1534.875 203.915 ;
        RECT 1533.325 131.665 1533.495 155.635 ;
      LAYER mcon ;
        RECT 1534.245 1586.865 1534.415 1587.035 ;
        RECT 1533.785 1241.765 1533.955 1241.935 ;
        RECT 1534.245 903.805 1534.415 903.975 ;
        RECT 1534.705 203.745 1534.875 203.915 ;
        RECT 1533.325 155.465 1533.495 155.635 ;
      LAYER met1 ;
        RECT 1533.710 1594.160 1534.030 1594.220 ;
        RECT 1534.170 1594.160 1534.490 1594.220 ;
        RECT 1533.710 1594.020 1534.490 1594.160 ;
        RECT 1533.710 1593.960 1534.030 1594.020 ;
        RECT 1534.170 1593.960 1534.490 1594.020 ;
        RECT 1534.170 1587.020 1534.490 1587.080 ;
        RECT 1533.975 1586.880 1534.490 1587.020 ;
        RECT 1534.170 1586.820 1534.490 1586.880 ;
        RECT 1534.170 1497.600 1534.490 1497.660 ;
        RECT 1533.975 1497.460 1534.490 1497.600 ;
        RECT 1534.170 1497.400 1534.490 1497.460 ;
        RECT 1534.170 1463.060 1534.490 1463.320 ;
        RECT 1534.260 1462.640 1534.400 1463.060 ;
        RECT 1534.170 1462.380 1534.490 1462.640 ;
        RECT 1533.710 1249.060 1534.030 1249.120 ;
        RECT 1534.630 1249.060 1534.950 1249.120 ;
        RECT 1533.710 1248.920 1534.950 1249.060 ;
        RECT 1533.710 1248.860 1534.030 1248.920 ;
        RECT 1534.630 1248.860 1534.950 1248.920 ;
        RECT 1533.710 1241.920 1534.030 1241.980 ;
        RECT 1533.515 1241.780 1534.030 1241.920 ;
        RECT 1533.710 1241.720 1534.030 1241.780 ;
        RECT 1533.725 1200.440 1534.015 1200.485 ;
        RECT 1534.170 1200.440 1534.490 1200.500 ;
        RECT 1533.725 1200.300 1534.490 1200.440 ;
        RECT 1533.725 1200.255 1534.015 1200.300 ;
        RECT 1534.170 1200.240 1534.490 1200.300 ;
        RECT 1534.630 1159.640 1534.950 1159.700 ;
        RECT 1534.260 1159.500 1534.950 1159.640 ;
        RECT 1534.260 1159.020 1534.400 1159.500 ;
        RECT 1534.630 1159.440 1534.950 1159.500 ;
        RECT 1534.170 1158.760 1534.490 1159.020 ;
        RECT 1533.710 1068.520 1534.030 1068.580 ;
        RECT 1534.630 1068.520 1534.950 1068.580 ;
        RECT 1533.710 1068.380 1534.950 1068.520 ;
        RECT 1533.710 1068.320 1534.030 1068.380 ;
        RECT 1534.630 1068.320 1534.950 1068.380 ;
        RECT 1533.710 1014.460 1534.030 1014.520 ;
        RECT 1534.170 1014.460 1534.490 1014.520 ;
        RECT 1533.710 1014.320 1534.490 1014.460 ;
        RECT 1533.710 1014.260 1534.030 1014.320 ;
        RECT 1534.170 1014.260 1534.490 1014.320 ;
        RECT 1534.170 1007.320 1534.490 1007.380 ;
        RECT 1534.630 1007.320 1534.950 1007.380 ;
        RECT 1534.170 1007.180 1534.950 1007.320 ;
        RECT 1534.170 1007.120 1534.490 1007.180 ;
        RECT 1534.630 1007.120 1534.950 1007.180 ;
        RECT 1534.170 917.900 1534.490 917.960 ;
        RECT 1534.630 917.900 1534.950 917.960 ;
        RECT 1534.170 917.760 1534.950 917.900 ;
        RECT 1534.170 917.700 1534.490 917.760 ;
        RECT 1534.630 917.700 1534.950 917.760 ;
        RECT 1534.170 903.960 1534.490 904.020 ;
        RECT 1533.975 903.820 1534.490 903.960 ;
        RECT 1534.170 903.760 1534.490 903.820 ;
        RECT 1534.170 855.680 1534.490 855.740 ;
        RECT 1533.975 855.540 1534.490 855.680 ;
        RECT 1534.170 855.480 1534.490 855.540 ;
        RECT 1533.710 641.620 1534.030 641.880 ;
        RECT 1533.800 641.480 1533.940 641.620 ;
        RECT 1534.170 641.480 1534.490 641.540 ;
        RECT 1533.800 641.340 1534.490 641.480 ;
        RECT 1534.170 641.280 1534.490 641.340 ;
        RECT 1534.170 427.960 1534.490 428.020 ;
        RECT 1534.630 427.960 1534.950 428.020 ;
        RECT 1534.170 427.820 1534.950 427.960 ;
        RECT 1534.170 427.760 1534.490 427.820 ;
        RECT 1534.630 427.760 1534.950 427.820 ;
        RECT 1533.710 386.480 1534.030 386.540 ;
        RECT 1534.170 386.480 1534.490 386.540 ;
        RECT 1533.710 386.340 1534.490 386.480 ;
        RECT 1533.710 386.280 1534.030 386.340 ;
        RECT 1534.170 386.280 1534.490 386.340 ;
        RECT 1533.710 331.060 1534.030 331.120 ;
        RECT 1534.630 331.060 1534.950 331.120 ;
        RECT 1533.710 330.920 1534.950 331.060 ;
        RECT 1533.710 330.860 1534.030 330.920 ;
        RECT 1534.630 330.860 1534.950 330.920 ;
        RECT 1534.630 203.900 1534.950 203.960 ;
        RECT 1534.435 203.760 1534.950 203.900 ;
        RECT 1534.630 203.700 1534.950 203.760 ;
        RECT 1533.710 179.760 1534.030 179.820 ;
        RECT 1534.645 179.760 1534.935 179.805 ;
        RECT 1533.710 179.620 1534.935 179.760 ;
        RECT 1533.710 179.560 1534.030 179.620 ;
        RECT 1534.645 179.575 1534.935 179.620 ;
        RECT 1533.265 155.620 1533.555 155.665 ;
        RECT 1533.710 155.620 1534.030 155.680 ;
        RECT 1533.265 155.480 1534.030 155.620 ;
        RECT 1533.265 155.435 1533.555 155.480 ;
        RECT 1533.710 155.420 1534.030 155.480 ;
        RECT 1533.250 131.820 1533.570 131.880 ;
        RECT 1533.055 131.680 1533.570 131.820 ;
        RECT 1533.250 131.620 1533.570 131.680 ;
        RECT 1534.170 76.060 1534.490 76.120 ;
        RECT 1535.090 76.060 1535.410 76.120 ;
        RECT 1534.170 75.920 1535.410 76.060 ;
        RECT 1534.170 75.860 1534.490 75.920 ;
        RECT 1535.090 75.860 1535.410 75.920 ;
        RECT 1533.250 34.580 1533.570 34.640 ;
        RECT 1534.170 34.580 1534.490 34.640 ;
        RECT 1533.250 34.440 1534.490 34.580 ;
        RECT 1533.250 34.380 1533.570 34.440 ;
        RECT 1534.170 34.380 1534.490 34.440 ;
        RECT 942.150 29.140 942.470 29.200 ;
        RECT 1533.250 29.140 1533.570 29.200 ;
        RECT 942.150 29.000 1533.570 29.140 ;
        RECT 942.150 28.940 942.470 29.000 ;
        RECT 1533.250 28.940 1533.570 29.000 ;
      LAYER via ;
        RECT 1533.740 1593.960 1534.000 1594.220 ;
        RECT 1534.200 1593.960 1534.460 1594.220 ;
        RECT 1534.200 1586.820 1534.460 1587.080 ;
        RECT 1534.200 1497.400 1534.460 1497.660 ;
        RECT 1534.200 1463.060 1534.460 1463.320 ;
        RECT 1534.200 1462.380 1534.460 1462.640 ;
        RECT 1533.740 1248.860 1534.000 1249.120 ;
        RECT 1534.660 1248.860 1534.920 1249.120 ;
        RECT 1533.740 1241.720 1534.000 1241.980 ;
        RECT 1534.200 1200.240 1534.460 1200.500 ;
        RECT 1534.660 1159.440 1534.920 1159.700 ;
        RECT 1534.200 1158.760 1534.460 1159.020 ;
        RECT 1533.740 1068.320 1534.000 1068.580 ;
        RECT 1534.660 1068.320 1534.920 1068.580 ;
        RECT 1533.740 1014.260 1534.000 1014.520 ;
        RECT 1534.200 1014.260 1534.460 1014.520 ;
        RECT 1534.200 1007.120 1534.460 1007.380 ;
        RECT 1534.660 1007.120 1534.920 1007.380 ;
        RECT 1534.200 917.700 1534.460 917.960 ;
        RECT 1534.660 917.700 1534.920 917.960 ;
        RECT 1534.200 903.760 1534.460 904.020 ;
        RECT 1534.200 855.480 1534.460 855.740 ;
        RECT 1533.740 641.620 1534.000 641.880 ;
        RECT 1534.200 641.280 1534.460 641.540 ;
        RECT 1534.200 427.760 1534.460 428.020 ;
        RECT 1534.660 427.760 1534.920 428.020 ;
        RECT 1533.740 386.280 1534.000 386.540 ;
        RECT 1534.200 386.280 1534.460 386.540 ;
        RECT 1533.740 330.860 1534.000 331.120 ;
        RECT 1534.660 330.860 1534.920 331.120 ;
        RECT 1534.660 203.700 1534.920 203.960 ;
        RECT 1533.740 179.560 1534.000 179.820 ;
        RECT 1533.740 155.420 1534.000 155.680 ;
        RECT 1533.280 131.620 1533.540 131.880 ;
        RECT 1534.200 75.860 1534.460 76.120 ;
        RECT 1535.120 75.860 1535.380 76.120 ;
        RECT 1533.280 34.380 1533.540 34.640 ;
        RECT 1534.200 34.380 1534.460 34.640 ;
        RECT 942.180 28.940 942.440 29.200 ;
        RECT 1533.280 28.940 1533.540 29.200 ;
      LAYER met2 ;
        RECT 1536.885 1700.410 1537.165 1704.000 ;
        RECT 1535.180 1700.270 1537.165 1700.410 ;
        RECT 1535.180 1656.210 1535.320 1700.270 ;
        RECT 1536.885 1700.000 1537.165 1700.270 ;
        RECT 1533.800 1656.070 1535.320 1656.210 ;
        RECT 1533.800 1594.250 1533.940 1656.070 ;
        RECT 1533.740 1593.930 1534.000 1594.250 ;
        RECT 1534.200 1593.930 1534.460 1594.250 ;
        RECT 1534.260 1587.110 1534.400 1593.930 ;
        RECT 1534.200 1586.790 1534.460 1587.110 ;
        RECT 1534.200 1497.370 1534.460 1497.690 ;
        RECT 1534.260 1463.350 1534.400 1497.370 ;
        RECT 1534.200 1463.030 1534.460 1463.350 ;
        RECT 1534.200 1462.350 1534.460 1462.670 ;
        RECT 1534.260 1376.730 1534.400 1462.350 ;
        RECT 1533.800 1376.590 1534.400 1376.730 ;
        RECT 1533.800 1322.330 1533.940 1376.590 ;
        RECT 1533.800 1322.190 1534.860 1322.330 ;
        RECT 1534.720 1317.570 1534.860 1322.190 ;
        RECT 1534.260 1317.430 1534.860 1317.570 ;
        RECT 1534.260 1273.370 1534.400 1317.430 ;
        RECT 1534.260 1273.230 1534.860 1273.370 ;
        RECT 1534.720 1249.150 1534.860 1273.230 ;
        RECT 1533.740 1248.830 1534.000 1249.150 ;
        RECT 1534.660 1248.830 1534.920 1249.150 ;
        RECT 1533.800 1242.010 1533.940 1248.830 ;
        RECT 1533.740 1241.690 1534.000 1242.010 ;
        RECT 1534.200 1200.210 1534.460 1200.530 ;
        RECT 1534.260 1193.810 1534.400 1200.210 ;
        RECT 1534.260 1193.670 1534.860 1193.810 ;
        RECT 1534.720 1159.730 1534.860 1193.670 ;
        RECT 1534.660 1159.410 1534.920 1159.730 ;
        RECT 1534.200 1158.730 1534.460 1159.050 ;
        RECT 1534.260 1104.050 1534.400 1158.730 ;
        RECT 1534.260 1103.910 1534.860 1104.050 ;
        RECT 1534.720 1068.610 1534.860 1103.910 ;
        RECT 1533.740 1068.290 1534.000 1068.610 ;
        RECT 1534.660 1068.290 1534.920 1068.610 ;
        RECT 1533.800 1014.550 1533.940 1068.290 ;
        RECT 1533.740 1014.230 1534.000 1014.550 ;
        RECT 1534.200 1014.230 1534.460 1014.550 ;
        RECT 1534.260 1007.410 1534.400 1014.230 ;
        RECT 1534.200 1007.090 1534.460 1007.410 ;
        RECT 1534.660 1007.090 1534.920 1007.410 ;
        RECT 1534.720 917.990 1534.860 1007.090 ;
        RECT 1534.200 917.670 1534.460 917.990 ;
        RECT 1534.660 917.670 1534.920 917.990 ;
        RECT 1534.260 904.050 1534.400 917.670 ;
        RECT 1534.200 903.730 1534.460 904.050 ;
        RECT 1534.200 855.450 1534.460 855.770 ;
        RECT 1534.260 806.890 1534.400 855.450 ;
        RECT 1534.260 806.750 1534.860 806.890 ;
        RECT 1534.720 772.890 1534.860 806.750 ;
        RECT 1533.800 772.750 1534.860 772.890 ;
        RECT 1533.800 748.410 1533.940 772.750 ;
        RECT 1533.800 748.270 1534.400 748.410 ;
        RECT 1534.260 676.330 1534.400 748.270 ;
        RECT 1533.800 676.190 1534.400 676.330 ;
        RECT 1533.800 641.910 1533.940 676.190 ;
        RECT 1533.740 641.590 1534.000 641.910 ;
        RECT 1534.200 641.250 1534.460 641.570 ;
        RECT 1534.260 579.770 1534.400 641.250 ;
        RECT 1533.800 579.630 1534.400 579.770 ;
        RECT 1533.800 549.170 1533.940 579.630 ;
        RECT 1533.800 549.030 1534.400 549.170 ;
        RECT 1534.260 497.490 1534.400 549.030 ;
        RECT 1534.260 497.350 1534.860 497.490 ;
        RECT 1534.720 428.050 1534.860 497.350 ;
        RECT 1534.200 427.730 1534.460 428.050 ;
        RECT 1534.660 427.730 1534.920 428.050 ;
        RECT 1534.260 386.570 1534.400 427.730 ;
        RECT 1533.740 386.250 1534.000 386.570 ;
        RECT 1534.200 386.250 1534.460 386.570 ;
        RECT 1533.800 331.150 1533.940 386.250 ;
        RECT 1533.740 330.830 1534.000 331.150 ;
        RECT 1534.660 330.830 1534.920 331.150 ;
        RECT 1534.720 203.990 1534.860 330.830 ;
        RECT 1534.660 203.670 1534.920 203.990 ;
        RECT 1533.740 179.530 1534.000 179.850 ;
        RECT 1533.800 155.710 1533.940 179.530 ;
        RECT 1533.740 155.390 1534.000 155.710 ;
        RECT 1533.280 131.590 1533.540 131.910 ;
        RECT 1533.340 124.285 1533.480 131.590 ;
        RECT 1533.270 123.915 1533.550 124.285 ;
        RECT 1535.110 123.915 1535.390 124.285 ;
        RECT 1535.180 76.150 1535.320 123.915 ;
        RECT 1534.200 75.830 1534.460 76.150 ;
        RECT 1535.120 75.830 1535.380 76.150 ;
        RECT 1534.260 34.670 1534.400 75.830 ;
        RECT 1533.280 34.350 1533.540 34.670 ;
        RECT 1534.200 34.350 1534.460 34.670 ;
        RECT 1533.340 29.230 1533.480 34.350 ;
        RECT 942.180 28.910 942.440 29.230 ;
        RECT 1533.280 28.910 1533.540 29.230 ;
        RECT 942.240 2.400 942.380 28.910 ;
        RECT 942.030 -4.800 942.590 2.400 ;
      LAYER via2 ;
        RECT 1533.270 123.960 1533.550 124.240 ;
        RECT 1535.110 123.960 1535.390 124.240 ;
      LAYER met3 ;
        RECT 1533.245 124.250 1533.575 124.265 ;
        RECT 1535.085 124.250 1535.415 124.265 ;
        RECT 1533.245 123.950 1535.415 124.250 ;
        RECT 1533.245 123.935 1533.575 123.950 ;
        RECT 1535.085 123.935 1535.415 123.950 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1538.770 1678.140 1539.090 1678.200 ;
        RECT 1542.910 1678.140 1543.230 1678.200 ;
        RECT 1538.770 1678.000 1543.230 1678.140 ;
        RECT 1538.770 1677.940 1539.090 1678.000 ;
        RECT 1542.910 1677.940 1543.230 1678.000 ;
        RECT 960.090 28.800 960.410 28.860 ;
        RECT 1538.770 28.800 1539.090 28.860 ;
        RECT 960.090 28.660 1539.090 28.800 ;
        RECT 960.090 28.600 960.410 28.660 ;
        RECT 1538.770 28.600 1539.090 28.660 ;
      LAYER via ;
        RECT 1538.800 1677.940 1539.060 1678.200 ;
        RECT 1542.940 1677.940 1543.200 1678.200 ;
        RECT 960.120 28.600 960.380 28.860 ;
        RECT 1538.800 28.600 1539.060 28.860 ;
      LAYER met2 ;
        RECT 1544.245 1700.410 1544.525 1704.000 ;
        RECT 1543.000 1700.270 1544.525 1700.410 ;
        RECT 1543.000 1678.230 1543.140 1700.270 ;
        RECT 1544.245 1700.000 1544.525 1700.270 ;
        RECT 1538.800 1677.910 1539.060 1678.230 ;
        RECT 1542.940 1677.910 1543.200 1678.230 ;
        RECT 1538.860 28.890 1539.000 1677.910 ;
        RECT 960.120 28.570 960.380 28.890 ;
        RECT 1538.800 28.570 1539.060 28.890 ;
        RECT 960.180 2.400 960.320 28.570 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1545.670 1678.140 1545.990 1678.200 ;
        RECT 1550.270 1678.140 1550.590 1678.200 ;
        RECT 1545.670 1678.000 1550.590 1678.140 ;
        RECT 1545.670 1677.940 1545.990 1678.000 ;
        RECT 1550.270 1677.940 1550.590 1678.000 ;
        RECT 978.030 28.460 978.350 28.520 ;
        RECT 1545.670 28.460 1545.990 28.520 ;
        RECT 978.030 28.320 1545.990 28.460 ;
        RECT 978.030 28.260 978.350 28.320 ;
        RECT 1545.670 28.260 1545.990 28.320 ;
      LAYER via ;
        RECT 1545.700 1677.940 1545.960 1678.200 ;
        RECT 1550.300 1677.940 1550.560 1678.200 ;
        RECT 978.060 28.260 978.320 28.520 ;
        RECT 1545.700 28.260 1545.960 28.520 ;
      LAYER met2 ;
        RECT 1551.605 1700.410 1551.885 1704.000 ;
        RECT 1550.360 1700.270 1551.885 1700.410 ;
        RECT 1550.360 1678.230 1550.500 1700.270 ;
        RECT 1551.605 1700.000 1551.885 1700.270 ;
        RECT 1545.700 1677.910 1545.960 1678.230 ;
        RECT 1550.300 1677.910 1550.560 1678.230 ;
        RECT 1545.760 28.550 1545.900 1677.910 ;
        RECT 978.060 28.230 978.320 28.550 ;
        RECT 1545.700 28.230 1545.960 28.550 ;
        RECT 978.120 2.400 978.260 28.230 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1415.030 1678.140 1415.350 1678.200 ;
        RECT 1417.790 1678.140 1418.110 1678.200 ;
        RECT 1415.030 1678.000 1418.110 1678.140 ;
        RECT 1415.030 1677.940 1415.350 1678.000 ;
        RECT 1417.790 1677.940 1418.110 1678.000 ;
        RECT 656.950 33.220 657.270 33.280 ;
        RECT 1415.030 33.220 1415.350 33.280 ;
        RECT 656.950 33.080 1415.350 33.220 ;
        RECT 656.950 33.020 657.270 33.080 ;
        RECT 1415.030 33.020 1415.350 33.080 ;
      LAYER via ;
        RECT 1415.060 1677.940 1415.320 1678.200 ;
        RECT 1417.820 1677.940 1418.080 1678.200 ;
        RECT 656.980 33.020 657.240 33.280 ;
        RECT 1415.060 33.020 1415.320 33.280 ;
      LAYER met2 ;
        RECT 1419.125 1700.410 1419.405 1704.000 ;
        RECT 1417.880 1700.270 1419.405 1700.410 ;
        RECT 1417.880 1678.230 1418.020 1700.270 ;
        RECT 1419.125 1700.000 1419.405 1700.270 ;
        RECT 1415.060 1677.910 1415.320 1678.230 ;
        RECT 1417.820 1677.910 1418.080 1678.230 ;
        RECT 1415.120 33.310 1415.260 1677.910 ;
        RECT 656.980 32.990 657.240 33.310 ;
        RECT 1415.060 32.990 1415.320 33.310 ;
        RECT 657.040 2.400 657.180 32.990 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1552.570 1678.140 1552.890 1678.200 ;
        RECT 1557.630 1678.140 1557.950 1678.200 ;
        RECT 1552.570 1678.000 1557.950 1678.140 ;
        RECT 1552.570 1677.940 1552.890 1678.000 ;
        RECT 1557.630 1677.940 1557.950 1678.000 ;
        RECT 995.970 27.780 996.290 27.840 ;
        RECT 1552.570 27.780 1552.890 27.840 ;
        RECT 995.970 27.640 1552.890 27.780 ;
        RECT 995.970 27.580 996.290 27.640 ;
        RECT 1552.570 27.580 1552.890 27.640 ;
      LAYER via ;
        RECT 1552.600 1677.940 1552.860 1678.200 ;
        RECT 1557.660 1677.940 1557.920 1678.200 ;
        RECT 996.000 27.580 996.260 27.840 ;
        RECT 1552.600 27.580 1552.860 27.840 ;
      LAYER met2 ;
        RECT 1558.965 1700.410 1559.245 1704.000 ;
        RECT 1557.720 1700.270 1559.245 1700.410 ;
        RECT 1557.720 1678.230 1557.860 1700.270 ;
        RECT 1558.965 1700.000 1559.245 1700.270 ;
        RECT 1552.600 1677.910 1552.860 1678.230 ;
        RECT 1557.660 1677.910 1557.920 1678.230 ;
        RECT 1552.660 27.870 1552.800 1677.910 ;
        RECT 996.000 27.550 996.260 27.870 ;
        RECT 1552.600 27.550 1552.860 27.870 ;
        RECT 996.060 2.400 996.200 27.550 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.450 28.120 1013.770 28.180 ;
        RECT 1566.370 28.120 1566.690 28.180 ;
        RECT 1013.450 27.980 1566.690 28.120 ;
        RECT 1013.450 27.920 1013.770 27.980 ;
        RECT 1566.370 27.920 1566.690 27.980 ;
      LAYER via ;
        RECT 1013.480 27.920 1013.740 28.180 ;
        RECT 1566.400 27.920 1566.660 28.180 ;
      LAYER met2 ;
        RECT 1566.325 1700.000 1566.605 1704.000 ;
        RECT 1566.460 28.210 1566.600 1700.000 ;
        RECT 1013.480 27.890 1013.740 28.210 ;
        RECT 1566.400 27.890 1566.660 28.210 ;
        RECT 1013.540 2.400 1013.680 27.890 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1034.610 64.840 1034.930 64.900 ;
        RECT 1574.190 64.840 1574.510 64.900 ;
        RECT 1034.610 64.700 1574.510 64.840 ;
        RECT 1034.610 64.640 1034.930 64.700 ;
        RECT 1574.190 64.640 1574.510 64.700 ;
      LAYER via ;
        RECT 1034.640 64.640 1034.900 64.900 ;
        RECT 1574.220 64.640 1574.480 64.900 ;
      LAYER met2 ;
        RECT 1573.685 1700.410 1573.965 1704.000 ;
        RECT 1573.685 1700.270 1574.420 1700.410 ;
        RECT 1573.685 1700.000 1573.965 1700.270 ;
        RECT 1574.280 64.930 1574.420 1700.270 ;
        RECT 1034.640 64.610 1034.900 64.930 ;
        RECT 1574.220 64.610 1574.480 64.930 ;
        RECT 1034.700 16.730 1034.840 64.610 ;
        RECT 1031.480 16.590 1034.840 16.730 ;
        RECT 1031.480 2.400 1031.620 16.590 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1055.310 64.500 1055.630 64.560 ;
        RECT 1581.090 64.500 1581.410 64.560 ;
        RECT 1055.310 64.360 1581.410 64.500 ;
        RECT 1055.310 64.300 1055.630 64.360 ;
        RECT 1581.090 64.300 1581.410 64.360 ;
        RECT 1049.330 20.980 1049.650 21.040 ;
        RECT 1055.310 20.980 1055.630 21.040 ;
        RECT 1049.330 20.840 1055.630 20.980 ;
        RECT 1049.330 20.780 1049.650 20.840 ;
        RECT 1055.310 20.780 1055.630 20.840 ;
      LAYER via ;
        RECT 1055.340 64.300 1055.600 64.560 ;
        RECT 1581.120 64.300 1581.380 64.560 ;
        RECT 1049.360 20.780 1049.620 21.040 ;
        RECT 1055.340 20.780 1055.600 21.040 ;
      LAYER met2 ;
        RECT 1581.045 1700.000 1581.325 1704.000 ;
        RECT 1581.180 64.590 1581.320 1700.000 ;
        RECT 1055.340 64.270 1055.600 64.590 ;
        RECT 1581.120 64.270 1581.380 64.590 ;
        RECT 1055.400 21.070 1055.540 64.270 ;
        RECT 1049.360 20.750 1049.620 21.070 ;
        RECT 1055.340 20.750 1055.600 21.070 ;
        RECT 1049.420 2.400 1049.560 20.750 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1069.110 64.160 1069.430 64.220 ;
        RECT 1587.990 64.160 1588.310 64.220 ;
        RECT 1069.110 64.020 1588.310 64.160 ;
        RECT 1069.110 63.960 1069.430 64.020 ;
        RECT 1587.990 63.960 1588.310 64.020 ;
      LAYER via ;
        RECT 1069.140 63.960 1069.400 64.220 ;
        RECT 1588.020 63.960 1588.280 64.220 ;
      LAYER met2 ;
        RECT 1588.405 1700.410 1588.685 1704.000 ;
        RECT 1588.080 1700.270 1588.685 1700.410 ;
        RECT 1588.080 64.250 1588.220 1700.270 ;
        RECT 1588.405 1700.000 1588.685 1700.270 ;
        RECT 1069.140 63.930 1069.400 64.250 ;
        RECT 1588.020 63.930 1588.280 64.250 ;
        RECT 1069.200 16.730 1069.340 63.930 ;
        RECT 1067.360 16.590 1069.340 16.730 ;
        RECT 1067.360 2.400 1067.500 16.590 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1089.810 63.820 1090.130 63.880 ;
        RECT 1594.890 63.820 1595.210 63.880 ;
        RECT 1089.810 63.680 1595.210 63.820 ;
        RECT 1089.810 63.620 1090.130 63.680 ;
        RECT 1594.890 63.620 1595.210 63.680 ;
      LAYER via ;
        RECT 1089.840 63.620 1090.100 63.880 ;
        RECT 1594.920 63.620 1595.180 63.880 ;
      LAYER met2 ;
        RECT 1595.765 1700.410 1596.045 1704.000 ;
        RECT 1594.980 1700.270 1596.045 1700.410 ;
        RECT 1594.980 63.910 1595.120 1700.270 ;
        RECT 1595.765 1700.000 1596.045 1700.270 ;
        RECT 1089.840 63.590 1090.100 63.910 ;
        RECT 1594.920 63.590 1595.180 63.910 ;
        RECT 1089.900 16.730 1090.040 63.590 ;
        RECT 1085.300 16.590 1090.040 16.730 ;
        RECT 1085.300 2.400 1085.440 16.590 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1103.610 63.480 1103.930 63.540 ;
        RECT 1601.330 63.480 1601.650 63.540 ;
        RECT 1103.610 63.340 1601.650 63.480 ;
        RECT 1103.610 63.280 1103.930 63.340 ;
        RECT 1601.330 63.280 1601.650 63.340 ;
      LAYER via ;
        RECT 1103.640 63.280 1103.900 63.540 ;
        RECT 1601.360 63.280 1601.620 63.540 ;
      LAYER met2 ;
        RECT 1603.125 1700.410 1603.405 1704.000 ;
        RECT 1601.420 1700.270 1603.405 1700.410 ;
        RECT 1601.420 63.570 1601.560 1700.270 ;
        RECT 1603.125 1700.000 1603.405 1700.270 ;
        RECT 1103.640 63.250 1103.900 63.570 ;
        RECT 1601.360 63.250 1601.620 63.570 ;
        RECT 1103.700 16.730 1103.840 63.250 ;
        RECT 1102.780 16.590 1103.840 16.730 ;
        RECT 1102.780 2.400 1102.920 16.590 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1124.310 63.140 1124.630 63.200 ;
        RECT 1608.690 63.140 1609.010 63.200 ;
        RECT 1124.310 63.000 1609.010 63.140 ;
        RECT 1124.310 62.940 1124.630 63.000 ;
        RECT 1608.690 62.940 1609.010 63.000 ;
      LAYER via ;
        RECT 1124.340 62.940 1124.600 63.200 ;
        RECT 1608.720 62.940 1608.980 63.200 ;
      LAYER met2 ;
        RECT 1610.485 1700.410 1610.765 1704.000 ;
        RECT 1608.780 1700.270 1610.765 1700.410 ;
        RECT 1608.780 63.230 1608.920 1700.270 ;
        RECT 1610.485 1700.000 1610.765 1700.270 ;
        RECT 1124.340 62.910 1124.600 63.230 ;
        RECT 1608.720 62.910 1608.980 63.230 ;
        RECT 1124.400 16.730 1124.540 62.910 ;
        RECT 1120.720 16.590 1124.540 16.730 ;
        RECT 1120.720 2.400 1120.860 16.590 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.010 62.800 1145.330 62.860 ;
        RECT 1615.590 62.800 1615.910 62.860 ;
        RECT 1145.010 62.660 1615.910 62.800 ;
        RECT 1145.010 62.600 1145.330 62.660 ;
        RECT 1615.590 62.600 1615.910 62.660 ;
        RECT 1138.570 37.980 1138.890 38.040 ;
        RECT 1145.010 37.980 1145.330 38.040 ;
        RECT 1138.570 37.840 1145.330 37.980 ;
        RECT 1138.570 37.780 1138.890 37.840 ;
        RECT 1145.010 37.780 1145.330 37.840 ;
      LAYER via ;
        RECT 1145.040 62.600 1145.300 62.860 ;
        RECT 1615.620 62.600 1615.880 62.860 ;
        RECT 1138.600 37.780 1138.860 38.040 ;
        RECT 1145.040 37.780 1145.300 38.040 ;
      LAYER met2 ;
        RECT 1617.385 1700.410 1617.665 1704.000 ;
        RECT 1615.680 1700.270 1617.665 1700.410 ;
        RECT 1615.680 62.890 1615.820 1700.270 ;
        RECT 1617.385 1700.000 1617.665 1700.270 ;
        RECT 1145.040 62.570 1145.300 62.890 ;
        RECT 1615.620 62.570 1615.880 62.890 ;
        RECT 1145.100 38.070 1145.240 62.570 ;
        RECT 1138.600 37.750 1138.860 38.070 ;
        RECT 1145.040 37.750 1145.300 38.070 ;
        RECT 1138.660 2.400 1138.800 37.750 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1156.510 37.980 1156.830 38.040 ;
        RECT 1622.030 37.980 1622.350 38.040 ;
        RECT 1156.510 37.840 1622.350 37.980 ;
        RECT 1156.510 37.780 1156.830 37.840 ;
        RECT 1622.030 37.780 1622.350 37.840 ;
      LAYER via ;
        RECT 1156.540 37.780 1156.800 38.040 ;
        RECT 1622.060 37.780 1622.320 38.040 ;
      LAYER met2 ;
        RECT 1624.745 1700.410 1625.025 1704.000 ;
        RECT 1623.500 1700.270 1625.025 1700.410 ;
        RECT 1623.500 1678.650 1623.640 1700.270 ;
        RECT 1624.745 1700.000 1625.025 1700.270 ;
        RECT 1622.120 1678.510 1623.640 1678.650 ;
        RECT 1622.120 38.070 1622.260 1678.510 ;
        RECT 1156.540 37.750 1156.800 38.070 ;
        RECT 1622.060 37.750 1622.320 38.070 ;
        RECT 1156.600 2.400 1156.740 37.750 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1423.385 1193.825 1423.555 1241.935 ;
        RECT 1423.845 186.405 1424.015 234.515 ;
      LAYER mcon ;
        RECT 1423.385 1241.765 1423.555 1241.935 ;
        RECT 1423.845 234.345 1424.015 234.515 ;
      LAYER met1 ;
        RECT 1423.770 1559.620 1424.090 1559.880 ;
        RECT 1423.860 1559.200 1424.000 1559.620 ;
        RECT 1423.770 1558.940 1424.090 1559.200 ;
        RECT 1423.310 1497.260 1423.630 1497.320 ;
        RECT 1423.770 1497.260 1424.090 1497.320 ;
        RECT 1423.310 1497.120 1424.090 1497.260 ;
        RECT 1423.310 1497.060 1423.630 1497.120 ;
        RECT 1423.770 1497.060 1424.090 1497.120 ;
        RECT 1423.310 1490.460 1423.630 1490.520 ;
        RECT 1423.770 1490.460 1424.090 1490.520 ;
        RECT 1423.310 1490.320 1424.090 1490.460 ;
        RECT 1423.310 1490.260 1423.630 1490.320 ;
        RECT 1423.770 1490.260 1424.090 1490.320 ;
        RECT 1423.770 1400.700 1424.090 1400.760 ;
        RECT 1424.230 1400.700 1424.550 1400.760 ;
        RECT 1423.770 1400.560 1424.550 1400.700 ;
        RECT 1423.770 1400.500 1424.090 1400.560 ;
        RECT 1424.230 1400.500 1424.550 1400.560 ;
        RECT 1423.770 1297.340 1424.090 1297.400 ;
        RECT 1424.230 1297.340 1424.550 1297.400 ;
        RECT 1423.770 1297.200 1424.550 1297.340 ;
        RECT 1423.770 1297.140 1424.090 1297.200 ;
        RECT 1424.230 1297.140 1424.550 1297.200 ;
        RECT 1423.310 1255.860 1423.630 1255.920 ;
        RECT 1423.770 1255.860 1424.090 1255.920 ;
        RECT 1423.310 1255.720 1424.090 1255.860 ;
        RECT 1423.310 1255.660 1423.630 1255.720 ;
        RECT 1423.770 1255.660 1424.090 1255.720 ;
        RECT 1423.310 1241.920 1423.630 1241.980 ;
        RECT 1423.115 1241.780 1423.630 1241.920 ;
        RECT 1423.310 1241.720 1423.630 1241.780 ;
        RECT 1423.325 1193.980 1423.615 1194.025 ;
        RECT 1423.770 1193.980 1424.090 1194.040 ;
        RECT 1423.325 1193.840 1424.090 1193.980 ;
        RECT 1423.325 1193.795 1423.615 1193.840 ;
        RECT 1423.770 1193.780 1424.090 1193.840 ;
        RECT 1423.310 1062.740 1423.630 1062.800 ;
        RECT 1424.230 1062.740 1424.550 1062.800 ;
        RECT 1423.310 1062.600 1424.550 1062.740 ;
        RECT 1423.310 1062.540 1423.630 1062.600 ;
        RECT 1424.230 1062.540 1424.550 1062.600 ;
        RECT 1423.310 1028.200 1423.630 1028.460 ;
        RECT 1423.400 1027.720 1423.540 1028.200 ;
        RECT 1423.770 1027.720 1424.090 1027.780 ;
        RECT 1423.400 1027.580 1424.090 1027.720 ;
        RECT 1423.770 1027.520 1424.090 1027.580 ;
        RECT 1423.310 966.180 1423.630 966.240 ;
        RECT 1424.230 966.180 1424.550 966.240 ;
        RECT 1423.310 966.040 1424.550 966.180 ;
        RECT 1423.310 965.980 1423.630 966.040 ;
        RECT 1424.230 965.980 1424.550 966.040 ;
        RECT 1423.310 869.620 1423.630 869.680 ;
        RECT 1424.230 869.620 1424.550 869.680 ;
        RECT 1423.310 869.480 1424.550 869.620 ;
        RECT 1423.310 869.420 1423.630 869.480 ;
        RECT 1424.230 869.420 1424.550 869.480 ;
        RECT 1423.310 724.440 1423.630 724.500 ;
        RECT 1423.770 724.440 1424.090 724.500 ;
        RECT 1423.310 724.300 1424.090 724.440 ;
        RECT 1423.310 724.240 1423.630 724.300 ;
        RECT 1423.770 724.240 1424.090 724.300 ;
        RECT 1423.770 531.320 1424.090 531.380 ;
        RECT 1424.230 531.320 1424.550 531.380 ;
        RECT 1423.770 531.180 1424.550 531.320 ;
        RECT 1423.770 531.120 1424.090 531.180 ;
        RECT 1424.230 531.120 1424.550 531.180 ;
        RECT 1424.230 483.380 1424.550 483.440 ;
        RECT 1423.860 483.240 1424.550 483.380 ;
        RECT 1423.860 483.100 1424.000 483.240 ;
        RECT 1424.230 483.180 1424.550 483.240 ;
        RECT 1423.770 482.840 1424.090 483.100 ;
        RECT 1422.850 434.760 1423.170 434.820 ;
        RECT 1423.770 434.760 1424.090 434.820 ;
        RECT 1422.850 434.620 1424.090 434.760 ;
        RECT 1422.850 434.560 1423.170 434.620 ;
        RECT 1423.770 434.560 1424.090 434.620 ;
        RECT 1423.770 290.060 1424.090 290.320 ;
        RECT 1423.860 289.640 1424.000 290.060 ;
        RECT 1423.770 289.380 1424.090 289.640 ;
        RECT 1423.310 241.640 1423.630 241.700 ;
        RECT 1423.770 241.640 1424.090 241.700 ;
        RECT 1423.310 241.500 1424.090 241.640 ;
        RECT 1423.310 241.440 1423.630 241.500 ;
        RECT 1423.770 241.440 1424.090 241.500 ;
        RECT 1423.310 234.500 1423.630 234.560 ;
        RECT 1423.785 234.500 1424.075 234.545 ;
        RECT 1423.310 234.360 1424.075 234.500 ;
        RECT 1423.310 234.300 1423.630 234.360 ;
        RECT 1423.785 234.315 1424.075 234.360 ;
        RECT 1423.770 186.560 1424.090 186.620 ;
        RECT 1423.770 186.420 1424.285 186.560 ;
        RECT 1423.770 186.360 1424.090 186.420 ;
        RECT 1422.850 144.740 1423.170 144.800 ;
        RECT 1423.770 144.740 1424.090 144.800 ;
        RECT 1422.850 144.600 1424.090 144.740 ;
        RECT 1422.850 144.540 1423.170 144.600 ;
        RECT 1423.770 144.540 1424.090 144.600 ;
        RECT 674.430 37.640 674.750 37.700 ;
        RECT 1422.850 37.640 1423.170 37.700 ;
        RECT 674.430 37.500 1423.170 37.640 ;
        RECT 674.430 37.440 674.750 37.500 ;
        RECT 1422.850 37.440 1423.170 37.500 ;
      LAYER via ;
        RECT 1423.800 1559.620 1424.060 1559.880 ;
        RECT 1423.800 1558.940 1424.060 1559.200 ;
        RECT 1423.340 1497.060 1423.600 1497.320 ;
        RECT 1423.800 1497.060 1424.060 1497.320 ;
        RECT 1423.340 1490.260 1423.600 1490.520 ;
        RECT 1423.800 1490.260 1424.060 1490.520 ;
        RECT 1423.800 1400.500 1424.060 1400.760 ;
        RECT 1424.260 1400.500 1424.520 1400.760 ;
        RECT 1423.800 1297.140 1424.060 1297.400 ;
        RECT 1424.260 1297.140 1424.520 1297.400 ;
        RECT 1423.340 1255.660 1423.600 1255.920 ;
        RECT 1423.800 1255.660 1424.060 1255.920 ;
        RECT 1423.340 1241.720 1423.600 1241.980 ;
        RECT 1423.800 1193.780 1424.060 1194.040 ;
        RECT 1423.340 1062.540 1423.600 1062.800 ;
        RECT 1424.260 1062.540 1424.520 1062.800 ;
        RECT 1423.340 1028.200 1423.600 1028.460 ;
        RECT 1423.800 1027.520 1424.060 1027.780 ;
        RECT 1423.340 965.980 1423.600 966.240 ;
        RECT 1424.260 965.980 1424.520 966.240 ;
        RECT 1423.340 869.420 1423.600 869.680 ;
        RECT 1424.260 869.420 1424.520 869.680 ;
        RECT 1423.340 724.240 1423.600 724.500 ;
        RECT 1423.800 724.240 1424.060 724.500 ;
        RECT 1423.800 531.120 1424.060 531.380 ;
        RECT 1424.260 531.120 1424.520 531.380 ;
        RECT 1424.260 483.180 1424.520 483.440 ;
        RECT 1423.800 482.840 1424.060 483.100 ;
        RECT 1422.880 434.560 1423.140 434.820 ;
        RECT 1423.800 434.560 1424.060 434.820 ;
        RECT 1423.800 290.060 1424.060 290.320 ;
        RECT 1423.800 289.380 1424.060 289.640 ;
        RECT 1423.340 241.440 1423.600 241.700 ;
        RECT 1423.800 241.440 1424.060 241.700 ;
        RECT 1423.340 234.300 1423.600 234.560 ;
        RECT 1423.800 186.360 1424.060 186.620 ;
        RECT 1422.880 144.540 1423.140 144.800 ;
        RECT 1423.800 144.540 1424.060 144.800 ;
        RECT 674.460 37.440 674.720 37.700 ;
        RECT 1422.880 37.440 1423.140 37.700 ;
      LAYER met2 ;
        RECT 1426.485 1700.410 1426.765 1704.000 ;
        RECT 1425.700 1700.270 1426.765 1700.410 ;
        RECT 1425.700 1656.210 1425.840 1700.270 ;
        RECT 1426.485 1700.000 1426.765 1700.270 ;
        RECT 1423.860 1656.070 1425.840 1656.210 ;
        RECT 1423.860 1559.910 1424.000 1656.070 ;
        RECT 1423.800 1559.590 1424.060 1559.910 ;
        RECT 1423.800 1558.910 1424.060 1559.230 ;
        RECT 1423.860 1497.350 1424.000 1558.910 ;
        RECT 1423.340 1497.030 1423.600 1497.350 ;
        RECT 1423.800 1497.030 1424.060 1497.350 ;
        RECT 1423.400 1490.550 1423.540 1497.030 ;
        RECT 1423.340 1490.230 1423.600 1490.550 ;
        RECT 1423.800 1490.230 1424.060 1490.550 ;
        RECT 1423.860 1400.790 1424.000 1490.230 ;
        RECT 1423.800 1400.470 1424.060 1400.790 ;
        RECT 1424.260 1400.470 1424.520 1400.790 ;
        RECT 1424.320 1393.845 1424.460 1400.470 ;
        RECT 1423.330 1393.475 1423.610 1393.845 ;
        RECT 1424.250 1393.475 1424.530 1393.845 ;
        RECT 1423.400 1349.530 1423.540 1393.475 ;
        RECT 1423.400 1349.390 1424.460 1349.530 ;
        RECT 1424.320 1297.430 1424.460 1349.390 ;
        RECT 1423.800 1297.110 1424.060 1297.430 ;
        RECT 1424.260 1297.110 1424.520 1297.430 ;
        RECT 1423.860 1255.950 1424.000 1297.110 ;
        RECT 1423.340 1255.630 1423.600 1255.950 ;
        RECT 1423.800 1255.630 1424.060 1255.950 ;
        RECT 1423.400 1242.010 1423.540 1255.630 ;
        RECT 1423.340 1241.690 1423.600 1242.010 ;
        RECT 1423.800 1193.750 1424.060 1194.070 ;
        RECT 1423.860 1087.050 1424.000 1193.750 ;
        RECT 1423.860 1086.910 1424.460 1087.050 ;
        RECT 1424.320 1062.830 1424.460 1086.910 ;
        RECT 1423.340 1062.510 1423.600 1062.830 ;
        RECT 1424.260 1062.510 1424.520 1062.830 ;
        RECT 1423.400 1028.490 1423.540 1062.510 ;
        RECT 1423.340 1028.170 1423.600 1028.490 ;
        RECT 1423.800 1027.490 1424.060 1027.810 ;
        RECT 1423.860 990.490 1424.000 1027.490 ;
        RECT 1423.860 990.350 1424.460 990.490 ;
        RECT 1424.320 966.270 1424.460 990.350 ;
        RECT 1423.340 966.125 1423.600 966.270 ;
        RECT 1424.260 966.125 1424.520 966.270 ;
        RECT 1423.330 965.755 1423.610 966.125 ;
        RECT 1424.250 965.755 1424.530 966.125 ;
        RECT 1424.320 931.330 1424.460 965.755 ;
        RECT 1423.860 931.190 1424.460 931.330 ;
        RECT 1423.860 893.930 1424.000 931.190 ;
        RECT 1423.860 893.790 1424.460 893.930 ;
        RECT 1424.320 869.710 1424.460 893.790 ;
        RECT 1423.340 869.565 1423.600 869.710 ;
        RECT 1424.260 869.565 1424.520 869.710 ;
        RECT 1423.330 869.195 1423.610 869.565 ;
        RECT 1424.250 869.195 1424.530 869.565 ;
        RECT 1424.320 834.090 1424.460 869.195 ;
        RECT 1423.860 833.950 1424.460 834.090 ;
        RECT 1423.860 787.170 1424.000 833.950 ;
        RECT 1423.400 787.030 1424.000 787.170 ;
        RECT 1423.400 748.410 1423.540 787.030 ;
        RECT 1422.940 748.270 1423.540 748.410 ;
        RECT 1422.940 736.850 1423.080 748.270 ;
        RECT 1422.940 736.710 1424.000 736.850 ;
        RECT 1423.860 724.530 1424.000 736.710 ;
        RECT 1423.340 724.210 1423.600 724.530 ;
        RECT 1423.800 724.210 1424.060 724.530 ;
        RECT 1423.400 699.450 1423.540 724.210 ;
        RECT 1423.400 699.310 1424.000 699.450 ;
        RECT 1423.860 628.845 1424.000 699.310 ;
        RECT 1423.790 628.475 1424.070 628.845 ;
        RECT 1423.330 627.795 1423.610 628.165 ;
        RECT 1423.400 597.450 1423.540 627.795 ;
        RECT 1423.400 597.310 1424.460 597.450 ;
        RECT 1424.320 593.370 1424.460 597.310 ;
        RECT 1423.860 593.230 1424.460 593.370 ;
        RECT 1423.860 531.410 1424.000 593.230 ;
        RECT 1423.800 531.090 1424.060 531.410 ;
        RECT 1424.260 531.090 1424.520 531.410 ;
        RECT 1424.320 483.470 1424.460 531.090 ;
        RECT 1424.260 483.150 1424.520 483.470 ;
        RECT 1423.800 482.810 1424.060 483.130 ;
        RECT 1423.860 434.850 1424.000 482.810 ;
        RECT 1422.880 434.530 1423.140 434.850 ;
        RECT 1423.800 434.530 1424.060 434.850 ;
        RECT 1422.940 362.170 1423.080 434.530 ;
        RECT 1422.940 362.030 1424.000 362.170 ;
        RECT 1423.860 290.350 1424.000 362.030 ;
        RECT 1423.800 290.030 1424.060 290.350 ;
        RECT 1423.800 289.350 1424.060 289.670 ;
        RECT 1423.860 241.730 1424.000 289.350 ;
        RECT 1423.340 241.410 1423.600 241.730 ;
        RECT 1423.800 241.410 1424.060 241.730 ;
        RECT 1423.400 234.590 1423.540 241.410 ;
        RECT 1423.340 234.270 1423.600 234.590 ;
        RECT 1423.800 186.330 1424.060 186.650 ;
        RECT 1423.860 144.830 1424.000 186.330 ;
        RECT 1422.880 144.510 1423.140 144.830 ;
        RECT 1423.800 144.510 1424.060 144.830 ;
        RECT 1422.940 96.970 1423.080 144.510 ;
        RECT 1422.940 96.830 1423.540 96.970 ;
        RECT 1423.400 62.290 1423.540 96.830 ;
        RECT 1423.400 62.150 1424.000 62.290 ;
        RECT 1423.860 61.610 1424.000 62.150 ;
        RECT 1422.940 61.470 1424.000 61.610 ;
        RECT 1422.940 37.730 1423.080 61.470 ;
        RECT 674.460 37.410 674.720 37.730 ;
        RECT 1422.880 37.410 1423.140 37.730 ;
        RECT 674.520 2.400 674.660 37.410 ;
        RECT 674.310 -4.800 674.870 2.400 ;
      LAYER via2 ;
        RECT 1423.330 1393.520 1423.610 1393.800 ;
        RECT 1424.250 1393.520 1424.530 1393.800 ;
        RECT 1423.330 965.800 1423.610 966.080 ;
        RECT 1424.250 965.800 1424.530 966.080 ;
        RECT 1423.330 869.240 1423.610 869.520 ;
        RECT 1424.250 869.240 1424.530 869.520 ;
        RECT 1423.790 628.520 1424.070 628.800 ;
        RECT 1423.330 627.840 1423.610 628.120 ;
      LAYER met3 ;
        RECT 1423.305 1393.810 1423.635 1393.825 ;
        RECT 1424.225 1393.810 1424.555 1393.825 ;
        RECT 1423.305 1393.510 1424.555 1393.810 ;
        RECT 1423.305 1393.495 1423.635 1393.510 ;
        RECT 1424.225 1393.495 1424.555 1393.510 ;
        RECT 1423.305 966.090 1423.635 966.105 ;
        RECT 1424.225 966.090 1424.555 966.105 ;
        RECT 1423.305 965.790 1424.555 966.090 ;
        RECT 1423.305 965.775 1423.635 965.790 ;
        RECT 1424.225 965.775 1424.555 965.790 ;
        RECT 1423.305 869.530 1423.635 869.545 ;
        RECT 1424.225 869.530 1424.555 869.545 ;
        RECT 1423.305 869.230 1424.555 869.530 ;
        RECT 1423.305 869.215 1423.635 869.230 ;
        RECT 1424.225 869.215 1424.555 869.230 ;
        RECT 1423.765 628.810 1424.095 628.825 ;
        RECT 1423.550 628.495 1424.095 628.810 ;
        RECT 1423.550 628.145 1423.850 628.495 ;
        RECT 1423.305 627.830 1423.850 628.145 ;
        RECT 1423.305 627.815 1423.635 627.830 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1173.990 38.320 1174.310 38.380 ;
        RECT 1628.930 38.320 1629.250 38.380 ;
        RECT 1173.990 38.180 1629.250 38.320 ;
        RECT 1173.990 38.120 1174.310 38.180 ;
        RECT 1628.930 38.120 1629.250 38.180 ;
      LAYER via ;
        RECT 1174.020 38.120 1174.280 38.380 ;
        RECT 1628.960 38.120 1629.220 38.380 ;
      LAYER met2 ;
        RECT 1632.105 1700.410 1632.385 1704.000 ;
        RECT 1630.400 1700.270 1632.385 1700.410 ;
        RECT 1630.400 1677.970 1630.540 1700.270 ;
        RECT 1632.105 1700.000 1632.385 1700.270 ;
        RECT 1629.020 1677.830 1630.540 1677.970 ;
        RECT 1629.020 38.410 1629.160 1677.830 ;
        RECT 1174.020 38.090 1174.280 38.410 ;
        RECT 1628.960 38.090 1629.220 38.410 ;
        RECT 1174.080 2.400 1174.220 38.090 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1636.365 1587.205 1636.535 1635.315 ;
        RECT 1635.905 1393.745 1636.075 1401.055 ;
        RECT 1635.905 965.685 1636.075 1007.335 ;
        RECT 1635.905 482.885 1636.075 517.395 ;
        RECT 1635.905 282.965 1636.075 331.075 ;
        RECT 1636.825 234.685 1636.995 241.655 ;
      LAYER mcon ;
        RECT 1636.365 1635.145 1636.535 1635.315 ;
        RECT 1635.905 1400.885 1636.075 1401.055 ;
        RECT 1635.905 1007.165 1636.075 1007.335 ;
        RECT 1635.905 517.225 1636.075 517.395 ;
        RECT 1635.905 330.905 1636.075 331.075 ;
        RECT 1636.825 241.485 1636.995 241.655 ;
      LAYER met1 ;
        RECT 1636.750 1692.080 1637.070 1692.140 ;
        RECT 1639.510 1692.080 1639.830 1692.140 ;
        RECT 1636.750 1691.940 1639.830 1692.080 ;
        RECT 1636.750 1691.880 1637.070 1691.940 ;
        RECT 1639.510 1691.880 1639.830 1691.940 ;
        RECT 1636.290 1635.300 1636.610 1635.360 ;
        RECT 1636.095 1635.160 1636.610 1635.300 ;
        RECT 1636.290 1635.100 1636.610 1635.160 ;
        RECT 1636.290 1587.360 1636.610 1587.420 ;
        RECT 1636.095 1587.220 1636.610 1587.360 ;
        RECT 1636.290 1587.160 1636.610 1587.220 ;
        RECT 1635.830 1545.680 1636.150 1545.940 ;
        RECT 1635.920 1545.260 1636.060 1545.680 ;
        RECT 1635.830 1545.000 1636.150 1545.260 ;
        RECT 1635.830 1401.040 1636.150 1401.100 ;
        RECT 1635.635 1400.900 1636.150 1401.040 ;
        RECT 1635.830 1400.840 1636.150 1400.900 ;
        RECT 1635.830 1393.900 1636.150 1393.960 ;
        RECT 1635.635 1393.760 1636.150 1393.900 ;
        RECT 1635.830 1393.700 1636.150 1393.760 ;
        RECT 1635.830 1352.760 1636.150 1352.820 ;
        RECT 1636.290 1352.760 1636.610 1352.820 ;
        RECT 1635.830 1352.620 1636.610 1352.760 ;
        RECT 1635.830 1352.560 1636.150 1352.620 ;
        RECT 1636.290 1352.560 1636.610 1352.620 ;
        RECT 1636.290 1304.820 1636.610 1304.880 ;
        RECT 1635.920 1304.680 1636.610 1304.820 ;
        RECT 1635.920 1303.860 1636.060 1304.680 ;
        RECT 1636.290 1304.620 1636.610 1304.680 ;
        RECT 1635.830 1303.600 1636.150 1303.860 ;
        RECT 1636.290 1159.300 1636.610 1159.360 ;
        RECT 1636.750 1159.300 1637.070 1159.360 ;
        RECT 1636.290 1159.160 1637.070 1159.300 ;
        RECT 1636.290 1159.100 1636.610 1159.160 ;
        RECT 1636.750 1159.100 1637.070 1159.160 ;
        RECT 1636.290 1111.360 1636.610 1111.420 ;
        RECT 1635.920 1111.220 1636.610 1111.360 ;
        RECT 1635.920 1111.080 1636.060 1111.220 ;
        RECT 1636.290 1111.160 1636.610 1111.220 ;
        RECT 1635.830 1110.820 1636.150 1111.080 ;
        RECT 1635.830 1062.740 1636.150 1062.800 ;
        RECT 1636.290 1062.740 1636.610 1062.800 ;
        RECT 1635.830 1062.600 1636.610 1062.740 ;
        RECT 1635.830 1062.540 1636.150 1062.600 ;
        RECT 1636.290 1062.540 1636.610 1062.600 ;
        RECT 1636.290 1014.800 1636.610 1014.860 ;
        RECT 1635.920 1014.660 1636.610 1014.800 ;
        RECT 1635.920 1014.520 1636.060 1014.660 ;
        RECT 1636.290 1014.600 1636.610 1014.660 ;
        RECT 1635.830 1014.260 1636.150 1014.520 ;
        RECT 1635.830 1007.320 1636.150 1007.380 ;
        RECT 1635.635 1007.180 1636.150 1007.320 ;
        RECT 1635.830 1007.120 1636.150 1007.180 ;
        RECT 1635.845 965.840 1636.135 965.885 ;
        RECT 1636.290 965.840 1636.610 965.900 ;
        RECT 1635.845 965.700 1636.610 965.840 ;
        RECT 1635.845 965.655 1636.135 965.700 ;
        RECT 1636.290 965.640 1636.610 965.700 ;
        RECT 1635.830 917.900 1636.150 917.960 ;
        RECT 1636.750 917.900 1637.070 917.960 ;
        RECT 1635.830 917.760 1637.070 917.900 ;
        RECT 1635.830 917.700 1636.150 917.760 ;
        RECT 1636.750 917.700 1637.070 917.760 ;
        RECT 1635.830 869.620 1636.150 869.680 ;
        RECT 1636.290 869.620 1636.610 869.680 ;
        RECT 1635.830 869.480 1636.610 869.620 ;
        RECT 1635.830 869.420 1636.150 869.480 ;
        RECT 1636.290 869.420 1636.610 869.480 ;
        RECT 1635.830 517.380 1636.150 517.440 ;
        RECT 1635.635 517.240 1636.150 517.380 ;
        RECT 1635.830 517.180 1636.150 517.240 ;
        RECT 1635.830 483.040 1636.150 483.100 ;
        RECT 1635.635 482.900 1636.150 483.040 ;
        RECT 1635.830 482.840 1636.150 482.900 ;
        RECT 1635.830 434.560 1636.150 434.820 ;
        RECT 1635.920 434.420 1636.060 434.560 ;
        RECT 1636.290 434.420 1636.610 434.480 ;
        RECT 1635.920 434.280 1636.610 434.420 ;
        RECT 1636.290 434.220 1636.610 434.280 ;
        RECT 1636.290 352.480 1636.610 352.540 ;
        RECT 1635.920 352.340 1636.610 352.480 ;
        RECT 1635.920 351.860 1636.060 352.340 ;
        RECT 1636.290 352.280 1636.610 352.340 ;
        RECT 1635.830 351.600 1636.150 351.860 ;
        RECT 1635.830 331.060 1636.150 331.120 ;
        RECT 1635.635 330.920 1636.150 331.060 ;
        RECT 1635.830 330.860 1636.150 330.920 ;
        RECT 1635.845 283.120 1636.135 283.165 ;
        RECT 1637.210 283.120 1637.530 283.180 ;
        RECT 1635.845 282.980 1637.530 283.120 ;
        RECT 1635.845 282.935 1636.135 282.980 ;
        RECT 1637.210 282.920 1637.530 282.980 ;
        RECT 1636.750 241.640 1637.070 241.700 ;
        RECT 1636.555 241.500 1637.070 241.640 ;
        RECT 1636.750 241.440 1637.070 241.500 ;
        RECT 1636.750 234.840 1637.070 234.900 ;
        RECT 1636.555 234.700 1637.070 234.840 ;
        RECT 1636.750 234.640 1637.070 234.700 ;
        RECT 1636.290 193.360 1636.610 193.420 ;
        RECT 1636.750 193.360 1637.070 193.420 ;
        RECT 1636.290 193.220 1637.070 193.360 ;
        RECT 1636.290 193.160 1636.610 193.220 ;
        RECT 1636.750 193.160 1637.070 193.220 ;
        RECT 1191.930 34.920 1192.250 34.980 ;
        RECT 1636.290 34.920 1636.610 34.980 ;
        RECT 1191.930 34.780 1636.610 34.920 ;
        RECT 1191.930 34.720 1192.250 34.780 ;
        RECT 1636.290 34.720 1636.610 34.780 ;
      LAYER via ;
        RECT 1636.780 1691.880 1637.040 1692.140 ;
        RECT 1639.540 1691.880 1639.800 1692.140 ;
        RECT 1636.320 1635.100 1636.580 1635.360 ;
        RECT 1636.320 1587.160 1636.580 1587.420 ;
        RECT 1635.860 1545.680 1636.120 1545.940 ;
        RECT 1635.860 1545.000 1636.120 1545.260 ;
        RECT 1635.860 1400.840 1636.120 1401.100 ;
        RECT 1635.860 1393.700 1636.120 1393.960 ;
        RECT 1635.860 1352.560 1636.120 1352.820 ;
        RECT 1636.320 1352.560 1636.580 1352.820 ;
        RECT 1636.320 1304.620 1636.580 1304.880 ;
        RECT 1635.860 1303.600 1636.120 1303.860 ;
        RECT 1636.320 1159.100 1636.580 1159.360 ;
        RECT 1636.780 1159.100 1637.040 1159.360 ;
        RECT 1636.320 1111.160 1636.580 1111.420 ;
        RECT 1635.860 1110.820 1636.120 1111.080 ;
        RECT 1635.860 1062.540 1636.120 1062.800 ;
        RECT 1636.320 1062.540 1636.580 1062.800 ;
        RECT 1636.320 1014.600 1636.580 1014.860 ;
        RECT 1635.860 1014.260 1636.120 1014.520 ;
        RECT 1635.860 1007.120 1636.120 1007.380 ;
        RECT 1636.320 965.640 1636.580 965.900 ;
        RECT 1635.860 917.700 1636.120 917.960 ;
        RECT 1636.780 917.700 1637.040 917.960 ;
        RECT 1635.860 869.420 1636.120 869.680 ;
        RECT 1636.320 869.420 1636.580 869.680 ;
        RECT 1635.860 517.180 1636.120 517.440 ;
        RECT 1635.860 482.840 1636.120 483.100 ;
        RECT 1635.860 434.560 1636.120 434.820 ;
        RECT 1636.320 434.220 1636.580 434.480 ;
        RECT 1636.320 352.280 1636.580 352.540 ;
        RECT 1635.860 351.600 1636.120 351.860 ;
        RECT 1635.860 330.860 1636.120 331.120 ;
        RECT 1637.240 282.920 1637.500 283.180 ;
        RECT 1636.780 241.440 1637.040 241.700 ;
        RECT 1636.780 234.640 1637.040 234.900 ;
        RECT 1636.320 193.160 1636.580 193.420 ;
        RECT 1636.780 193.160 1637.040 193.420 ;
        RECT 1191.960 34.720 1192.220 34.980 ;
        RECT 1636.320 34.720 1636.580 34.980 ;
      LAYER met2 ;
        RECT 1639.465 1700.000 1639.745 1704.000 ;
        RECT 1639.600 1692.170 1639.740 1700.000 ;
        RECT 1636.780 1691.850 1637.040 1692.170 ;
        RECT 1639.540 1691.850 1639.800 1692.170 ;
        RECT 1636.840 1655.530 1636.980 1691.850 ;
        RECT 1636.380 1655.390 1636.980 1655.530 ;
        RECT 1636.380 1635.390 1636.520 1655.390 ;
        RECT 1636.320 1635.070 1636.580 1635.390 ;
        RECT 1636.320 1587.130 1636.580 1587.450 ;
        RECT 1636.380 1586.850 1636.520 1587.130 ;
        RECT 1635.920 1586.710 1636.520 1586.850 ;
        RECT 1635.920 1545.970 1636.060 1586.710 ;
        RECT 1635.860 1545.650 1636.120 1545.970 ;
        RECT 1635.860 1544.970 1636.120 1545.290 ;
        RECT 1635.920 1401.130 1636.060 1544.970 ;
        RECT 1635.860 1400.810 1636.120 1401.130 ;
        RECT 1635.860 1393.670 1636.120 1393.990 ;
        RECT 1635.920 1352.850 1636.060 1393.670 ;
        RECT 1635.860 1352.530 1636.120 1352.850 ;
        RECT 1636.320 1352.530 1636.580 1352.850 ;
        RECT 1636.380 1304.910 1636.520 1352.530 ;
        RECT 1636.320 1304.590 1636.580 1304.910 ;
        RECT 1635.860 1303.570 1636.120 1303.890 ;
        RECT 1635.920 1297.285 1636.060 1303.570 ;
        RECT 1635.850 1296.915 1636.130 1297.285 ;
        RECT 1636.770 1296.235 1637.050 1296.605 ;
        RECT 1636.840 1159.390 1636.980 1296.235 ;
        RECT 1636.320 1159.070 1636.580 1159.390 ;
        RECT 1636.780 1159.070 1637.040 1159.390 ;
        RECT 1636.380 1111.450 1636.520 1159.070 ;
        RECT 1636.320 1111.130 1636.580 1111.450 ;
        RECT 1635.860 1110.790 1636.120 1111.110 ;
        RECT 1635.920 1062.830 1636.060 1110.790 ;
        RECT 1635.860 1062.510 1636.120 1062.830 ;
        RECT 1636.320 1062.510 1636.580 1062.830 ;
        RECT 1636.380 1014.890 1636.520 1062.510 ;
        RECT 1636.320 1014.570 1636.580 1014.890 ;
        RECT 1635.860 1014.230 1636.120 1014.550 ;
        RECT 1635.920 1007.410 1636.060 1014.230 ;
        RECT 1635.860 1007.090 1636.120 1007.410 ;
        RECT 1636.320 965.610 1636.580 965.930 ;
        RECT 1636.380 959.210 1636.520 965.610 ;
        RECT 1636.380 959.070 1636.980 959.210 ;
        RECT 1636.840 917.990 1636.980 959.070 ;
        RECT 1635.860 917.670 1636.120 917.990 ;
        RECT 1636.780 917.670 1637.040 917.990 ;
        RECT 1635.920 869.710 1636.060 917.670 ;
        RECT 1635.860 869.390 1636.120 869.710 ;
        RECT 1636.320 869.390 1636.580 869.710 ;
        RECT 1636.380 830.690 1636.520 869.390 ;
        RECT 1636.380 830.550 1637.440 830.690 ;
        RECT 1637.300 814.485 1637.440 830.550 ;
        RECT 1636.310 814.115 1636.590 814.485 ;
        RECT 1637.230 814.115 1637.510 814.485 ;
        RECT 1636.380 742.290 1636.520 814.115 ;
        RECT 1636.380 742.150 1636.980 742.290 ;
        RECT 1636.840 688.570 1636.980 742.150 ;
        RECT 1636.380 688.430 1636.980 688.570 ;
        RECT 1636.380 651.850 1636.520 688.430 ;
        RECT 1635.920 651.710 1636.520 651.850 ;
        RECT 1635.920 566.965 1636.060 651.710 ;
        RECT 1635.850 566.595 1636.130 566.965 ;
        RECT 1635.850 565.915 1636.130 566.285 ;
        RECT 1635.920 517.470 1636.060 565.915 ;
        RECT 1635.860 517.150 1636.120 517.470 ;
        RECT 1635.860 482.810 1636.120 483.130 ;
        RECT 1635.920 434.850 1636.060 482.810 ;
        RECT 1635.860 434.530 1636.120 434.850 ;
        RECT 1636.320 434.190 1636.580 434.510 ;
        RECT 1636.380 352.570 1636.520 434.190 ;
        RECT 1636.320 352.250 1636.580 352.570 ;
        RECT 1635.860 351.570 1636.120 351.890 ;
        RECT 1635.920 331.150 1636.060 351.570 ;
        RECT 1635.860 330.830 1636.120 331.150 ;
        RECT 1637.240 282.890 1637.500 283.210 ;
        RECT 1637.300 282.610 1637.440 282.890 ;
        RECT 1636.840 282.470 1637.440 282.610 ;
        RECT 1636.840 241.730 1636.980 282.470 ;
        RECT 1636.780 241.410 1637.040 241.730 ;
        RECT 1636.780 234.610 1637.040 234.930 ;
        RECT 1636.840 193.450 1636.980 234.610 ;
        RECT 1636.320 193.130 1636.580 193.450 ;
        RECT 1636.780 193.130 1637.040 193.450 ;
        RECT 1636.380 35.010 1636.520 193.130 ;
        RECT 1191.960 34.690 1192.220 35.010 ;
        RECT 1636.320 34.690 1636.580 35.010 ;
        RECT 1192.020 2.400 1192.160 34.690 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
      LAYER via2 ;
        RECT 1635.850 1296.960 1636.130 1297.240 ;
        RECT 1636.770 1296.280 1637.050 1296.560 ;
        RECT 1636.310 814.160 1636.590 814.440 ;
        RECT 1637.230 814.160 1637.510 814.440 ;
        RECT 1635.850 566.640 1636.130 566.920 ;
        RECT 1635.850 565.960 1636.130 566.240 ;
      LAYER met3 ;
        RECT 1635.825 1297.250 1636.155 1297.265 ;
        RECT 1635.150 1296.950 1636.155 1297.250 ;
        RECT 1635.150 1296.570 1635.450 1296.950 ;
        RECT 1635.825 1296.935 1636.155 1296.950 ;
        RECT 1636.745 1296.570 1637.075 1296.585 ;
        RECT 1635.150 1296.270 1637.075 1296.570 ;
        RECT 1636.745 1296.255 1637.075 1296.270 ;
        RECT 1636.285 814.450 1636.615 814.465 ;
        RECT 1637.205 814.450 1637.535 814.465 ;
        RECT 1636.285 814.150 1637.535 814.450 ;
        RECT 1636.285 814.135 1636.615 814.150 ;
        RECT 1637.205 814.135 1637.535 814.150 ;
        RECT 1635.825 566.930 1636.155 566.945 ;
        RECT 1635.825 566.615 1636.370 566.930 ;
        RECT 1636.070 566.265 1636.370 566.615 ;
        RECT 1635.825 565.950 1636.370 566.265 ;
        RECT 1635.825 565.935 1636.155 565.950 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1642.730 1658.420 1643.050 1658.480 ;
        RECT 1645.030 1658.420 1645.350 1658.480 ;
        RECT 1642.730 1658.280 1645.350 1658.420 ;
        RECT 1642.730 1658.220 1643.050 1658.280 ;
        RECT 1645.030 1658.220 1645.350 1658.280 ;
        RECT 1209.870 38.660 1210.190 38.720 ;
        RECT 1642.730 38.660 1643.050 38.720 ;
        RECT 1209.870 38.520 1643.050 38.660 ;
        RECT 1209.870 38.460 1210.190 38.520 ;
        RECT 1642.730 38.460 1643.050 38.520 ;
      LAYER via ;
        RECT 1642.760 1658.220 1643.020 1658.480 ;
        RECT 1645.060 1658.220 1645.320 1658.480 ;
        RECT 1209.900 38.460 1210.160 38.720 ;
        RECT 1642.760 38.460 1643.020 38.720 ;
      LAYER met2 ;
        RECT 1646.825 1700.410 1647.105 1704.000 ;
        RECT 1645.120 1700.270 1647.105 1700.410 ;
        RECT 1645.120 1658.510 1645.260 1700.270 ;
        RECT 1646.825 1700.000 1647.105 1700.270 ;
        RECT 1642.760 1658.190 1643.020 1658.510 ;
        RECT 1645.060 1658.190 1645.320 1658.510 ;
        RECT 1642.820 38.750 1642.960 1658.190 ;
        RECT 1209.900 38.430 1210.160 38.750 ;
        RECT 1642.760 38.430 1643.020 38.750 ;
        RECT 1209.960 2.400 1210.100 38.430 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1651.085 1538.925 1651.255 1587.035 ;
        RECT 1650.625 1013.965 1650.795 1055.615 ;
        RECT 1651.085 724.625 1651.255 813.875 ;
        RECT 1650.625 493.425 1650.795 517.055 ;
        RECT 1649.705 421.005 1649.875 469.115 ;
        RECT 1650.625 289.085 1650.795 307.275 ;
        RECT 1651.085 48.365 1651.255 129.455 ;
      LAYER mcon ;
        RECT 1651.085 1586.865 1651.255 1587.035 ;
        RECT 1650.625 1055.445 1650.795 1055.615 ;
        RECT 1651.085 813.705 1651.255 813.875 ;
        RECT 1650.625 516.885 1650.795 517.055 ;
        RECT 1649.705 468.945 1649.875 469.115 ;
        RECT 1650.625 307.105 1650.795 307.275 ;
        RECT 1651.085 129.285 1651.255 129.455 ;
      LAYER met1 ;
        RECT 1651.010 1587.020 1651.330 1587.080 ;
        RECT 1650.815 1586.880 1651.330 1587.020 ;
        RECT 1651.010 1586.820 1651.330 1586.880 ;
        RECT 1651.010 1539.080 1651.330 1539.140 ;
        RECT 1650.815 1538.940 1651.330 1539.080 ;
        RECT 1651.010 1538.880 1651.330 1538.940 ;
        RECT 1650.550 1442.180 1650.870 1442.240 ;
        RECT 1651.010 1442.180 1651.330 1442.240 ;
        RECT 1650.550 1442.040 1651.330 1442.180 ;
        RECT 1650.550 1441.980 1650.870 1442.040 ;
        RECT 1651.010 1441.980 1651.330 1442.040 ;
        RECT 1649.630 1394.580 1649.950 1394.640 ;
        RECT 1651.010 1394.580 1651.330 1394.640 ;
        RECT 1649.630 1394.440 1651.330 1394.580 ;
        RECT 1649.630 1394.380 1649.950 1394.440 ;
        RECT 1651.010 1394.380 1651.330 1394.440 ;
        RECT 1649.630 1338.820 1649.950 1338.880 ;
        RECT 1650.550 1338.820 1650.870 1338.880 ;
        RECT 1649.630 1338.680 1650.870 1338.820 ;
        RECT 1649.630 1338.620 1649.950 1338.680 ;
        RECT 1650.550 1338.620 1650.870 1338.680 ;
        RECT 1650.550 1290.200 1650.870 1290.260 ;
        RECT 1651.470 1290.200 1651.790 1290.260 ;
        RECT 1650.550 1290.060 1651.790 1290.200 ;
        RECT 1650.550 1290.000 1650.870 1290.060 ;
        RECT 1651.470 1290.000 1651.790 1290.060 ;
        RECT 1649.630 1224.920 1649.950 1224.980 ;
        RECT 1651.010 1224.920 1651.330 1224.980 ;
        RECT 1649.630 1224.780 1651.330 1224.920 ;
        RECT 1649.630 1224.720 1649.950 1224.780 ;
        RECT 1651.010 1224.720 1651.330 1224.780 ;
        RECT 1651.010 1152.500 1651.330 1152.560 ;
        RECT 1651.930 1152.500 1652.250 1152.560 ;
        RECT 1651.010 1152.360 1652.250 1152.500 ;
        RECT 1651.010 1152.300 1651.330 1152.360 ;
        RECT 1651.930 1152.300 1652.250 1152.360 ;
        RECT 1650.550 1111.020 1650.870 1111.080 ;
        RECT 1651.010 1111.020 1651.330 1111.080 ;
        RECT 1650.550 1110.880 1651.330 1111.020 ;
        RECT 1650.550 1110.820 1650.870 1110.880 ;
        RECT 1651.010 1110.820 1651.330 1110.880 ;
        RECT 1651.010 1062.880 1651.330 1063.140 ;
        RECT 1651.100 1062.460 1651.240 1062.880 ;
        RECT 1651.010 1062.200 1651.330 1062.460 ;
        RECT 1650.565 1055.600 1650.855 1055.645 ;
        RECT 1651.470 1055.600 1651.790 1055.660 ;
        RECT 1650.565 1055.460 1651.790 1055.600 ;
        RECT 1650.565 1055.415 1650.855 1055.460 ;
        RECT 1651.470 1055.400 1651.790 1055.460 ;
        RECT 1650.550 1014.120 1650.870 1014.180 ;
        RECT 1650.355 1013.980 1650.870 1014.120 ;
        RECT 1650.550 1013.920 1650.870 1013.980 ;
        RECT 1650.550 1007.320 1650.870 1007.380 ;
        RECT 1651.470 1007.320 1651.790 1007.380 ;
        RECT 1650.550 1007.180 1651.790 1007.320 ;
        RECT 1650.550 1007.120 1650.870 1007.180 ;
        RECT 1651.470 1007.120 1651.790 1007.180 ;
        RECT 1651.470 1000.520 1651.790 1000.580 ;
        RECT 1652.390 1000.520 1652.710 1000.580 ;
        RECT 1651.470 1000.380 1652.710 1000.520 ;
        RECT 1651.470 1000.320 1651.790 1000.380 ;
        RECT 1652.390 1000.320 1652.710 1000.380 ;
        RECT 1649.630 910.420 1649.950 910.480 ;
        RECT 1650.550 910.420 1650.870 910.480 ;
        RECT 1649.630 910.280 1650.870 910.420 ;
        RECT 1649.630 910.220 1649.950 910.280 ;
        RECT 1650.550 910.220 1650.870 910.280 ;
        RECT 1649.630 862.480 1649.950 862.540 ;
        RECT 1651.010 862.480 1651.330 862.540 ;
        RECT 1649.630 862.340 1651.330 862.480 ;
        RECT 1649.630 862.280 1649.950 862.340 ;
        RECT 1651.010 862.280 1651.330 862.340 ;
        RECT 1650.550 813.860 1650.870 813.920 ;
        RECT 1651.025 813.860 1651.315 813.905 ;
        RECT 1650.550 813.720 1651.315 813.860 ;
        RECT 1650.550 813.660 1650.870 813.720 ;
        RECT 1651.025 813.675 1651.315 813.720 ;
        RECT 1651.010 724.780 1651.330 724.840 ;
        RECT 1650.815 724.640 1651.330 724.780 ;
        RECT 1651.010 724.580 1651.330 724.640 ;
        RECT 1649.630 717.640 1649.950 717.700 ;
        RECT 1651.010 717.640 1651.330 717.700 ;
        RECT 1649.630 717.500 1651.330 717.640 ;
        RECT 1649.630 717.440 1649.950 717.500 ;
        RECT 1651.010 717.440 1651.330 717.500 ;
        RECT 1650.550 627.880 1650.870 627.940 ;
        RECT 1651.470 627.880 1651.790 627.940 ;
        RECT 1650.550 627.740 1651.790 627.880 ;
        RECT 1650.550 627.680 1650.870 627.740 ;
        RECT 1651.470 627.680 1651.790 627.740 ;
        RECT 1650.550 517.040 1650.870 517.100 ;
        RECT 1650.355 516.900 1650.870 517.040 ;
        RECT 1650.550 516.840 1650.870 516.900 ;
        RECT 1650.565 493.580 1650.855 493.625 ;
        RECT 1651.010 493.580 1651.330 493.640 ;
        RECT 1650.565 493.440 1651.330 493.580 ;
        RECT 1650.565 493.395 1650.855 493.440 ;
        RECT 1651.010 493.380 1651.330 493.440 ;
        RECT 1649.645 469.100 1649.935 469.145 ;
        RECT 1650.550 469.100 1650.870 469.160 ;
        RECT 1649.645 468.960 1650.870 469.100 ;
        RECT 1649.645 468.915 1649.935 468.960 ;
        RECT 1650.550 468.900 1650.870 468.960 ;
        RECT 1649.630 421.160 1649.950 421.220 ;
        RECT 1649.435 421.020 1649.950 421.160 ;
        RECT 1649.630 420.960 1649.950 421.020 ;
        RECT 1649.630 338.200 1649.950 338.260 ;
        RECT 1650.550 338.200 1650.870 338.260 ;
        RECT 1649.630 338.060 1650.870 338.200 ;
        RECT 1649.630 338.000 1649.950 338.060 ;
        RECT 1650.550 338.000 1650.870 338.060 ;
        RECT 1650.550 307.260 1650.870 307.320 ;
        RECT 1650.355 307.120 1650.870 307.260 ;
        RECT 1650.550 307.060 1650.870 307.120 ;
        RECT 1650.565 289.240 1650.855 289.285 ;
        RECT 1651.470 289.240 1651.790 289.300 ;
        RECT 1650.565 289.100 1651.790 289.240 ;
        RECT 1650.565 289.055 1650.855 289.100 ;
        RECT 1651.470 289.040 1651.790 289.100 ;
        RECT 1649.630 193.360 1649.950 193.420 ;
        RECT 1651.010 193.360 1651.330 193.420 ;
        RECT 1649.630 193.220 1651.330 193.360 ;
        RECT 1649.630 193.160 1649.950 193.220 ;
        RECT 1651.010 193.160 1651.330 193.220 ;
        RECT 1649.630 131.480 1649.950 131.540 ;
        RECT 1651.010 131.480 1651.330 131.540 ;
        RECT 1649.630 131.340 1651.330 131.480 ;
        RECT 1649.630 131.280 1649.950 131.340 ;
        RECT 1651.010 131.280 1651.330 131.340 ;
        RECT 1649.630 129.440 1649.950 129.500 ;
        RECT 1651.025 129.440 1651.315 129.485 ;
        RECT 1649.630 129.300 1651.315 129.440 ;
        RECT 1649.630 129.240 1649.950 129.300 ;
        RECT 1651.025 129.255 1651.315 129.300 ;
        RECT 1651.010 48.520 1651.330 48.580 ;
        RECT 1650.815 48.380 1651.330 48.520 ;
        RECT 1651.010 48.320 1651.330 48.380 ;
        RECT 1227.810 39.000 1228.130 39.060 ;
        RECT 1651.010 39.000 1651.330 39.060 ;
        RECT 1227.810 38.860 1651.330 39.000 ;
        RECT 1227.810 38.800 1228.130 38.860 ;
        RECT 1651.010 38.800 1651.330 38.860 ;
      LAYER via ;
        RECT 1651.040 1586.820 1651.300 1587.080 ;
        RECT 1651.040 1538.880 1651.300 1539.140 ;
        RECT 1650.580 1441.980 1650.840 1442.240 ;
        RECT 1651.040 1441.980 1651.300 1442.240 ;
        RECT 1649.660 1394.380 1649.920 1394.640 ;
        RECT 1651.040 1394.380 1651.300 1394.640 ;
        RECT 1649.660 1338.620 1649.920 1338.880 ;
        RECT 1650.580 1338.620 1650.840 1338.880 ;
        RECT 1650.580 1290.000 1650.840 1290.260 ;
        RECT 1651.500 1290.000 1651.760 1290.260 ;
        RECT 1649.660 1224.720 1649.920 1224.980 ;
        RECT 1651.040 1224.720 1651.300 1224.980 ;
        RECT 1651.040 1152.300 1651.300 1152.560 ;
        RECT 1651.960 1152.300 1652.220 1152.560 ;
        RECT 1650.580 1110.820 1650.840 1111.080 ;
        RECT 1651.040 1110.820 1651.300 1111.080 ;
        RECT 1651.040 1062.880 1651.300 1063.140 ;
        RECT 1651.040 1062.200 1651.300 1062.460 ;
        RECT 1651.500 1055.400 1651.760 1055.660 ;
        RECT 1650.580 1013.920 1650.840 1014.180 ;
        RECT 1650.580 1007.120 1650.840 1007.380 ;
        RECT 1651.500 1007.120 1651.760 1007.380 ;
        RECT 1651.500 1000.320 1651.760 1000.580 ;
        RECT 1652.420 1000.320 1652.680 1000.580 ;
        RECT 1649.660 910.220 1649.920 910.480 ;
        RECT 1650.580 910.220 1650.840 910.480 ;
        RECT 1649.660 862.280 1649.920 862.540 ;
        RECT 1651.040 862.280 1651.300 862.540 ;
        RECT 1650.580 813.660 1650.840 813.920 ;
        RECT 1651.040 724.580 1651.300 724.840 ;
        RECT 1649.660 717.440 1649.920 717.700 ;
        RECT 1651.040 717.440 1651.300 717.700 ;
        RECT 1650.580 627.680 1650.840 627.940 ;
        RECT 1651.500 627.680 1651.760 627.940 ;
        RECT 1650.580 516.840 1650.840 517.100 ;
        RECT 1651.040 493.380 1651.300 493.640 ;
        RECT 1650.580 468.900 1650.840 469.160 ;
        RECT 1649.660 420.960 1649.920 421.220 ;
        RECT 1649.660 338.000 1649.920 338.260 ;
        RECT 1650.580 338.000 1650.840 338.260 ;
        RECT 1650.580 307.060 1650.840 307.320 ;
        RECT 1651.500 289.040 1651.760 289.300 ;
        RECT 1649.660 193.160 1649.920 193.420 ;
        RECT 1651.040 193.160 1651.300 193.420 ;
        RECT 1649.660 131.280 1649.920 131.540 ;
        RECT 1651.040 131.280 1651.300 131.540 ;
        RECT 1649.660 129.240 1649.920 129.500 ;
        RECT 1651.040 48.320 1651.300 48.580 ;
        RECT 1227.840 38.800 1228.100 39.060 ;
        RECT 1651.040 38.800 1651.300 39.060 ;
      LAYER met2 ;
        RECT 1654.185 1700.410 1654.465 1704.000 ;
        RECT 1652.940 1700.270 1654.465 1700.410 ;
        RECT 1652.940 1658.930 1653.080 1700.270 ;
        RECT 1654.185 1700.000 1654.465 1700.270 ;
        RECT 1651.100 1658.790 1653.080 1658.930 ;
        RECT 1651.100 1587.110 1651.240 1658.790 ;
        RECT 1651.040 1586.790 1651.300 1587.110 ;
        RECT 1651.040 1538.850 1651.300 1539.170 ;
        RECT 1651.100 1497.770 1651.240 1538.850 ;
        RECT 1650.640 1497.630 1651.240 1497.770 ;
        RECT 1650.640 1442.270 1650.780 1497.630 ;
        RECT 1650.580 1441.950 1650.840 1442.270 ;
        RECT 1651.040 1441.950 1651.300 1442.270 ;
        RECT 1651.100 1394.670 1651.240 1441.950 ;
        RECT 1649.660 1394.350 1649.920 1394.670 ;
        RECT 1651.040 1394.350 1651.300 1394.670 ;
        RECT 1649.720 1338.910 1649.860 1394.350 ;
        RECT 1649.660 1338.590 1649.920 1338.910 ;
        RECT 1650.580 1338.590 1650.840 1338.910 ;
        RECT 1650.640 1290.290 1650.780 1338.590 ;
        RECT 1650.580 1289.970 1650.840 1290.290 ;
        RECT 1651.500 1289.970 1651.760 1290.290 ;
        RECT 1651.560 1242.205 1651.700 1289.970 ;
        RECT 1649.650 1241.835 1649.930 1242.205 ;
        RECT 1651.490 1241.835 1651.770 1242.205 ;
        RECT 1649.720 1225.010 1649.860 1241.835 ;
        RECT 1649.660 1224.690 1649.920 1225.010 ;
        RECT 1651.040 1224.690 1651.300 1225.010 ;
        RECT 1651.100 1200.725 1651.240 1224.690 ;
        RECT 1651.030 1200.355 1651.310 1200.725 ;
        RECT 1651.950 1200.355 1652.230 1200.725 ;
        RECT 1652.020 1152.590 1652.160 1200.355 ;
        RECT 1651.040 1152.270 1651.300 1152.590 ;
        RECT 1651.960 1152.270 1652.220 1152.590 ;
        RECT 1650.640 1111.110 1650.780 1111.265 ;
        RECT 1651.100 1111.110 1651.240 1152.270 ;
        RECT 1650.580 1110.850 1650.840 1111.110 ;
        RECT 1651.040 1110.850 1651.300 1111.110 ;
        RECT 1650.580 1110.790 1651.300 1110.850 ;
        RECT 1650.640 1110.710 1651.240 1110.790 ;
        RECT 1651.100 1063.170 1651.240 1110.710 ;
        RECT 1651.040 1062.850 1651.300 1063.170 ;
        RECT 1651.040 1062.170 1651.300 1062.490 ;
        RECT 1651.100 1055.770 1651.240 1062.170 ;
        RECT 1651.100 1055.690 1651.700 1055.770 ;
        RECT 1651.100 1055.630 1651.760 1055.690 ;
        RECT 1651.500 1055.370 1651.760 1055.630 ;
        RECT 1651.560 1055.215 1651.700 1055.370 ;
        RECT 1650.580 1013.890 1650.840 1014.210 ;
        RECT 1650.640 1007.410 1650.780 1013.890 ;
        RECT 1650.580 1007.090 1650.840 1007.410 ;
        RECT 1651.500 1007.090 1651.760 1007.410 ;
        RECT 1651.560 1000.610 1651.700 1007.090 ;
        RECT 1651.500 1000.290 1651.760 1000.610 ;
        RECT 1652.420 1000.290 1652.680 1000.610 ;
        RECT 1652.480 952.525 1652.620 1000.290 ;
        RECT 1651.490 952.155 1651.770 952.525 ;
        RECT 1652.410 952.155 1652.690 952.525 ;
        RECT 1651.560 911.045 1651.700 952.155 ;
        RECT 1650.570 910.675 1650.850 911.045 ;
        RECT 1651.490 910.675 1651.770 911.045 ;
        RECT 1650.640 910.510 1650.780 910.675 ;
        RECT 1649.660 910.190 1649.920 910.510 ;
        RECT 1650.580 910.190 1650.840 910.510 ;
        RECT 1649.720 862.765 1649.860 910.190 ;
        RECT 1649.650 862.395 1649.930 862.765 ;
        RECT 1651.030 862.395 1651.310 862.765 ;
        RECT 1649.660 862.250 1649.920 862.395 ;
        RECT 1651.040 862.250 1651.300 862.395 ;
        RECT 1649.720 814.485 1649.860 862.250 ;
        RECT 1649.650 814.115 1649.930 814.485 ;
        RECT 1650.570 814.115 1650.850 814.485 ;
        RECT 1650.640 813.950 1650.780 814.115 ;
        RECT 1650.580 813.630 1650.840 813.950 ;
        RECT 1651.040 724.550 1651.300 724.870 ;
        RECT 1651.100 717.730 1651.240 724.550 ;
        RECT 1649.660 717.410 1649.920 717.730 ;
        RECT 1651.040 717.410 1651.300 717.730 ;
        RECT 1649.720 628.165 1649.860 717.410 ;
        RECT 1649.650 627.795 1649.930 628.165 ;
        RECT 1650.570 627.795 1650.850 628.165 ;
        RECT 1650.580 627.650 1650.840 627.795 ;
        RECT 1651.500 627.650 1651.760 627.970 ;
        RECT 1651.560 572.460 1651.700 627.650 ;
        RECT 1650.640 572.320 1651.700 572.460 ;
        RECT 1650.640 517.130 1650.780 572.320 ;
        RECT 1650.580 516.810 1650.840 517.130 ;
        RECT 1651.040 493.350 1651.300 493.670 ;
        RECT 1651.100 469.610 1651.240 493.350 ;
        RECT 1650.640 469.470 1651.240 469.610 ;
        RECT 1650.640 469.190 1650.780 469.470 ;
        RECT 1650.580 468.870 1650.840 469.190 ;
        RECT 1649.660 420.930 1649.920 421.250 ;
        RECT 1649.720 338.290 1649.860 420.930 ;
        RECT 1649.660 337.970 1649.920 338.290 ;
        RECT 1650.580 337.970 1650.840 338.290 ;
        RECT 1650.640 307.350 1650.780 337.970 ;
        RECT 1650.580 307.030 1650.840 307.350 ;
        RECT 1651.500 289.010 1651.760 289.330 ;
        RECT 1651.560 241.925 1651.700 289.010 ;
        RECT 1651.490 241.555 1651.770 241.925 ;
        RECT 1649.650 240.875 1649.930 241.245 ;
        RECT 1649.720 193.450 1649.860 240.875 ;
        RECT 1649.660 193.130 1649.920 193.450 ;
        RECT 1651.040 193.130 1651.300 193.450 ;
        RECT 1651.100 131.570 1651.240 193.130 ;
        RECT 1649.660 131.250 1649.920 131.570 ;
        RECT 1651.040 131.250 1651.300 131.570 ;
        RECT 1649.720 129.530 1649.860 131.250 ;
        RECT 1649.660 129.210 1649.920 129.530 ;
        RECT 1651.040 48.290 1651.300 48.610 ;
        RECT 1651.100 39.090 1651.240 48.290 ;
        RECT 1227.840 38.770 1228.100 39.090 ;
        RECT 1651.040 38.770 1651.300 39.090 ;
        RECT 1227.900 2.400 1228.040 38.770 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
      LAYER via2 ;
        RECT 1649.650 1241.880 1649.930 1242.160 ;
        RECT 1651.490 1241.880 1651.770 1242.160 ;
        RECT 1651.030 1200.400 1651.310 1200.680 ;
        RECT 1651.950 1200.400 1652.230 1200.680 ;
        RECT 1651.490 952.200 1651.770 952.480 ;
        RECT 1652.410 952.200 1652.690 952.480 ;
        RECT 1650.570 910.720 1650.850 911.000 ;
        RECT 1651.490 910.720 1651.770 911.000 ;
        RECT 1649.650 862.440 1649.930 862.720 ;
        RECT 1651.030 862.440 1651.310 862.720 ;
        RECT 1649.650 814.160 1649.930 814.440 ;
        RECT 1650.570 814.160 1650.850 814.440 ;
        RECT 1649.650 627.840 1649.930 628.120 ;
        RECT 1650.570 627.840 1650.850 628.120 ;
        RECT 1651.490 241.600 1651.770 241.880 ;
        RECT 1649.650 240.920 1649.930 241.200 ;
      LAYER met3 ;
        RECT 1649.625 1242.170 1649.955 1242.185 ;
        RECT 1651.465 1242.170 1651.795 1242.185 ;
        RECT 1649.625 1241.870 1651.795 1242.170 ;
        RECT 1649.625 1241.855 1649.955 1241.870 ;
        RECT 1651.465 1241.855 1651.795 1241.870 ;
        RECT 1651.005 1200.690 1651.335 1200.705 ;
        RECT 1651.925 1200.690 1652.255 1200.705 ;
        RECT 1651.005 1200.390 1652.255 1200.690 ;
        RECT 1651.005 1200.375 1651.335 1200.390 ;
        RECT 1651.925 1200.375 1652.255 1200.390 ;
        RECT 1651.465 952.490 1651.795 952.505 ;
        RECT 1652.385 952.490 1652.715 952.505 ;
        RECT 1651.465 952.190 1652.715 952.490 ;
        RECT 1651.465 952.175 1651.795 952.190 ;
        RECT 1652.385 952.175 1652.715 952.190 ;
        RECT 1650.545 911.010 1650.875 911.025 ;
        RECT 1651.465 911.010 1651.795 911.025 ;
        RECT 1650.545 910.710 1651.795 911.010 ;
        RECT 1650.545 910.695 1650.875 910.710 ;
        RECT 1651.465 910.695 1651.795 910.710 ;
        RECT 1649.625 862.730 1649.955 862.745 ;
        RECT 1651.005 862.730 1651.335 862.745 ;
        RECT 1649.625 862.430 1651.335 862.730 ;
        RECT 1649.625 862.415 1649.955 862.430 ;
        RECT 1651.005 862.415 1651.335 862.430 ;
        RECT 1649.625 814.450 1649.955 814.465 ;
        RECT 1650.545 814.450 1650.875 814.465 ;
        RECT 1649.625 814.150 1650.875 814.450 ;
        RECT 1649.625 814.135 1649.955 814.150 ;
        RECT 1650.545 814.135 1650.875 814.150 ;
        RECT 1649.625 628.130 1649.955 628.145 ;
        RECT 1650.545 628.130 1650.875 628.145 ;
        RECT 1649.625 627.830 1650.875 628.130 ;
        RECT 1649.625 627.815 1649.955 627.830 ;
        RECT 1650.545 627.815 1650.875 627.830 ;
        RECT 1651.465 241.890 1651.795 241.905 ;
        RECT 1649.870 241.590 1651.795 241.890 ;
        RECT 1649.870 241.225 1650.170 241.590 ;
        RECT 1651.465 241.575 1651.795 241.590 ;
        RECT 1649.625 240.910 1650.170 241.225 ;
        RECT 1649.625 240.895 1649.955 240.910 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1656.530 1678.480 1656.850 1678.540 ;
        RECT 1659.750 1678.480 1660.070 1678.540 ;
        RECT 1656.530 1678.340 1660.070 1678.480 ;
        RECT 1656.530 1678.280 1656.850 1678.340 ;
        RECT 1659.750 1678.280 1660.070 1678.340 ;
        RECT 1245.750 39.340 1246.070 39.400 ;
        RECT 1656.530 39.340 1656.850 39.400 ;
        RECT 1245.750 39.200 1656.850 39.340 ;
        RECT 1245.750 39.140 1246.070 39.200 ;
        RECT 1656.530 39.140 1656.850 39.200 ;
      LAYER via ;
        RECT 1656.560 1678.280 1656.820 1678.540 ;
        RECT 1659.780 1678.280 1660.040 1678.540 ;
        RECT 1245.780 39.140 1246.040 39.400 ;
        RECT 1656.560 39.140 1656.820 39.400 ;
      LAYER met2 ;
        RECT 1661.545 1700.410 1661.825 1704.000 ;
        RECT 1659.840 1700.270 1661.825 1700.410 ;
        RECT 1659.840 1678.570 1659.980 1700.270 ;
        RECT 1661.545 1700.000 1661.825 1700.270 ;
        RECT 1656.560 1678.250 1656.820 1678.570 ;
        RECT 1659.780 1678.250 1660.040 1678.570 ;
        RECT 1656.620 39.430 1656.760 1678.250 ;
        RECT 1245.780 39.110 1246.040 39.430 ;
        RECT 1656.560 39.110 1656.820 39.430 ;
        RECT 1245.840 2.400 1245.980 39.110 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1663.430 1675.420 1663.750 1675.480 ;
        RECT 1667.110 1675.420 1667.430 1675.480 ;
        RECT 1663.430 1675.280 1667.430 1675.420 ;
        RECT 1663.430 1675.220 1663.750 1675.280 ;
        RECT 1667.110 1675.220 1667.430 1675.280 ;
        RECT 1263.230 39.680 1263.550 39.740 ;
        RECT 1663.430 39.680 1663.750 39.740 ;
        RECT 1263.230 39.540 1663.750 39.680 ;
        RECT 1263.230 39.480 1263.550 39.540 ;
        RECT 1663.430 39.480 1663.750 39.540 ;
      LAYER via ;
        RECT 1663.460 1675.220 1663.720 1675.480 ;
        RECT 1667.140 1675.220 1667.400 1675.480 ;
        RECT 1263.260 39.480 1263.520 39.740 ;
        RECT 1663.460 39.480 1663.720 39.740 ;
      LAYER met2 ;
        RECT 1668.905 1700.410 1669.185 1704.000 ;
        RECT 1667.200 1700.270 1669.185 1700.410 ;
        RECT 1667.200 1675.510 1667.340 1700.270 ;
        RECT 1668.905 1700.000 1669.185 1700.270 ;
        RECT 1663.460 1675.190 1663.720 1675.510 ;
        RECT 1667.140 1675.190 1667.400 1675.510 ;
        RECT 1663.520 39.770 1663.660 1675.190 ;
        RECT 1263.260 39.450 1263.520 39.770 ;
        RECT 1663.460 39.450 1663.720 39.770 ;
        RECT 1263.320 2.400 1263.460 39.450 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1670.330 1678.480 1670.650 1678.540 ;
        RECT 1674.470 1678.480 1674.790 1678.540 ;
        RECT 1670.330 1678.340 1674.790 1678.480 ;
        RECT 1670.330 1678.280 1670.650 1678.340 ;
        RECT 1674.470 1678.280 1674.790 1678.340 ;
        RECT 1281.170 40.020 1281.490 40.080 ;
        RECT 1670.330 40.020 1670.650 40.080 ;
        RECT 1281.170 39.880 1670.650 40.020 ;
        RECT 1281.170 39.820 1281.490 39.880 ;
        RECT 1670.330 39.820 1670.650 39.880 ;
      LAYER via ;
        RECT 1670.360 1678.280 1670.620 1678.540 ;
        RECT 1674.500 1678.280 1674.760 1678.540 ;
        RECT 1281.200 39.820 1281.460 40.080 ;
        RECT 1670.360 39.820 1670.620 40.080 ;
      LAYER met2 ;
        RECT 1676.265 1700.410 1676.545 1704.000 ;
        RECT 1674.560 1700.270 1676.545 1700.410 ;
        RECT 1674.560 1678.570 1674.700 1700.270 ;
        RECT 1676.265 1700.000 1676.545 1700.270 ;
        RECT 1670.360 1678.250 1670.620 1678.570 ;
        RECT 1674.500 1678.250 1674.760 1678.570 ;
        RECT 1670.420 40.110 1670.560 1678.250 ;
        RECT 1281.200 39.790 1281.460 40.110 ;
        RECT 1670.360 39.790 1670.620 40.110 ;
        RECT 1281.260 2.400 1281.400 39.790 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1683.670 1659.440 1683.990 1659.500 ;
        RECT 1684.590 1659.440 1684.910 1659.500 ;
        RECT 1683.670 1659.300 1684.910 1659.440 ;
        RECT 1683.670 1659.240 1683.990 1659.300 ;
        RECT 1684.590 1659.240 1684.910 1659.300 ;
        RECT 1299.110 40.360 1299.430 40.420 ;
        RECT 1684.590 40.360 1684.910 40.420 ;
        RECT 1299.110 40.220 1684.910 40.360 ;
        RECT 1299.110 40.160 1299.430 40.220 ;
        RECT 1684.590 40.160 1684.910 40.220 ;
      LAYER via ;
        RECT 1683.700 1659.240 1683.960 1659.500 ;
        RECT 1684.620 1659.240 1684.880 1659.500 ;
        RECT 1299.140 40.160 1299.400 40.420 ;
        RECT 1684.620 40.160 1684.880 40.420 ;
      LAYER met2 ;
        RECT 1683.625 1700.000 1683.905 1704.000 ;
        RECT 1683.760 1659.530 1683.900 1700.000 ;
        RECT 1683.700 1659.210 1683.960 1659.530 ;
        RECT 1684.620 1659.210 1684.880 1659.530 ;
        RECT 1684.680 40.450 1684.820 1659.210 ;
        RECT 1299.140 40.130 1299.400 40.450 ;
        RECT 1684.620 40.130 1684.880 40.450 ;
        RECT 1299.200 2.400 1299.340 40.130 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.050 40.700 1317.370 40.760 ;
        RECT 1691.490 40.700 1691.810 40.760 ;
        RECT 1317.050 40.560 1691.810 40.700 ;
        RECT 1317.050 40.500 1317.370 40.560 ;
        RECT 1691.490 40.500 1691.810 40.560 ;
      LAYER via ;
        RECT 1317.080 40.500 1317.340 40.760 ;
        RECT 1691.520 40.500 1691.780 40.760 ;
      LAYER met2 ;
        RECT 1690.985 1700.410 1691.265 1704.000 ;
        RECT 1690.985 1700.270 1691.720 1700.410 ;
        RECT 1690.985 1700.000 1691.265 1700.270 ;
        RECT 1691.580 40.790 1691.720 1700.270 ;
        RECT 1317.080 40.470 1317.340 40.790 ;
        RECT 1691.520 40.470 1691.780 40.790 ;
        RECT 1317.140 2.400 1317.280 40.470 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1334.990 41.040 1335.310 41.100 ;
        RECT 1697.930 41.040 1698.250 41.100 ;
        RECT 1334.990 40.900 1698.250 41.040 ;
        RECT 1334.990 40.840 1335.310 40.900 ;
        RECT 1697.930 40.840 1698.250 40.900 ;
      LAYER via ;
        RECT 1335.020 40.840 1335.280 41.100 ;
        RECT 1697.960 40.840 1698.220 41.100 ;
      LAYER met2 ;
        RECT 1698.345 1700.410 1698.625 1704.000 ;
        RECT 1698.020 1700.270 1698.625 1700.410 ;
        RECT 1698.020 41.130 1698.160 1700.270 ;
        RECT 1698.345 1700.000 1698.625 1700.270 ;
        RECT 1335.020 40.810 1335.280 41.130 ;
        RECT 1697.960 40.810 1698.220 41.130 ;
        RECT 1335.080 2.400 1335.220 40.810 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1430.285 1235.305 1430.455 1279.675 ;
        RECT 1430.285 1014.305 1430.455 1062.415 ;
        RECT 1429.825 758.965 1429.995 807.075 ;
        RECT 1429.825 517.565 1429.995 565.675 ;
        RECT 1430.285 379.525 1430.455 424.915 ;
      LAYER mcon ;
        RECT 1430.285 1279.505 1430.455 1279.675 ;
        RECT 1430.285 1062.245 1430.455 1062.415 ;
        RECT 1429.825 806.905 1429.995 807.075 ;
        RECT 1429.825 565.505 1429.995 565.675 ;
        RECT 1430.285 424.745 1430.455 424.915 ;
      LAYER met1 ;
        RECT 1429.750 1677.460 1430.070 1677.520 ;
        RECT 1432.970 1677.460 1433.290 1677.520 ;
        RECT 1429.750 1677.320 1433.290 1677.460 ;
        RECT 1429.750 1677.260 1430.070 1677.320 ;
        RECT 1432.970 1677.260 1433.290 1677.320 ;
        RECT 1428.830 1580.220 1429.150 1580.280 ;
        RECT 1430.210 1580.220 1430.530 1580.280 ;
        RECT 1428.830 1580.080 1430.530 1580.220 ;
        RECT 1428.830 1580.020 1429.150 1580.080 ;
        RECT 1430.210 1580.020 1430.530 1580.080 ;
        RECT 1430.670 1531.940 1430.990 1532.000 ;
        RECT 1431.130 1531.940 1431.450 1532.000 ;
        RECT 1430.670 1531.800 1431.450 1531.940 ;
        RECT 1430.670 1531.740 1430.990 1531.800 ;
        RECT 1431.130 1531.740 1431.450 1531.800 ;
        RECT 1430.210 1491.140 1430.530 1491.200 ;
        RECT 1430.670 1491.140 1430.990 1491.200 ;
        RECT 1430.210 1491.000 1430.990 1491.140 ;
        RECT 1430.210 1490.940 1430.530 1491.000 ;
        RECT 1430.670 1490.940 1430.990 1491.000 ;
        RECT 1430.210 1490.460 1430.530 1490.520 ;
        RECT 1430.670 1490.460 1430.990 1490.520 ;
        RECT 1430.210 1490.320 1430.990 1490.460 ;
        RECT 1430.210 1490.260 1430.530 1490.320 ;
        RECT 1430.670 1490.260 1430.990 1490.320 ;
        RECT 1430.210 1352.420 1430.530 1352.480 ;
        RECT 1430.670 1352.420 1430.990 1352.480 ;
        RECT 1430.210 1352.280 1430.990 1352.420 ;
        RECT 1430.210 1352.220 1430.530 1352.280 ;
        RECT 1430.670 1352.220 1430.990 1352.280 ;
        RECT 1430.225 1279.660 1430.515 1279.705 ;
        RECT 1430.670 1279.660 1430.990 1279.720 ;
        RECT 1430.225 1279.520 1430.990 1279.660 ;
        RECT 1430.225 1279.475 1430.515 1279.520 ;
        RECT 1430.670 1279.460 1430.990 1279.520 ;
        RECT 1430.210 1235.460 1430.530 1235.520 ;
        RECT 1430.015 1235.320 1430.530 1235.460 ;
        RECT 1430.210 1235.260 1430.530 1235.320 ;
        RECT 1429.750 1193.440 1430.070 1193.700 ;
        RECT 1429.840 1192.960 1429.980 1193.440 ;
        RECT 1430.670 1192.960 1430.990 1193.020 ;
        RECT 1429.840 1192.820 1430.990 1192.960 ;
        RECT 1430.670 1192.760 1430.990 1192.820 ;
        RECT 1430.210 1062.400 1430.530 1062.460 ;
        RECT 1430.015 1062.260 1430.530 1062.400 ;
        RECT 1430.210 1062.200 1430.530 1062.260 ;
        RECT 1430.225 1014.460 1430.515 1014.505 ;
        RECT 1430.670 1014.460 1430.990 1014.520 ;
        RECT 1430.225 1014.320 1430.990 1014.460 ;
        RECT 1430.225 1014.275 1430.515 1014.320 ;
        RECT 1430.670 1014.260 1430.990 1014.320 ;
        RECT 1429.750 959.040 1430.070 959.100 ;
        RECT 1430.210 959.040 1430.530 959.100 ;
        RECT 1429.750 958.900 1430.530 959.040 ;
        RECT 1429.750 958.840 1430.070 958.900 ;
        RECT 1430.210 958.840 1430.530 958.900 ;
        RECT 1429.750 821.140 1430.070 821.400 ;
        RECT 1429.840 820.660 1429.980 821.140 ;
        RECT 1430.670 820.660 1430.990 820.720 ;
        RECT 1429.840 820.520 1430.990 820.660 ;
        RECT 1430.670 820.460 1430.990 820.520 ;
        RECT 1429.765 807.060 1430.055 807.105 ;
        RECT 1430.670 807.060 1430.990 807.120 ;
        RECT 1429.765 806.920 1430.990 807.060 ;
        RECT 1429.765 806.875 1430.055 806.920 ;
        RECT 1430.670 806.860 1430.990 806.920 ;
        RECT 1429.750 759.120 1430.070 759.180 ;
        RECT 1429.555 758.980 1430.070 759.120 ;
        RECT 1429.750 758.920 1430.070 758.980 ;
        RECT 1428.830 688.740 1429.150 688.800 ;
        RECT 1430.670 688.740 1430.990 688.800 ;
        RECT 1428.830 688.600 1430.990 688.740 ;
        RECT 1428.830 688.540 1429.150 688.600 ;
        RECT 1430.670 688.540 1430.990 688.600 ;
        RECT 1429.750 613.940 1430.070 614.000 ;
        RECT 1430.210 613.940 1430.530 614.000 ;
        RECT 1429.750 613.800 1430.530 613.940 ;
        RECT 1429.750 613.740 1430.070 613.800 ;
        RECT 1430.210 613.740 1430.530 613.800 ;
        RECT 1429.750 565.660 1430.070 565.720 ;
        RECT 1429.555 565.520 1430.070 565.660 ;
        RECT 1429.750 565.460 1430.070 565.520 ;
        RECT 1429.765 517.720 1430.055 517.765 ;
        RECT 1430.210 517.720 1430.530 517.780 ;
        RECT 1429.765 517.580 1430.530 517.720 ;
        RECT 1429.765 517.535 1430.055 517.580 ;
        RECT 1430.210 517.520 1430.530 517.580 ;
        RECT 1430.225 424.900 1430.515 424.945 ;
        RECT 1430.670 424.900 1430.990 424.960 ;
        RECT 1430.225 424.760 1430.990 424.900 ;
        RECT 1430.225 424.715 1430.515 424.760 ;
        RECT 1430.670 424.700 1430.990 424.760 ;
        RECT 1430.225 379.680 1430.515 379.725 ;
        RECT 1430.670 379.680 1430.990 379.740 ;
        RECT 1430.225 379.540 1430.990 379.680 ;
        RECT 1430.225 379.495 1430.515 379.540 ;
        RECT 1430.670 379.480 1430.990 379.540 ;
        RECT 1430.210 234.500 1430.530 234.560 ;
        RECT 1430.670 234.500 1430.990 234.560 ;
        RECT 1430.210 234.360 1430.990 234.500 ;
        RECT 1430.210 234.300 1430.530 234.360 ;
        RECT 1430.670 234.300 1430.990 234.360 ;
        RECT 692.370 37.300 692.690 37.360 ;
        RECT 1429.750 37.300 1430.070 37.360 ;
        RECT 692.370 37.160 1430.070 37.300 ;
        RECT 692.370 37.100 692.690 37.160 ;
        RECT 1429.750 37.100 1430.070 37.160 ;
      LAYER via ;
        RECT 1429.780 1677.260 1430.040 1677.520 ;
        RECT 1433.000 1677.260 1433.260 1677.520 ;
        RECT 1428.860 1580.020 1429.120 1580.280 ;
        RECT 1430.240 1580.020 1430.500 1580.280 ;
        RECT 1430.700 1531.740 1430.960 1532.000 ;
        RECT 1431.160 1531.740 1431.420 1532.000 ;
        RECT 1430.240 1490.940 1430.500 1491.200 ;
        RECT 1430.700 1490.940 1430.960 1491.200 ;
        RECT 1430.240 1490.260 1430.500 1490.520 ;
        RECT 1430.700 1490.260 1430.960 1490.520 ;
        RECT 1430.240 1352.220 1430.500 1352.480 ;
        RECT 1430.700 1352.220 1430.960 1352.480 ;
        RECT 1430.700 1279.460 1430.960 1279.720 ;
        RECT 1430.240 1235.260 1430.500 1235.520 ;
        RECT 1429.780 1193.440 1430.040 1193.700 ;
        RECT 1430.700 1192.760 1430.960 1193.020 ;
        RECT 1430.240 1062.200 1430.500 1062.460 ;
        RECT 1430.700 1014.260 1430.960 1014.520 ;
        RECT 1429.780 958.840 1430.040 959.100 ;
        RECT 1430.240 958.840 1430.500 959.100 ;
        RECT 1429.780 821.140 1430.040 821.400 ;
        RECT 1430.700 820.460 1430.960 820.720 ;
        RECT 1430.700 806.860 1430.960 807.120 ;
        RECT 1429.780 758.920 1430.040 759.180 ;
        RECT 1428.860 688.540 1429.120 688.800 ;
        RECT 1430.700 688.540 1430.960 688.800 ;
        RECT 1429.780 613.740 1430.040 614.000 ;
        RECT 1430.240 613.740 1430.500 614.000 ;
        RECT 1429.780 565.460 1430.040 565.720 ;
        RECT 1430.240 517.520 1430.500 517.780 ;
        RECT 1430.700 424.700 1430.960 424.960 ;
        RECT 1430.700 379.480 1430.960 379.740 ;
        RECT 1430.240 234.300 1430.500 234.560 ;
        RECT 1430.700 234.300 1430.960 234.560 ;
        RECT 692.400 37.100 692.660 37.360 ;
        RECT 1429.780 37.100 1430.040 37.360 ;
      LAYER met2 ;
        RECT 1433.845 1700.410 1434.125 1704.000 ;
        RECT 1433.060 1700.270 1434.125 1700.410 ;
        RECT 1433.060 1677.550 1433.200 1700.270 ;
        RECT 1433.845 1700.000 1434.125 1700.270 ;
        RECT 1429.780 1677.230 1430.040 1677.550 ;
        RECT 1433.000 1677.230 1433.260 1677.550 ;
        RECT 1429.840 1628.445 1429.980 1677.230 ;
        RECT 1428.850 1628.075 1429.130 1628.445 ;
        RECT 1429.770 1628.075 1430.050 1628.445 ;
        RECT 1428.920 1580.310 1429.060 1628.075 ;
        RECT 1428.860 1579.990 1429.120 1580.310 ;
        RECT 1430.240 1580.165 1430.500 1580.310 ;
        RECT 1430.230 1579.795 1430.510 1580.165 ;
        RECT 1431.150 1579.795 1431.430 1580.165 ;
        RECT 1431.220 1532.030 1431.360 1579.795 ;
        RECT 1430.700 1531.710 1430.960 1532.030 ;
        RECT 1431.160 1531.710 1431.420 1532.030 ;
        RECT 1430.760 1491.230 1430.900 1531.710 ;
        RECT 1430.240 1490.910 1430.500 1491.230 ;
        RECT 1430.700 1490.910 1430.960 1491.230 ;
        RECT 1430.300 1490.550 1430.440 1490.910 ;
        RECT 1430.240 1490.230 1430.500 1490.550 ;
        RECT 1430.700 1490.230 1430.960 1490.550 ;
        RECT 1430.760 1376.050 1430.900 1490.230 ;
        RECT 1430.300 1375.910 1430.900 1376.050 ;
        RECT 1430.300 1352.510 1430.440 1375.910 ;
        RECT 1430.240 1352.190 1430.500 1352.510 ;
        RECT 1430.700 1352.190 1430.960 1352.510 ;
        RECT 1430.760 1279.750 1430.900 1352.190 ;
        RECT 1430.700 1279.430 1430.960 1279.750 ;
        RECT 1430.240 1235.230 1430.500 1235.550 ;
        RECT 1430.300 1194.605 1430.440 1235.230 ;
        RECT 1430.230 1194.235 1430.510 1194.605 ;
        RECT 1429.770 1193.555 1430.050 1193.925 ;
        RECT 1429.780 1193.410 1430.040 1193.555 ;
        RECT 1430.700 1192.730 1430.960 1193.050 ;
        RECT 1430.760 1086.370 1430.900 1192.730 ;
        RECT 1430.300 1086.230 1430.900 1086.370 ;
        RECT 1430.300 1062.490 1430.440 1086.230 ;
        RECT 1430.240 1062.170 1430.500 1062.490 ;
        RECT 1430.700 1014.230 1430.960 1014.550 ;
        RECT 1430.760 989.810 1430.900 1014.230 ;
        RECT 1430.300 989.670 1430.900 989.810 ;
        RECT 1430.300 959.130 1430.440 989.670 ;
        RECT 1429.780 958.810 1430.040 959.130 ;
        RECT 1430.240 958.810 1430.500 959.130 ;
        RECT 1429.840 911.045 1429.980 958.810 ;
        RECT 1429.770 910.675 1430.050 911.045 ;
        RECT 1430.690 910.675 1430.970 911.045 ;
        RECT 1430.760 869.565 1430.900 910.675 ;
        RECT 1429.770 869.195 1430.050 869.565 ;
        RECT 1430.690 869.195 1430.970 869.565 ;
        RECT 1429.840 821.430 1429.980 869.195 ;
        RECT 1429.780 821.110 1430.040 821.430 ;
        RECT 1430.700 820.430 1430.960 820.750 ;
        RECT 1430.760 807.150 1430.900 820.430 ;
        RECT 1430.700 806.830 1430.960 807.150 ;
        RECT 1429.780 758.890 1430.040 759.210 ;
        RECT 1429.840 738.890 1429.980 758.890 ;
        RECT 1429.840 738.750 1430.440 738.890 ;
        RECT 1430.300 717.810 1430.440 738.750 ;
        RECT 1430.300 717.670 1430.900 717.810 ;
        RECT 1430.760 688.830 1430.900 717.670 ;
        RECT 1428.860 688.510 1429.120 688.830 ;
        RECT 1430.700 688.510 1430.960 688.830 ;
        RECT 1428.920 621.365 1429.060 688.510 ;
        RECT 1428.850 620.995 1429.130 621.365 ;
        RECT 1429.770 620.995 1430.050 621.365 ;
        RECT 1429.840 614.030 1429.980 620.995 ;
        RECT 1429.780 613.710 1430.040 614.030 ;
        RECT 1430.240 613.710 1430.500 614.030 ;
        RECT 1430.300 566.170 1430.440 613.710 ;
        RECT 1429.840 566.030 1430.440 566.170 ;
        RECT 1429.840 565.750 1429.980 566.030 ;
        RECT 1429.780 565.430 1430.040 565.750 ;
        RECT 1430.240 517.490 1430.500 517.810 ;
        RECT 1430.300 468.930 1430.440 517.490 ;
        RECT 1430.300 468.790 1430.900 468.930 ;
        RECT 1430.760 424.990 1430.900 468.790 ;
        RECT 1430.700 424.670 1430.960 424.990 ;
        RECT 1430.700 379.450 1430.960 379.770 ;
        RECT 1430.760 379.170 1430.900 379.450 ;
        RECT 1430.760 379.030 1431.360 379.170 ;
        RECT 1431.220 283.405 1431.360 379.030 ;
        RECT 1430.230 283.035 1430.510 283.405 ;
        RECT 1431.150 283.035 1431.430 283.405 ;
        RECT 1430.300 234.590 1430.440 283.035 ;
        RECT 1430.240 234.270 1430.500 234.590 ;
        RECT 1430.700 234.270 1430.960 234.590 ;
        RECT 1430.760 130.290 1430.900 234.270 ;
        RECT 1430.300 130.150 1430.900 130.290 ;
        RECT 1430.300 61.610 1430.440 130.150 ;
        RECT 1429.840 61.470 1430.440 61.610 ;
        RECT 1429.840 37.390 1429.980 61.470 ;
        RECT 692.400 37.070 692.660 37.390 ;
        RECT 1429.780 37.070 1430.040 37.390 ;
        RECT 692.460 2.400 692.600 37.070 ;
        RECT 692.250 -4.800 692.810 2.400 ;
      LAYER via2 ;
        RECT 1428.850 1628.120 1429.130 1628.400 ;
        RECT 1429.770 1628.120 1430.050 1628.400 ;
        RECT 1430.230 1579.840 1430.510 1580.120 ;
        RECT 1431.150 1579.840 1431.430 1580.120 ;
        RECT 1430.230 1194.280 1430.510 1194.560 ;
        RECT 1429.770 1193.600 1430.050 1193.880 ;
        RECT 1429.770 910.720 1430.050 911.000 ;
        RECT 1430.690 910.720 1430.970 911.000 ;
        RECT 1429.770 869.240 1430.050 869.520 ;
        RECT 1430.690 869.240 1430.970 869.520 ;
        RECT 1428.850 621.040 1429.130 621.320 ;
        RECT 1429.770 621.040 1430.050 621.320 ;
        RECT 1430.230 283.080 1430.510 283.360 ;
        RECT 1431.150 283.080 1431.430 283.360 ;
      LAYER met3 ;
        RECT 1428.825 1628.410 1429.155 1628.425 ;
        RECT 1429.745 1628.410 1430.075 1628.425 ;
        RECT 1428.825 1628.110 1430.075 1628.410 ;
        RECT 1428.825 1628.095 1429.155 1628.110 ;
        RECT 1429.745 1628.095 1430.075 1628.110 ;
        RECT 1430.205 1580.130 1430.535 1580.145 ;
        RECT 1431.125 1580.130 1431.455 1580.145 ;
        RECT 1430.205 1579.830 1431.455 1580.130 ;
        RECT 1430.205 1579.815 1430.535 1579.830 ;
        RECT 1431.125 1579.815 1431.455 1579.830 ;
        RECT 1430.205 1194.570 1430.535 1194.585 ;
        RECT 1429.990 1194.255 1430.535 1194.570 ;
        RECT 1429.990 1193.905 1430.290 1194.255 ;
        RECT 1429.745 1193.590 1430.290 1193.905 ;
        RECT 1429.745 1193.575 1430.075 1193.590 ;
        RECT 1429.745 911.010 1430.075 911.025 ;
        RECT 1430.665 911.010 1430.995 911.025 ;
        RECT 1429.745 910.710 1430.995 911.010 ;
        RECT 1429.745 910.695 1430.075 910.710 ;
        RECT 1430.665 910.695 1430.995 910.710 ;
        RECT 1429.745 869.530 1430.075 869.545 ;
        RECT 1430.665 869.530 1430.995 869.545 ;
        RECT 1429.745 869.230 1430.995 869.530 ;
        RECT 1429.745 869.215 1430.075 869.230 ;
        RECT 1430.665 869.215 1430.995 869.230 ;
        RECT 1428.825 621.330 1429.155 621.345 ;
        RECT 1429.745 621.330 1430.075 621.345 ;
        RECT 1428.825 621.030 1430.075 621.330 ;
        RECT 1428.825 621.015 1429.155 621.030 ;
        RECT 1429.745 621.015 1430.075 621.030 ;
        RECT 1430.205 283.370 1430.535 283.385 ;
        RECT 1431.125 283.370 1431.455 283.385 ;
        RECT 1430.205 283.070 1431.455 283.370 ;
        RECT 1430.205 283.055 1430.535 283.070 ;
        RECT 1431.125 283.055 1431.455 283.070 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.470 41.380 1352.790 41.440 ;
        RECT 1704.830 41.380 1705.150 41.440 ;
        RECT 1352.470 41.240 1705.150 41.380 ;
        RECT 1352.470 41.180 1352.790 41.240 ;
        RECT 1704.830 41.180 1705.150 41.240 ;
      LAYER via ;
        RECT 1352.500 41.180 1352.760 41.440 ;
        RECT 1704.860 41.180 1705.120 41.440 ;
      LAYER met2 ;
        RECT 1705.705 1700.410 1705.985 1704.000 ;
        RECT 1704.920 1700.270 1705.985 1700.410 ;
        RECT 1704.920 41.470 1705.060 1700.270 ;
        RECT 1705.705 1700.000 1705.985 1700.270 ;
        RECT 1352.500 41.150 1352.760 41.470 ;
        RECT 1704.860 41.150 1705.120 41.470 ;
        RECT 1352.560 2.400 1352.700 41.150 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1370.410 30.840 1370.730 30.900 ;
        RECT 1711.730 30.840 1712.050 30.900 ;
        RECT 1370.410 30.700 1712.050 30.840 ;
        RECT 1370.410 30.640 1370.730 30.700 ;
        RECT 1711.730 30.640 1712.050 30.700 ;
      LAYER via ;
        RECT 1370.440 30.640 1370.700 30.900 ;
        RECT 1711.760 30.640 1712.020 30.900 ;
      LAYER met2 ;
        RECT 1713.065 1700.410 1713.345 1704.000 ;
        RECT 1711.820 1700.270 1713.345 1700.410 ;
        RECT 1711.820 30.930 1711.960 1700.270 ;
        RECT 1713.065 1700.000 1713.345 1700.270 ;
        RECT 1370.440 30.610 1370.700 30.930 ;
        RECT 1711.760 30.610 1712.020 30.930 ;
        RECT 1370.500 2.400 1370.640 30.610 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1452.290 1683.920 1452.610 1683.980 ;
        RECT 1720.470 1683.920 1720.790 1683.980 ;
        RECT 1452.290 1683.780 1720.790 1683.920 ;
        RECT 1452.290 1683.720 1452.610 1683.780 ;
        RECT 1720.470 1683.720 1720.790 1683.780 ;
        RECT 1388.350 15.880 1388.670 15.940 ;
        RECT 1452.290 15.880 1452.610 15.940 ;
        RECT 1388.350 15.740 1452.610 15.880 ;
        RECT 1388.350 15.680 1388.670 15.740 ;
        RECT 1452.290 15.680 1452.610 15.740 ;
      LAYER via ;
        RECT 1452.320 1683.720 1452.580 1683.980 ;
        RECT 1720.500 1683.720 1720.760 1683.980 ;
        RECT 1388.380 15.680 1388.640 15.940 ;
        RECT 1452.320 15.680 1452.580 15.940 ;
      LAYER met2 ;
        RECT 1720.425 1700.000 1720.705 1704.000 ;
        RECT 1720.560 1684.010 1720.700 1700.000 ;
        RECT 1452.320 1683.690 1452.580 1684.010 ;
        RECT 1720.500 1683.690 1720.760 1684.010 ;
        RECT 1452.380 15.970 1452.520 1683.690 ;
        RECT 1388.380 15.650 1388.640 15.970 ;
        RECT 1452.320 15.650 1452.580 15.970 ;
        RECT 1388.440 2.400 1388.580 15.650 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1407.210 1688.000 1407.530 1688.060 ;
        RECT 1726.450 1688.000 1726.770 1688.060 ;
        RECT 1407.210 1687.860 1726.770 1688.000 ;
        RECT 1407.210 1687.800 1407.530 1687.860 ;
        RECT 1726.450 1687.800 1726.770 1687.860 ;
        RECT 1406.290 2.960 1406.610 3.020 ;
        RECT 1407.210 2.960 1407.530 3.020 ;
        RECT 1406.290 2.820 1407.530 2.960 ;
        RECT 1406.290 2.760 1406.610 2.820 ;
        RECT 1407.210 2.760 1407.530 2.820 ;
      LAYER via ;
        RECT 1407.240 1687.800 1407.500 1688.060 ;
        RECT 1726.480 1687.800 1726.740 1688.060 ;
        RECT 1406.320 2.760 1406.580 3.020 ;
        RECT 1407.240 2.760 1407.500 3.020 ;
      LAYER met2 ;
        RECT 1727.785 1700.410 1728.065 1704.000 ;
        RECT 1726.540 1700.270 1728.065 1700.410 ;
        RECT 1726.540 1688.090 1726.680 1700.270 ;
        RECT 1727.785 1700.000 1728.065 1700.270 ;
        RECT 1407.240 1687.770 1407.500 1688.090 ;
        RECT 1726.480 1687.770 1726.740 1688.090 ;
        RECT 1407.300 3.050 1407.440 1687.770 ;
        RECT 1406.320 2.730 1406.580 3.050 ;
        RECT 1407.240 2.730 1407.500 3.050 ;
        RECT 1406.380 2.400 1406.520 2.730 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1427.910 1688.340 1428.230 1688.400 ;
        RECT 1735.190 1688.340 1735.510 1688.400 ;
        RECT 1427.910 1688.200 1735.510 1688.340 ;
        RECT 1427.910 1688.140 1428.230 1688.200 ;
        RECT 1735.190 1688.140 1735.510 1688.200 ;
        RECT 1423.770 20.640 1424.090 20.700 ;
        RECT 1427.910 20.640 1428.230 20.700 ;
        RECT 1423.770 20.500 1428.230 20.640 ;
        RECT 1423.770 20.440 1424.090 20.500 ;
        RECT 1427.910 20.440 1428.230 20.500 ;
      LAYER via ;
        RECT 1427.940 1688.140 1428.200 1688.400 ;
        RECT 1735.220 1688.140 1735.480 1688.400 ;
        RECT 1423.800 20.440 1424.060 20.700 ;
        RECT 1427.940 20.440 1428.200 20.700 ;
      LAYER met2 ;
        RECT 1735.145 1700.000 1735.425 1704.000 ;
        RECT 1735.280 1688.430 1735.420 1700.000 ;
        RECT 1427.940 1688.110 1428.200 1688.430 ;
        RECT 1735.220 1688.110 1735.480 1688.430 ;
        RECT 1428.000 20.730 1428.140 1688.110 ;
        RECT 1423.800 20.410 1424.060 20.730 ;
        RECT 1427.940 20.410 1428.200 20.730 ;
        RECT 1423.860 2.400 1424.000 20.410 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1732.045 1688.525 1732.215 1693.455 ;
      LAYER mcon ;
        RECT 1732.045 1693.285 1732.215 1693.455 ;
      LAYER met1 ;
        RECT 1731.985 1693.440 1732.275 1693.485 ;
        RECT 1742.550 1693.440 1742.870 1693.500 ;
        RECT 1731.985 1693.300 1742.870 1693.440 ;
        RECT 1731.985 1693.255 1732.275 1693.300 ;
        RECT 1742.550 1693.240 1742.870 1693.300 ;
        RECT 1441.250 1689.020 1441.570 1689.080 ;
        RECT 1441.250 1688.880 1510.480 1689.020 ;
        RECT 1441.250 1688.820 1441.570 1688.880 ;
        RECT 1510.340 1688.680 1510.480 1688.880 ;
        RECT 1635.830 1688.680 1636.150 1688.740 ;
        RECT 1510.340 1688.540 1636.150 1688.680 ;
        RECT 1635.830 1688.480 1636.150 1688.540 ;
        RECT 1680.910 1688.680 1681.230 1688.740 ;
        RECT 1731.985 1688.680 1732.275 1688.725 ;
        RECT 1680.910 1688.540 1732.275 1688.680 ;
        RECT 1680.910 1688.480 1681.230 1688.540 ;
        RECT 1731.985 1688.495 1732.275 1688.540 ;
      LAYER via ;
        RECT 1742.580 1693.240 1742.840 1693.500 ;
        RECT 1441.280 1688.820 1441.540 1689.080 ;
        RECT 1635.860 1688.480 1636.120 1688.740 ;
        RECT 1680.940 1688.480 1681.200 1688.740 ;
      LAYER met2 ;
        RECT 1742.505 1700.000 1742.785 1704.000 ;
        RECT 1742.640 1693.530 1742.780 1700.000 ;
        RECT 1742.580 1693.210 1742.840 1693.530 ;
        RECT 1441.280 1688.790 1441.540 1689.110 ;
        RECT 1441.340 3.130 1441.480 1688.790 ;
        RECT 1635.850 1688.595 1636.130 1688.965 ;
        RECT 1680.930 1688.595 1681.210 1688.965 ;
        RECT 1635.860 1688.450 1636.120 1688.595 ;
        RECT 1680.940 1688.450 1681.200 1688.595 ;
        RECT 1441.340 2.990 1441.940 3.130 ;
        RECT 1441.800 2.400 1441.940 2.990 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
      LAYER via2 ;
        RECT 1635.850 1688.640 1636.130 1688.920 ;
        RECT 1680.930 1688.640 1681.210 1688.920 ;
      LAYER met3 ;
        RECT 1635.825 1688.930 1636.155 1688.945 ;
        RECT 1680.905 1688.930 1681.235 1688.945 ;
        RECT 1635.825 1688.630 1681.235 1688.930 ;
        RECT 1635.825 1688.615 1636.155 1688.630 ;
        RECT 1680.905 1688.615 1681.235 1688.630 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1708.585 1685.465 1708.755 1687.675 ;
        RECT 1714.105 1687.505 1714.275 1690.735 ;
        RECT 1723.305 1689.205 1723.475 1690.735 ;
      LAYER mcon ;
        RECT 1714.105 1690.565 1714.275 1690.735 ;
        RECT 1723.305 1690.565 1723.475 1690.735 ;
        RECT 1708.585 1687.505 1708.755 1687.675 ;
      LAYER met1 ;
        RECT 1714.045 1690.720 1714.335 1690.765 ;
        RECT 1723.245 1690.720 1723.535 1690.765 ;
        RECT 1714.045 1690.580 1723.535 1690.720 ;
        RECT 1714.045 1690.535 1714.335 1690.580 ;
        RECT 1723.245 1690.535 1723.535 1690.580 ;
        RECT 1723.245 1689.360 1723.535 1689.405 ;
        RECT 1749.910 1689.360 1750.230 1689.420 ;
        RECT 1723.245 1689.220 1750.230 1689.360 ;
        RECT 1723.245 1689.175 1723.535 1689.220 ;
        RECT 1749.910 1689.160 1750.230 1689.220 ;
        RECT 1708.525 1687.660 1708.815 1687.705 ;
        RECT 1714.045 1687.660 1714.335 1687.705 ;
        RECT 1708.525 1687.520 1714.335 1687.660 ;
        RECT 1708.525 1687.475 1708.815 1687.520 ;
        RECT 1714.045 1687.475 1714.335 1687.520 ;
        RECT 1583.390 1685.620 1583.710 1685.680 ;
        RECT 1708.525 1685.620 1708.815 1685.665 ;
        RECT 1583.390 1685.480 1708.815 1685.620 ;
        RECT 1583.390 1685.420 1583.710 1685.480 ;
        RECT 1708.525 1685.435 1708.815 1685.480 ;
        RECT 1459.650 16.220 1459.970 16.280 ;
        RECT 1583.390 16.220 1583.710 16.280 ;
        RECT 1459.650 16.080 1583.710 16.220 ;
        RECT 1459.650 16.020 1459.970 16.080 ;
        RECT 1583.390 16.020 1583.710 16.080 ;
      LAYER via ;
        RECT 1749.940 1689.160 1750.200 1689.420 ;
        RECT 1583.420 1685.420 1583.680 1685.680 ;
        RECT 1459.680 16.020 1459.940 16.280 ;
        RECT 1583.420 16.020 1583.680 16.280 ;
      LAYER met2 ;
        RECT 1749.865 1700.000 1750.145 1704.000 ;
        RECT 1750.000 1689.450 1750.140 1700.000 ;
        RECT 1749.940 1689.130 1750.200 1689.450 ;
        RECT 1583.420 1685.390 1583.680 1685.710 ;
        RECT 1583.480 16.310 1583.620 1685.390 ;
        RECT 1459.680 15.990 1459.940 16.310 ;
        RECT 1583.420 15.990 1583.680 16.310 ;
        RECT 1459.740 2.400 1459.880 15.990 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1727.905 1684.785 1728.075 1688.015 ;
      LAYER mcon ;
        RECT 1727.905 1687.845 1728.075 1688.015 ;
      LAYER met1 ;
        RECT 1727.845 1688.000 1728.135 1688.045 ;
        RECT 1757.270 1688.000 1757.590 1688.060 ;
        RECT 1727.845 1687.860 1757.590 1688.000 ;
        RECT 1727.845 1687.815 1728.135 1687.860 ;
        RECT 1757.270 1687.800 1757.590 1687.860 ;
        RECT 1597.190 1684.940 1597.510 1685.000 ;
        RECT 1727.845 1684.940 1728.135 1684.985 ;
        RECT 1597.190 1684.800 1728.135 1684.940 ;
        RECT 1597.190 1684.740 1597.510 1684.800 ;
        RECT 1727.845 1684.755 1728.135 1684.800 ;
        RECT 1477.590 15.540 1477.910 15.600 ;
        RECT 1597.190 15.540 1597.510 15.600 ;
        RECT 1477.590 15.400 1597.510 15.540 ;
        RECT 1477.590 15.340 1477.910 15.400 ;
        RECT 1597.190 15.340 1597.510 15.400 ;
      LAYER via ;
        RECT 1757.300 1687.800 1757.560 1688.060 ;
        RECT 1597.220 1684.740 1597.480 1685.000 ;
        RECT 1477.620 15.340 1477.880 15.600 ;
        RECT 1597.220 15.340 1597.480 15.600 ;
      LAYER met2 ;
        RECT 1757.225 1700.000 1757.505 1704.000 ;
        RECT 1757.360 1688.090 1757.500 1700.000 ;
        RECT 1757.300 1687.770 1757.560 1688.090 ;
        RECT 1597.220 1684.710 1597.480 1685.030 ;
        RECT 1597.280 15.630 1597.420 1684.710 ;
        RECT 1477.620 15.310 1477.880 15.630 ;
        RECT 1597.220 15.310 1597.480 15.630 ;
        RECT 1477.680 2.400 1477.820 15.310 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1635.905 1689.545 1636.535 1689.715 ;
      LAYER mcon ;
        RECT 1636.365 1689.545 1636.535 1689.715 ;
      LAYER met1 ;
        RECT 1515.770 1689.700 1516.090 1689.760 ;
        RECT 1635.845 1689.700 1636.135 1689.745 ;
        RECT 1515.770 1689.560 1636.135 1689.700 ;
        RECT 1515.770 1689.500 1516.090 1689.560 ;
        RECT 1635.845 1689.515 1636.135 1689.560 ;
        RECT 1636.305 1689.700 1636.595 1689.745 ;
        RECT 1764.630 1689.700 1764.950 1689.760 ;
        RECT 1636.305 1689.560 1764.950 1689.700 ;
        RECT 1636.305 1689.515 1636.595 1689.560 ;
        RECT 1764.630 1689.500 1764.950 1689.560 ;
        RECT 1495.530 16.900 1495.850 16.960 ;
        RECT 1514.390 16.900 1514.710 16.960 ;
        RECT 1495.530 16.760 1514.710 16.900 ;
        RECT 1495.530 16.700 1495.850 16.760 ;
        RECT 1514.390 16.700 1514.710 16.760 ;
      LAYER via ;
        RECT 1515.800 1689.500 1516.060 1689.760 ;
        RECT 1764.660 1689.500 1764.920 1689.760 ;
        RECT 1495.560 16.700 1495.820 16.960 ;
        RECT 1514.420 16.700 1514.680 16.960 ;
      LAYER met2 ;
        RECT 1764.585 1700.000 1764.865 1704.000 ;
        RECT 1764.720 1689.790 1764.860 1700.000 ;
        RECT 1515.800 1689.470 1516.060 1689.790 ;
        RECT 1764.660 1689.470 1764.920 1689.790 ;
        RECT 1515.860 1673.210 1516.000 1689.470 ;
        RECT 1514.480 1673.070 1516.000 1673.210 ;
        RECT 1514.480 16.990 1514.620 1673.070 ;
        RECT 1495.560 16.670 1495.820 16.990 ;
        RECT 1514.420 16.670 1514.680 16.990 ;
        RECT 1495.620 2.400 1495.760 16.670 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1548.890 1690.380 1549.210 1690.440 ;
        RECT 1771.990 1690.380 1772.310 1690.440 ;
        RECT 1548.890 1690.240 1772.310 1690.380 ;
        RECT 1548.890 1690.180 1549.210 1690.240 ;
        RECT 1771.990 1690.180 1772.310 1690.240 ;
        RECT 1513.010 20.300 1513.330 20.360 ;
        RECT 1548.890 20.300 1549.210 20.360 ;
        RECT 1513.010 20.160 1549.210 20.300 ;
        RECT 1513.010 20.100 1513.330 20.160 ;
        RECT 1548.890 20.100 1549.210 20.160 ;
      LAYER via ;
        RECT 1548.920 1690.180 1549.180 1690.440 ;
        RECT 1772.020 1690.180 1772.280 1690.440 ;
        RECT 1513.040 20.100 1513.300 20.360 ;
        RECT 1548.920 20.100 1549.180 20.360 ;
      LAYER met2 ;
        RECT 1771.945 1700.000 1772.225 1704.000 ;
        RECT 1772.080 1690.470 1772.220 1700.000 ;
        RECT 1548.920 1690.150 1549.180 1690.470 ;
        RECT 1772.020 1690.150 1772.280 1690.470 ;
        RECT 1548.980 20.390 1549.120 1690.150 ;
        RECT 1513.040 20.070 1513.300 20.390 ;
        RECT 1548.920 20.070 1549.180 20.390 ;
        RECT 1513.100 2.400 1513.240 20.070 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1435.270 1678.140 1435.590 1678.200 ;
        RECT 1439.870 1678.140 1440.190 1678.200 ;
        RECT 1435.270 1678.000 1440.190 1678.140 ;
        RECT 1435.270 1677.940 1435.590 1678.000 ;
        RECT 1439.870 1677.940 1440.190 1678.000 ;
        RECT 709.850 36.960 710.170 37.020 ;
        RECT 1435.270 36.960 1435.590 37.020 ;
        RECT 709.850 36.820 1435.590 36.960 ;
        RECT 709.850 36.760 710.170 36.820 ;
        RECT 1435.270 36.760 1435.590 36.820 ;
      LAYER via ;
        RECT 1435.300 1677.940 1435.560 1678.200 ;
        RECT 1439.900 1677.940 1440.160 1678.200 ;
        RECT 709.880 36.760 710.140 37.020 ;
        RECT 1435.300 36.760 1435.560 37.020 ;
      LAYER met2 ;
        RECT 1441.205 1700.410 1441.485 1704.000 ;
        RECT 1439.960 1700.270 1441.485 1700.410 ;
        RECT 1439.960 1678.230 1440.100 1700.270 ;
        RECT 1441.205 1700.000 1441.485 1700.270 ;
        RECT 1435.300 1677.910 1435.560 1678.230 ;
        RECT 1439.900 1677.910 1440.160 1678.230 ;
        RECT 1435.360 37.050 1435.500 1677.910 ;
        RECT 709.880 36.730 710.140 37.050 ;
        RECT 1435.300 36.730 1435.560 37.050 ;
        RECT 709.940 17.410 710.080 36.730 ;
        RECT 709.940 17.270 710.540 17.410 ;
        RECT 710.400 2.400 710.540 17.270 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1530.950 1690.040 1531.270 1690.100 ;
        RECT 1779.350 1690.040 1779.670 1690.100 ;
        RECT 1530.950 1689.900 1779.670 1690.040 ;
        RECT 1530.950 1689.840 1531.270 1689.900 ;
        RECT 1779.350 1689.840 1779.670 1689.900 ;
      LAYER via ;
        RECT 1530.980 1689.840 1531.240 1690.100 ;
        RECT 1779.380 1689.840 1779.640 1690.100 ;
      LAYER met2 ;
        RECT 1779.305 1700.000 1779.585 1704.000 ;
        RECT 1779.440 1690.130 1779.580 1700.000 ;
        RECT 1530.980 1689.810 1531.240 1690.130 ;
        RECT 1779.380 1689.810 1779.640 1690.130 ;
        RECT 1531.040 2.400 1531.180 1689.810 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1752.745 1684.105 1752.915 1686.315 ;
        RECT 1769.765 1686.145 1769.935 1687.675 ;
        RECT 1679.145 14.705 1679.315 15.895 ;
      LAYER mcon ;
        RECT 1769.765 1687.505 1769.935 1687.675 ;
        RECT 1752.745 1686.145 1752.915 1686.315 ;
        RECT 1679.145 15.725 1679.315 15.895 ;
      LAYER met1 ;
        RECT 1769.705 1687.660 1769.995 1687.705 ;
        RECT 1786.710 1687.660 1787.030 1687.720 ;
        RECT 1769.705 1687.520 1787.030 1687.660 ;
        RECT 1769.705 1687.475 1769.995 1687.520 ;
        RECT 1786.710 1687.460 1787.030 1687.520 ;
        RECT 1752.685 1686.300 1752.975 1686.345 ;
        RECT 1769.705 1686.300 1769.995 1686.345 ;
        RECT 1752.685 1686.160 1769.995 1686.300 ;
        RECT 1752.685 1686.115 1752.975 1686.160 ;
        RECT 1769.705 1686.115 1769.995 1686.160 ;
        RECT 1721.390 1684.260 1721.710 1684.320 ;
        RECT 1752.685 1684.260 1752.975 1684.305 ;
        RECT 1721.390 1684.120 1752.975 1684.260 ;
        RECT 1721.390 1684.060 1721.710 1684.120 ;
        RECT 1752.685 1684.075 1752.975 1684.120 ;
        RECT 1548.890 15.880 1549.210 15.940 ;
        RECT 1679.085 15.880 1679.375 15.925 ;
        RECT 1548.890 15.740 1679.375 15.880 ;
        RECT 1548.890 15.680 1549.210 15.740 ;
        RECT 1679.085 15.695 1679.375 15.740 ;
        RECT 1679.085 14.860 1679.375 14.905 ;
        RECT 1721.850 14.860 1722.170 14.920 ;
        RECT 1679.085 14.720 1722.170 14.860 ;
        RECT 1679.085 14.675 1679.375 14.720 ;
        RECT 1721.850 14.660 1722.170 14.720 ;
      LAYER via ;
        RECT 1786.740 1687.460 1787.000 1687.720 ;
        RECT 1721.420 1684.060 1721.680 1684.320 ;
        RECT 1548.920 15.680 1549.180 15.940 ;
        RECT 1721.880 14.660 1722.140 14.920 ;
      LAYER met2 ;
        RECT 1786.665 1700.000 1786.945 1704.000 ;
        RECT 1786.800 1687.750 1786.940 1700.000 ;
        RECT 1786.740 1687.430 1787.000 1687.750 ;
        RECT 1721.420 1684.030 1721.680 1684.350 ;
        RECT 1548.920 15.650 1549.180 15.970 ;
        RECT 1548.980 2.400 1549.120 15.650 ;
        RECT 1721.480 15.370 1721.620 1684.030 ;
        RECT 1721.480 15.230 1722.080 15.370 ;
        RECT 1721.940 14.950 1722.080 15.230 ;
        RECT 1721.880 14.630 1722.140 14.950 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1761.945 19.805 1762.115 20.655 ;
      LAYER mcon ;
        RECT 1761.945 20.485 1762.115 20.655 ;
      LAYER met1 ;
        RECT 1761.885 20.640 1762.175 20.685 ;
        RECT 1794.530 20.640 1794.850 20.700 ;
        RECT 1761.885 20.500 1794.850 20.640 ;
        RECT 1761.885 20.455 1762.175 20.500 ;
        RECT 1794.530 20.440 1794.850 20.500 ;
        RECT 1566.830 19.960 1567.150 20.020 ;
        RECT 1761.885 19.960 1762.175 20.005 ;
        RECT 1566.830 19.820 1762.175 19.960 ;
        RECT 1566.830 19.760 1567.150 19.820 ;
        RECT 1761.885 19.775 1762.175 19.820 ;
      LAYER via ;
        RECT 1794.560 20.440 1794.820 20.700 ;
        RECT 1566.860 19.760 1567.120 20.020 ;
      LAYER met2 ;
        RECT 1794.025 1700.410 1794.305 1704.000 ;
        RECT 1794.025 1700.270 1794.760 1700.410 ;
        RECT 1794.025 1700.000 1794.305 1700.270 ;
        RECT 1794.620 20.730 1794.760 1700.270 ;
        RECT 1794.560 20.410 1794.820 20.730 ;
        RECT 1566.860 19.730 1567.120 20.050 ;
        RECT 1566.920 2.400 1567.060 19.730 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1703.985 20.485 1704.615 20.655 ;
        RECT 1678.225 14.025 1678.395 14.875 ;
        RECT 1703.985 14.025 1704.155 20.485 ;
      LAYER mcon ;
        RECT 1704.445 20.485 1704.615 20.655 ;
        RECT 1678.225 14.705 1678.395 14.875 ;
      LAYER met1 ;
        RECT 1728.290 1684.600 1728.610 1684.660 ;
        RECT 1801.430 1684.600 1801.750 1684.660 ;
        RECT 1728.290 1684.460 1801.750 1684.600 ;
        RECT 1728.290 1684.400 1728.610 1684.460 ;
        RECT 1801.430 1684.400 1801.750 1684.460 ;
        RECT 1704.385 20.640 1704.675 20.685 ;
        RECT 1728.290 20.640 1728.610 20.700 ;
        RECT 1704.385 20.500 1728.610 20.640 ;
        RECT 1704.385 20.455 1704.675 20.500 ;
        RECT 1728.290 20.440 1728.610 20.500 ;
        RECT 1584.770 14.860 1585.090 14.920 ;
        RECT 1678.165 14.860 1678.455 14.905 ;
        RECT 1584.770 14.720 1678.455 14.860 ;
        RECT 1584.770 14.660 1585.090 14.720 ;
        RECT 1678.165 14.675 1678.455 14.720 ;
        RECT 1678.165 14.180 1678.455 14.225 ;
        RECT 1703.925 14.180 1704.215 14.225 ;
        RECT 1678.165 14.040 1704.215 14.180 ;
        RECT 1678.165 13.995 1678.455 14.040 ;
        RECT 1703.925 13.995 1704.215 14.040 ;
      LAYER via ;
        RECT 1728.320 1684.400 1728.580 1684.660 ;
        RECT 1801.460 1684.400 1801.720 1684.660 ;
        RECT 1728.320 20.440 1728.580 20.700 ;
        RECT 1584.800 14.660 1585.060 14.920 ;
      LAYER met2 ;
        RECT 1801.385 1700.000 1801.665 1704.000 ;
        RECT 1801.520 1684.690 1801.660 1700.000 ;
        RECT 1728.320 1684.370 1728.580 1684.690 ;
        RECT 1801.460 1684.370 1801.720 1684.690 ;
        RECT 1728.380 20.730 1728.520 1684.370 ;
        RECT 1728.320 20.410 1728.580 20.730 ;
        RECT 1584.800 14.630 1585.060 14.950 ;
        RECT 1584.860 2.400 1585.000 14.630 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1607.310 1686.640 1607.630 1686.700 ;
        RECT 1808.790 1686.640 1809.110 1686.700 ;
        RECT 1607.310 1686.500 1809.110 1686.640 ;
        RECT 1607.310 1686.440 1607.630 1686.500 ;
        RECT 1808.790 1686.440 1809.110 1686.500 ;
        RECT 1602.250 17.580 1602.570 17.640 ;
        RECT 1605.930 17.580 1606.250 17.640 ;
        RECT 1602.250 17.440 1606.250 17.580 ;
        RECT 1602.250 17.380 1602.570 17.440 ;
        RECT 1605.930 17.380 1606.250 17.440 ;
      LAYER via ;
        RECT 1607.340 1686.440 1607.600 1686.700 ;
        RECT 1808.820 1686.440 1809.080 1686.700 ;
        RECT 1602.280 17.380 1602.540 17.640 ;
        RECT 1605.960 17.380 1606.220 17.640 ;
      LAYER met2 ;
        RECT 1808.745 1700.000 1809.025 1704.000 ;
        RECT 1808.880 1686.730 1809.020 1700.000 ;
        RECT 1607.340 1686.410 1607.600 1686.730 ;
        RECT 1808.820 1686.410 1809.080 1686.730 ;
        RECT 1607.400 24.040 1607.540 1686.410 ;
        RECT 1606.020 23.900 1607.540 24.040 ;
        RECT 1606.020 17.670 1606.160 23.900 ;
        RECT 1602.280 17.350 1602.540 17.670 ;
        RECT 1605.960 17.350 1606.220 17.670 ;
        RECT 1602.340 2.400 1602.480 17.350 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1815.690 17.580 1816.010 17.640 ;
        RECT 1776.680 17.440 1816.010 17.580 ;
        RECT 1620.190 17.240 1620.510 17.300 ;
        RECT 1776.680 17.240 1776.820 17.440 ;
        RECT 1815.690 17.380 1816.010 17.440 ;
        RECT 1620.190 17.100 1776.820 17.240 ;
        RECT 1620.190 17.040 1620.510 17.100 ;
      LAYER via ;
        RECT 1620.220 17.040 1620.480 17.300 ;
        RECT 1815.720 17.380 1815.980 17.640 ;
      LAYER met2 ;
        RECT 1816.105 1700.410 1816.385 1704.000 ;
        RECT 1815.780 1700.270 1816.385 1700.410 ;
        RECT 1815.780 17.670 1815.920 1700.270 ;
        RECT 1816.105 1700.000 1816.385 1700.270 ;
        RECT 1815.720 17.350 1815.980 17.670 ;
        RECT 1620.220 17.010 1620.480 17.330 ;
        RECT 1620.280 2.400 1620.420 17.010 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1678.685 15.045 1678.855 17.935 ;
        RECT 1777.125 17.085 1777.295 18.275 ;
      LAYER mcon ;
        RECT 1777.125 18.105 1777.295 18.275 ;
        RECT 1678.685 17.765 1678.855 17.935 ;
      LAYER met1 ;
        RECT 1817.990 1683.920 1818.310 1683.980 ;
        RECT 1823.510 1683.920 1823.830 1683.980 ;
        RECT 1817.990 1683.780 1823.830 1683.920 ;
        RECT 1817.990 1683.720 1818.310 1683.780 ;
        RECT 1823.510 1683.720 1823.830 1683.780 ;
        RECT 1777.065 18.260 1777.355 18.305 ;
        RECT 1775.760 18.120 1777.355 18.260 ;
        RECT 1678.625 17.920 1678.915 17.965 ;
        RECT 1775.760 17.920 1775.900 18.120 ;
        RECT 1777.065 18.075 1777.355 18.120 ;
        RECT 1678.625 17.780 1775.900 17.920 ;
        RECT 1678.625 17.735 1678.915 17.780 ;
        RECT 1777.065 17.240 1777.355 17.285 ;
        RECT 1817.990 17.240 1818.310 17.300 ;
        RECT 1777.065 17.100 1818.310 17.240 ;
        RECT 1777.065 17.055 1777.355 17.100 ;
        RECT 1817.990 17.040 1818.310 17.100 ;
        RECT 1638.130 15.200 1638.450 15.260 ;
        RECT 1678.625 15.200 1678.915 15.245 ;
        RECT 1638.130 15.060 1678.915 15.200 ;
        RECT 1638.130 15.000 1638.450 15.060 ;
        RECT 1678.625 15.015 1678.915 15.060 ;
      LAYER via ;
        RECT 1818.020 1683.720 1818.280 1683.980 ;
        RECT 1823.540 1683.720 1823.800 1683.980 ;
        RECT 1818.020 17.040 1818.280 17.300 ;
        RECT 1638.160 15.000 1638.420 15.260 ;
      LAYER met2 ;
        RECT 1823.465 1700.000 1823.745 1704.000 ;
        RECT 1823.600 1684.010 1823.740 1700.000 ;
        RECT 1818.020 1683.690 1818.280 1684.010 ;
        RECT 1823.540 1683.690 1823.800 1684.010 ;
        RECT 1818.080 17.330 1818.220 1683.690 ;
        RECT 1818.020 17.010 1818.280 17.330 ;
        RECT 1638.160 14.970 1638.420 15.290 ;
        RECT 1638.220 2.400 1638.360 14.970 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1679.605 18.445 1679.775 19.635 ;
      LAYER mcon ;
        RECT 1679.605 19.465 1679.775 19.635 ;
      LAYER met1 ;
        RECT 1679.545 19.620 1679.835 19.665 ;
        RECT 1829.030 19.620 1829.350 19.680 ;
        RECT 1679.545 19.480 1829.350 19.620 ;
        RECT 1679.545 19.435 1679.835 19.480 ;
        RECT 1829.030 19.420 1829.350 19.480 ;
        RECT 1656.070 18.600 1656.390 18.660 ;
        RECT 1679.545 18.600 1679.835 18.645 ;
        RECT 1656.070 18.460 1679.835 18.600 ;
        RECT 1656.070 18.400 1656.390 18.460 ;
        RECT 1679.545 18.415 1679.835 18.460 ;
      LAYER via ;
        RECT 1829.060 19.420 1829.320 19.680 ;
        RECT 1656.100 18.400 1656.360 18.660 ;
      LAYER met2 ;
        RECT 1830.825 1700.410 1831.105 1704.000 ;
        RECT 1829.120 1700.270 1831.105 1700.410 ;
        RECT 1829.120 19.710 1829.260 1700.270 ;
        RECT 1830.825 1700.000 1831.105 1700.270 ;
        RECT 1829.060 19.390 1829.320 19.710 ;
        RECT 1656.100 18.370 1656.360 18.690 ;
        RECT 1656.160 2.400 1656.300 18.370 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1676.310 1685.280 1676.630 1685.340 ;
        RECT 1838.230 1685.280 1838.550 1685.340 ;
        RECT 1676.310 1685.140 1838.550 1685.280 ;
        RECT 1676.310 1685.080 1676.630 1685.140 ;
        RECT 1838.230 1685.080 1838.550 1685.140 ;
        RECT 1673.550 20.640 1673.870 20.700 ;
        RECT 1676.310 20.640 1676.630 20.700 ;
        RECT 1673.550 20.500 1676.630 20.640 ;
        RECT 1673.550 20.440 1673.870 20.500 ;
        RECT 1676.310 20.440 1676.630 20.500 ;
      LAYER via ;
        RECT 1676.340 1685.080 1676.600 1685.340 ;
        RECT 1838.260 1685.080 1838.520 1685.340 ;
        RECT 1673.580 20.440 1673.840 20.700 ;
        RECT 1676.340 20.440 1676.600 20.700 ;
      LAYER met2 ;
        RECT 1838.185 1700.000 1838.465 1704.000 ;
        RECT 1838.320 1685.370 1838.460 1700.000 ;
        RECT 1676.340 1685.050 1676.600 1685.370 ;
        RECT 1838.260 1685.050 1838.520 1685.370 ;
        RECT 1676.400 20.730 1676.540 1685.050 ;
        RECT 1673.580 20.410 1673.840 20.730 ;
        RECT 1676.340 20.410 1676.600 20.730 ;
        RECT 1673.640 2.400 1673.780 20.410 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1691.490 18.600 1691.810 18.660 ;
        RECT 1843.290 18.600 1843.610 18.660 ;
        RECT 1691.490 18.460 1843.610 18.600 ;
        RECT 1691.490 18.400 1691.810 18.460 ;
        RECT 1843.290 18.400 1843.610 18.460 ;
      LAYER via ;
        RECT 1691.520 18.400 1691.780 18.660 ;
        RECT 1843.320 18.400 1843.580 18.660 ;
      LAYER met2 ;
        RECT 1845.545 1700.410 1845.825 1704.000 ;
        RECT 1843.380 1700.270 1845.825 1700.410 ;
        RECT 1843.380 18.690 1843.520 1700.270 ;
        RECT 1845.545 1700.000 1845.825 1700.270 ;
        RECT 1691.520 18.370 1691.780 18.690 ;
        RECT 1843.320 18.370 1843.580 18.690 ;
        RECT 1691.580 2.400 1691.720 18.370 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1442.170 1678.140 1442.490 1678.200 ;
        RECT 1447.230 1678.140 1447.550 1678.200 ;
        RECT 1442.170 1678.000 1447.550 1678.140 ;
        RECT 1442.170 1677.940 1442.490 1678.000 ;
        RECT 1447.230 1677.940 1447.550 1678.000 ;
        RECT 728.250 36.620 728.570 36.680 ;
        RECT 1442.170 36.620 1442.490 36.680 ;
        RECT 728.250 36.480 1442.490 36.620 ;
        RECT 728.250 36.420 728.570 36.480 ;
        RECT 1442.170 36.420 1442.490 36.480 ;
      LAYER via ;
        RECT 1442.200 1677.940 1442.460 1678.200 ;
        RECT 1447.260 1677.940 1447.520 1678.200 ;
        RECT 728.280 36.420 728.540 36.680 ;
        RECT 1442.200 36.420 1442.460 36.680 ;
      LAYER met2 ;
        RECT 1448.565 1700.410 1448.845 1704.000 ;
        RECT 1447.320 1700.270 1448.845 1700.410 ;
        RECT 1447.320 1678.230 1447.460 1700.270 ;
        RECT 1448.565 1700.000 1448.845 1700.270 ;
        RECT 1442.200 1677.910 1442.460 1678.230 ;
        RECT 1447.260 1677.910 1447.520 1678.230 ;
        RECT 1442.260 36.710 1442.400 1677.910 ;
        RECT 728.280 36.390 728.540 36.710 ;
        RECT 1442.200 36.390 1442.460 36.710 ;
        RECT 728.340 2.400 728.480 36.390 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1709.430 18.940 1709.750 19.000 ;
        RECT 1850.650 18.940 1850.970 19.000 ;
        RECT 1709.430 18.800 1850.970 18.940 ;
        RECT 1709.430 18.740 1709.750 18.800 ;
        RECT 1850.650 18.740 1850.970 18.800 ;
      LAYER via ;
        RECT 1709.460 18.740 1709.720 19.000 ;
        RECT 1850.680 18.740 1850.940 19.000 ;
      LAYER met2 ;
        RECT 1852.905 1700.410 1853.185 1704.000 ;
        RECT 1850.740 1700.270 1853.185 1700.410 ;
        RECT 1850.740 19.030 1850.880 1700.270 ;
        RECT 1852.905 1700.000 1853.185 1700.270 ;
        RECT 1709.460 18.710 1709.720 19.030 ;
        RECT 1850.680 18.710 1850.940 19.030 ;
        RECT 1709.520 2.400 1709.660 18.710 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1841.065 1685.805 1841.235 1688.015 ;
        RECT 1745.845 14.705 1746.015 20.655 ;
      LAYER mcon ;
        RECT 1841.065 1687.845 1841.235 1688.015 ;
        RECT 1745.845 20.485 1746.015 20.655 ;
      LAYER met1 ;
        RECT 1758.190 1688.000 1758.510 1688.060 ;
        RECT 1841.005 1688.000 1841.295 1688.045 ;
        RECT 1758.190 1687.860 1841.295 1688.000 ;
        RECT 1758.190 1687.800 1758.510 1687.860 ;
        RECT 1841.005 1687.815 1841.295 1687.860 ;
        RECT 1841.005 1685.960 1841.295 1686.005 ;
        RECT 1860.310 1685.960 1860.630 1686.020 ;
        RECT 1841.005 1685.820 1860.630 1685.960 ;
        RECT 1841.005 1685.775 1841.295 1685.820 ;
        RECT 1860.310 1685.760 1860.630 1685.820 ;
        RECT 1755.890 1684.260 1756.210 1684.320 ;
        RECT 1758.190 1684.260 1758.510 1684.320 ;
        RECT 1755.890 1684.120 1758.510 1684.260 ;
        RECT 1755.890 1684.060 1756.210 1684.120 ;
        RECT 1758.190 1684.060 1758.510 1684.120 ;
        RECT 1745.785 20.640 1746.075 20.685 ;
        RECT 1755.890 20.640 1756.210 20.700 ;
        RECT 1745.785 20.500 1756.210 20.640 ;
        RECT 1745.785 20.455 1746.075 20.500 ;
        RECT 1755.890 20.440 1756.210 20.500 ;
        RECT 1727.370 14.860 1727.690 14.920 ;
        RECT 1745.785 14.860 1746.075 14.905 ;
        RECT 1727.370 14.720 1746.075 14.860 ;
        RECT 1727.370 14.660 1727.690 14.720 ;
        RECT 1745.785 14.675 1746.075 14.720 ;
      LAYER via ;
        RECT 1758.220 1687.800 1758.480 1688.060 ;
        RECT 1860.340 1685.760 1860.600 1686.020 ;
        RECT 1755.920 1684.060 1756.180 1684.320 ;
        RECT 1758.220 1684.060 1758.480 1684.320 ;
        RECT 1755.920 20.440 1756.180 20.700 ;
        RECT 1727.400 14.660 1727.660 14.920 ;
      LAYER met2 ;
        RECT 1860.265 1700.000 1860.545 1704.000 ;
        RECT 1758.220 1687.770 1758.480 1688.090 ;
        RECT 1758.280 1684.350 1758.420 1687.770 ;
        RECT 1860.400 1686.050 1860.540 1700.000 ;
        RECT 1860.340 1685.730 1860.600 1686.050 ;
        RECT 1755.920 1684.030 1756.180 1684.350 ;
        RECT 1758.220 1684.030 1758.480 1684.350 ;
        RECT 1755.980 20.730 1756.120 1684.030 ;
        RECT 1755.920 20.410 1756.180 20.730 ;
        RECT 1727.400 14.630 1727.660 14.950 ;
        RECT 1727.460 2.400 1727.600 14.630 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1863.605 1545.725 1863.775 1593.835 ;
        RECT 1863.605 1449.165 1863.775 1497.275 ;
        RECT 1863.605 1352.605 1863.775 1400.715 ;
        RECT 1863.605 1256.045 1863.775 1304.155 ;
        RECT 1864.065 565.845 1864.235 613.955 ;
        RECT 1863.605 386.325 1863.775 517.055 ;
        RECT 1824.965 15.385 1825.135 16.575 ;
      LAYER mcon ;
        RECT 1863.605 1593.665 1863.775 1593.835 ;
        RECT 1863.605 1497.105 1863.775 1497.275 ;
        RECT 1863.605 1400.545 1863.775 1400.715 ;
        RECT 1863.605 1303.985 1863.775 1304.155 ;
        RECT 1864.065 613.785 1864.235 613.955 ;
        RECT 1863.605 516.885 1863.775 517.055 ;
        RECT 1824.965 16.405 1825.135 16.575 ;
      LAYER met1 ;
        RECT 1863.530 1642.440 1863.850 1642.500 ;
        RECT 1865.370 1642.440 1865.690 1642.500 ;
        RECT 1863.530 1642.300 1865.690 1642.440 ;
        RECT 1863.530 1642.240 1863.850 1642.300 ;
        RECT 1865.370 1642.240 1865.690 1642.300 ;
        RECT 1863.530 1593.820 1863.850 1593.880 ;
        RECT 1863.335 1593.680 1863.850 1593.820 ;
        RECT 1863.530 1593.620 1863.850 1593.680 ;
        RECT 1863.530 1545.880 1863.850 1545.940 ;
        RECT 1863.335 1545.740 1863.850 1545.880 ;
        RECT 1863.530 1545.680 1863.850 1545.740 ;
        RECT 1863.530 1497.260 1863.850 1497.320 ;
        RECT 1863.335 1497.120 1863.850 1497.260 ;
        RECT 1863.530 1497.060 1863.850 1497.120 ;
        RECT 1863.530 1449.320 1863.850 1449.380 ;
        RECT 1863.335 1449.180 1863.850 1449.320 ;
        RECT 1863.530 1449.120 1863.850 1449.180 ;
        RECT 1863.530 1400.700 1863.850 1400.760 ;
        RECT 1863.335 1400.560 1863.850 1400.700 ;
        RECT 1863.530 1400.500 1863.850 1400.560 ;
        RECT 1863.530 1352.760 1863.850 1352.820 ;
        RECT 1863.335 1352.620 1863.850 1352.760 ;
        RECT 1863.530 1352.560 1863.850 1352.620 ;
        RECT 1863.530 1304.140 1863.850 1304.200 ;
        RECT 1863.335 1304.000 1863.850 1304.140 ;
        RECT 1863.530 1303.940 1863.850 1304.000 ;
        RECT 1863.530 1256.200 1863.850 1256.260 ;
        RECT 1863.335 1256.060 1863.850 1256.200 ;
        RECT 1863.530 1256.000 1863.850 1256.060 ;
        RECT 1862.610 1159.300 1862.930 1159.360 ;
        RECT 1863.530 1159.300 1863.850 1159.360 ;
        RECT 1862.610 1159.160 1863.850 1159.300 ;
        RECT 1862.610 1159.100 1862.930 1159.160 ;
        RECT 1863.530 1159.100 1863.850 1159.160 ;
        RECT 1862.610 1062.740 1862.930 1062.800 ;
        RECT 1863.530 1062.740 1863.850 1062.800 ;
        RECT 1862.610 1062.600 1863.850 1062.740 ;
        RECT 1862.610 1062.540 1862.930 1062.600 ;
        RECT 1863.530 1062.540 1863.850 1062.600 ;
        RECT 1862.610 966.180 1862.930 966.240 ;
        RECT 1863.530 966.180 1863.850 966.240 ;
        RECT 1862.610 966.040 1863.850 966.180 ;
        RECT 1862.610 965.980 1862.930 966.040 ;
        RECT 1863.530 965.980 1863.850 966.040 ;
        RECT 1863.530 882.200 1863.850 882.260 ;
        RECT 1863.990 882.200 1864.310 882.260 ;
        RECT 1863.530 882.060 1864.310 882.200 ;
        RECT 1863.530 882.000 1863.850 882.060 ;
        RECT 1863.990 882.000 1864.310 882.060 ;
        RECT 1862.610 821.000 1862.930 821.060 ;
        RECT 1863.990 821.000 1864.310 821.060 ;
        RECT 1862.610 820.860 1864.310 821.000 ;
        RECT 1862.610 820.800 1862.930 820.860 ;
        RECT 1863.990 820.800 1864.310 820.860 ;
        RECT 1863.990 613.940 1864.310 614.000 ;
        RECT 1863.795 613.800 1864.310 613.940 ;
        RECT 1863.990 613.740 1864.310 613.800 ;
        RECT 1863.990 566.000 1864.310 566.060 ;
        RECT 1863.795 565.860 1864.310 566.000 ;
        RECT 1863.990 565.800 1864.310 565.860 ;
        RECT 1863.990 517.180 1864.310 517.440 ;
        RECT 1863.545 517.040 1863.835 517.085 ;
        RECT 1864.080 517.040 1864.220 517.180 ;
        RECT 1863.545 516.900 1864.220 517.040 ;
        RECT 1863.545 516.855 1863.835 516.900 ;
        RECT 1863.530 386.480 1863.850 386.540 ;
        RECT 1863.335 386.340 1863.850 386.480 ;
        RECT 1863.530 386.280 1863.850 386.340 ;
        RECT 1863.530 193.020 1863.850 193.080 ;
        RECT 1863.990 193.020 1864.310 193.080 ;
        RECT 1863.530 192.880 1864.310 193.020 ;
        RECT 1863.530 192.820 1863.850 192.880 ;
        RECT 1863.990 192.820 1864.310 192.880 ;
        RECT 1745.310 16.560 1745.630 16.620 ;
        RECT 1824.905 16.560 1825.195 16.605 ;
        RECT 1745.310 16.420 1825.195 16.560 ;
        RECT 1745.310 16.360 1745.630 16.420 ;
        RECT 1824.905 16.375 1825.195 16.420 ;
        RECT 1824.905 15.540 1825.195 15.585 ;
        RECT 1864.910 15.540 1865.230 15.600 ;
        RECT 1824.905 15.400 1865.230 15.540 ;
        RECT 1824.905 15.355 1825.195 15.400 ;
        RECT 1864.910 15.340 1865.230 15.400 ;
      LAYER via ;
        RECT 1863.560 1642.240 1863.820 1642.500 ;
        RECT 1865.400 1642.240 1865.660 1642.500 ;
        RECT 1863.560 1593.620 1863.820 1593.880 ;
        RECT 1863.560 1545.680 1863.820 1545.940 ;
        RECT 1863.560 1497.060 1863.820 1497.320 ;
        RECT 1863.560 1449.120 1863.820 1449.380 ;
        RECT 1863.560 1400.500 1863.820 1400.760 ;
        RECT 1863.560 1352.560 1863.820 1352.820 ;
        RECT 1863.560 1303.940 1863.820 1304.200 ;
        RECT 1863.560 1256.000 1863.820 1256.260 ;
        RECT 1862.640 1159.100 1862.900 1159.360 ;
        RECT 1863.560 1159.100 1863.820 1159.360 ;
        RECT 1862.640 1062.540 1862.900 1062.800 ;
        RECT 1863.560 1062.540 1863.820 1062.800 ;
        RECT 1862.640 965.980 1862.900 966.240 ;
        RECT 1863.560 965.980 1863.820 966.240 ;
        RECT 1863.560 882.000 1863.820 882.260 ;
        RECT 1864.020 882.000 1864.280 882.260 ;
        RECT 1862.640 820.800 1862.900 821.060 ;
        RECT 1864.020 820.800 1864.280 821.060 ;
        RECT 1864.020 613.740 1864.280 614.000 ;
        RECT 1864.020 565.800 1864.280 566.060 ;
        RECT 1864.020 517.180 1864.280 517.440 ;
        RECT 1863.560 386.280 1863.820 386.540 ;
        RECT 1863.560 192.820 1863.820 193.080 ;
        RECT 1864.020 192.820 1864.280 193.080 ;
        RECT 1745.340 16.360 1745.600 16.620 ;
        RECT 1864.940 15.340 1865.200 15.600 ;
      LAYER met2 ;
        RECT 1867.625 1701.090 1867.905 1704.000 ;
        RECT 1865.460 1700.950 1867.905 1701.090 ;
        RECT 1865.460 1642.530 1865.600 1700.950 ;
        RECT 1867.625 1700.000 1867.905 1700.950 ;
        RECT 1863.560 1642.210 1863.820 1642.530 ;
        RECT 1865.400 1642.210 1865.660 1642.530 ;
        RECT 1863.620 1593.910 1863.760 1642.210 ;
        RECT 1863.560 1593.590 1863.820 1593.910 ;
        RECT 1863.560 1545.650 1863.820 1545.970 ;
        RECT 1863.620 1497.350 1863.760 1545.650 ;
        RECT 1863.560 1497.030 1863.820 1497.350 ;
        RECT 1863.560 1449.090 1863.820 1449.410 ;
        RECT 1863.620 1400.790 1863.760 1449.090 ;
        RECT 1863.560 1400.470 1863.820 1400.790 ;
        RECT 1863.560 1352.530 1863.820 1352.850 ;
        RECT 1863.620 1304.230 1863.760 1352.530 ;
        RECT 1863.560 1303.910 1863.820 1304.230 ;
        RECT 1863.560 1255.970 1863.820 1256.290 ;
        RECT 1863.620 1207.525 1863.760 1255.970 ;
        RECT 1862.630 1207.155 1862.910 1207.525 ;
        RECT 1863.550 1207.155 1863.830 1207.525 ;
        RECT 1862.700 1159.390 1862.840 1207.155 ;
        RECT 1862.640 1159.070 1862.900 1159.390 ;
        RECT 1863.560 1159.070 1863.820 1159.390 ;
        RECT 1863.620 1110.965 1863.760 1159.070 ;
        RECT 1862.630 1110.595 1862.910 1110.965 ;
        RECT 1863.550 1110.595 1863.830 1110.965 ;
        RECT 1862.700 1062.830 1862.840 1110.595 ;
        RECT 1862.640 1062.510 1862.900 1062.830 ;
        RECT 1863.560 1062.510 1863.820 1062.830 ;
        RECT 1863.620 1014.405 1863.760 1062.510 ;
        RECT 1862.630 1014.035 1862.910 1014.405 ;
        RECT 1863.550 1014.035 1863.830 1014.405 ;
        RECT 1862.700 966.270 1862.840 1014.035 ;
        RECT 1862.640 965.950 1862.900 966.270 ;
        RECT 1863.560 965.950 1863.820 966.270 ;
        RECT 1863.620 882.290 1863.760 965.950 ;
        RECT 1863.560 881.970 1863.820 882.290 ;
        RECT 1864.020 881.970 1864.280 882.290 ;
        RECT 1864.080 821.090 1864.220 881.970 ;
        RECT 1862.640 820.770 1862.900 821.090 ;
        RECT 1864.020 820.770 1864.280 821.090 ;
        RECT 1862.700 773.005 1862.840 820.770 ;
        RECT 1862.630 772.635 1862.910 773.005 ;
        RECT 1863.550 772.635 1863.830 773.005 ;
        RECT 1863.620 738.890 1863.760 772.635 ;
        RECT 1863.160 738.750 1863.760 738.890 ;
        RECT 1863.160 738.210 1863.300 738.750 ;
        RECT 1863.160 738.070 1863.760 738.210 ;
        RECT 1863.620 640.290 1863.760 738.070 ;
        RECT 1863.620 640.150 1864.220 640.290 ;
        RECT 1864.080 614.030 1864.220 640.150 ;
        RECT 1864.020 613.710 1864.280 614.030 ;
        RECT 1864.020 565.770 1864.280 566.090 ;
        RECT 1864.080 517.470 1864.220 565.770 ;
        RECT 1864.020 517.150 1864.280 517.470 ;
        RECT 1863.560 386.250 1863.820 386.570 ;
        RECT 1863.620 351.970 1863.760 386.250 ;
        RECT 1863.160 351.830 1863.760 351.970 ;
        RECT 1863.160 351.290 1863.300 351.830 ;
        RECT 1863.160 351.150 1863.760 351.290 ;
        RECT 1863.620 255.410 1863.760 351.150 ;
        RECT 1863.160 255.270 1863.760 255.410 ;
        RECT 1863.160 254.730 1863.300 255.270 ;
        RECT 1863.160 254.590 1863.760 254.730 ;
        RECT 1863.620 193.110 1863.760 254.590 ;
        RECT 1863.560 192.790 1863.820 193.110 ;
        RECT 1864.020 192.790 1864.280 193.110 ;
        RECT 1864.080 109.890 1864.220 192.790 ;
        RECT 1864.080 109.750 1865.140 109.890 ;
        RECT 1745.340 16.330 1745.600 16.650 ;
        RECT 1745.400 2.400 1745.540 16.330 ;
        RECT 1865.000 15.630 1865.140 109.750 ;
        RECT 1864.940 15.310 1865.200 15.630 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
      LAYER via2 ;
        RECT 1862.630 1207.200 1862.910 1207.480 ;
        RECT 1863.550 1207.200 1863.830 1207.480 ;
        RECT 1862.630 1110.640 1862.910 1110.920 ;
        RECT 1863.550 1110.640 1863.830 1110.920 ;
        RECT 1862.630 1014.080 1862.910 1014.360 ;
        RECT 1863.550 1014.080 1863.830 1014.360 ;
        RECT 1862.630 772.680 1862.910 772.960 ;
        RECT 1863.550 772.680 1863.830 772.960 ;
      LAYER met3 ;
        RECT 1862.605 1207.490 1862.935 1207.505 ;
        RECT 1863.525 1207.490 1863.855 1207.505 ;
        RECT 1862.605 1207.190 1863.855 1207.490 ;
        RECT 1862.605 1207.175 1862.935 1207.190 ;
        RECT 1863.525 1207.175 1863.855 1207.190 ;
        RECT 1862.605 1110.930 1862.935 1110.945 ;
        RECT 1863.525 1110.930 1863.855 1110.945 ;
        RECT 1862.605 1110.630 1863.855 1110.930 ;
        RECT 1862.605 1110.615 1862.935 1110.630 ;
        RECT 1863.525 1110.615 1863.855 1110.630 ;
        RECT 1862.605 1014.370 1862.935 1014.385 ;
        RECT 1863.525 1014.370 1863.855 1014.385 ;
        RECT 1862.605 1014.070 1863.855 1014.370 ;
        RECT 1862.605 1014.055 1862.935 1014.070 ;
        RECT 1863.525 1014.055 1863.855 1014.070 ;
        RECT 1862.605 772.970 1862.935 772.985 ;
        RECT 1863.525 772.970 1863.855 772.985 ;
        RECT 1862.605 772.670 1863.855 772.970 ;
        RECT 1862.605 772.655 1862.935 772.670 ;
        RECT 1863.525 772.655 1863.855 772.670 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1780.345 14.705 1780.515 16.235 ;
      LAYER mcon ;
        RECT 1780.345 16.065 1780.515 16.235 ;
      LAYER met1 ;
        RECT 1762.790 16.220 1763.110 16.280 ;
        RECT 1780.285 16.220 1780.575 16.265 ;
        RECT 1762.790 16.080 1780.575 16.220 ;
        RECT 1762.790 16.020 1763.110 16.080 ;
        RECT 1780.285 16.035 1780.575 16.080 ;
        RECT 1801.980 15.060 1822.360 15.200 ;
        RECT 1780.285 14.860 1780.575 14.905 ;
        RECT 1801.980 14.860 1802.120 15.060 ;
        RECT 1780.285 14.720 1802.120 14.860 ;
        RECT 1822.220 14.860 1822.360 15.060 ;
        RECT 1870.430 14.860 1870.750 14.920 ;
        RECT 1822.220 14.720 1870.750 14.860 ;
        RECT 1780.285 14.675 1780.575 14.720 ;
        RECT 1870.430 14.660 1870.750 14.720 ;
      LAYER via ;
        RECT 1762.820 16.020 1763.080 16.280 ;
        RECT 1870.460 14.660 1870.720 14.920 ;
      LAYER met2 ;
        RECT 1874.985 1701.090 1875.265 1704.000 ;
        RECT 1872.820 1700.950 1875.265 1701.090 ;
        RECT 1872.820 1656.210 1872.960 1700.950 ;
        RECT 1874.985 1700.000 1875.265 1700.950 ;
        RECT 1870.520 1656.070 1872.960 1656.210 ;
        RECT 1762.820 15.990 1763.080 16.310 ;
        RECT 1762.880 2.400 1763.020 15.990 ;
        RECT 1870.520 14.950 1870.660 1656.070 ;
        RECT 1870.460 14.630 1870.720 14.950 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1879.245 1352.605 1879.415 1400.715 ;
        RECT 1879.245 1256.045 1879.415 1304.155 ;
        RECT 1879.245 1159.145 1879.415 1207.255 ;
        RECT 1879.245 1062.585 1879.415 1110.695 ;
        RECT 1879.245 966.025 1879.415 1014.135 ;
        RECT 1879.245 772.905 1879.415 821.015 ;
        RECT 1878.785 579.785 1878.955 627.895 ;
        RECT 1879.245 386.325 1879.415 434.775 ;
        RECT 1879.245 104.125 1879.415 137.955 ;
      LAYER mcon ;
        RECT 1879.245 1400.545 1879.415 1400.715 ;
        RECT 1879.245 1303.985 1879.415 1304.155 ;
        RECT 1879.245 1207.085 1879.415 1207.255 ;
        RECT 1879.245 1110.525 1879.415 1110.695 ;
        RECT 1879.245 1013.965 1879.415 1014.135 ;
        RECT 1879.245 820.845 1879.415 821.015 ;
        RECT 1878.785 627.725 1878.955 627.895 ;
        RECT 1879.245 434.605 1879.415 434.775 ;
        RECT 1879.245 137.785 1879.415 137.955 ;
      LAYER met1 ;
        RECT 1879.170 1607.900 1879.490 1608.160 ;
        RECT 1879.260 1607.080 1879.400 1607.900 ;
        RECT 1879.630 1607.080 1879.950 1607.140 ;
        RECT 1879.260 1606.940 1879.950 1607.080 ;
        RECT 1879.630 1606.880 1879.950 1606.940 ;
        RECT 1879.170 1449.320 1879.490 1449.380 ;
        RECT 1879.630 1449.320 1879.950 1449.380 ;
        RECT 1879.170 1449.180 1879.950 1449.320 ;
        RECT 1879.170 1449.120 1879.490 1449.180 ;
        RECT 1879.630 1449.120 1879.950 1449.180 ;
        RECT 1879.170 1400.700 1879.490 1400.760 ;
        RECT 1878.975 1400.560 1879.490 1400.700 ;
        RECT 1879.170 1400.500 1879.490 1400.560 ;
        RECT 1879.170 1352.760 1879.490 1352.820 ;
        RECT 1878.975 1352.620 1879.490 1352.760 ;
        RECT 1879.170 1352.560 1879.490 1352.620 ;
        RECT 1879.170 1304.140 1879.490 1304.200 ;
        RECT 1878.975 1304.000 1879.490 1304.140 ;
        RECT 1879.170 1303.940 1879.490 1304.000 ;
        RECT 1879.170 1256.200 1879.490 1256.260 ;
        RECT 1878.975 1256.060 1879.490 1256.200 ;
        RECT 1879.170 1256.000 1879.490 1256.060 ;
        RECT 1879.170 1207.240 1879.490 1207.300 ;
        RECT 1878.975 1207.100 1879.490 1207.240 ;
        RECT 1879.170 1207.040 1879.490 1207.100 ;
        RECT 1879.170 1159.300 1879.490 1159.360 ;
        RECT 1878.975 1159.160 1879.490 1159.300 ;
        RECT 1879.170 1159.100 1879.490 1159.160 ;
        RECT 1879.170 1110.680 1879.490 1110.740 ;
        RECT 1878.975 1110.540 1879.490 1110.680 ;
        RECT 1879.170 1110.480 1879.490 1110.540 ;
        RECT 1879.170 1062.740 1879.490 1062.800 ;
        RECT 1878.975 1062.600 1879.490 1062.740 ;
        RECT 1879.170 1062.540 1879.490 1062.600 ;
        RECT 1879.170 1014.120 1879.490 1014.180 ;
        RECT 1878.975 1013.980 1879.490 1014.120 ;
        RECT 1879.170 1013.920 1879.490 1013.980 ;
        RECT 1879.170 966.180 1879.490 966.240 ;
        RECT 1878.975 966.040 1879.490 966.180 ;
        RECT 1879.170 965.980 1879.490 966.040 ;
        RECT 1879.170 882.200 1879.490 882.260 ;
        RECT 1879.630 882.200 1879.950 882.260 ;
        RECT 1879.170 882.060 1879.950 882.200 ;
        RECT 1879.170 882.000 1879.490 882.060 ;
        RECT 1879.630 882.000 1879.950 882.060 ;
        RECT 1879.185 821.000 1879.475 821.045 ;
        RECT 1879.630 821.000 1879.950 821.060 ;
        RECT 1879.185 820.860 1879.950 821.000 ;
        RECT 1879.185 820.815 1879.475 820.860 ;
        RECT 1879.630 820.800 1879.950 820.860 ;
        RECT 1879.170 773.060 1879.490 773.120 ;
        RECT 1878.975 772.920 1879.490 773.060 ;
        RECT 1879.170 772.860 1879.490 772.920 ;
        RECT 1879.170 652.020 1879.490 652.080 ;
        RECT 1880.550 652.020 1880.870 652.080 ;
        RECT 1879.170 651.880 1880.870 652.020 ;
        RECT 1879.170 651.820 1879.490 651.880 ;
        RECT 1880.550 651.820 1880.870 651.880 ;
        RECT 1878.725 627.880 1879.015 627.925 ;
        RECT 1879.170 627.880 1879.490 627.940 ;
        RECT 1878.725 627.740 1879.490 627.880 ;
        RECT 1878.725 627.695 1879.015 627.740 ;
        RECT 1879.170 627.680 1879.490 627.740 ;
        RECT 1878.710 579.940 1879.030 580.000 ;
        RECT 1878.515 579.800 1879.030 579.940 ;
        RECT 1878.710 579.740 1879.030 579.800 ;
        RECT 1878.710 545.060 1879.030 545.320 ;
        RECT 1878.800 544.920 1878.940 545.060 ;
        RECT 1879.170 544.920 1879.490 544.980 ;
        RECT 1878.800 544.780 1879.490 544.920 ;
        RECT 1879.170 544.720 1879.490 544.780 ;
        RECT 1879.170 434.760 1879.490 434.820 ;
        RECT 1878.975 434.620 1879.490 434.760 ;
        RECT 1879.170 434.560 1879.490 434.620 ;
        RECT 1879.170 386.480 1879.490 386.540 ;
        RECT 1878.975 386.340 1879.490 386.480 ;
        RECT 1879.170 386.280 1879.490 386.340 ;
        RECT 1879.170 352.280 1879.490 352.540 ;
        RECT 1879.260 351.860 1879.400 352.280 ;
        RECT 1879.170 351.600 1879.490 351.860 ;
        RECT 1879.170 255.720 1879.490 255.980 ;
        RECT 1879.260 255.300 1879.400 255.720 ;
        RECT 1879.170 255.040 1879.490 255.300 ;
        RECT 1878.710 234.500 1879.030 234.560 ;
        RECT 1879.170 234.500 1879.490 234.560 ;
        RECT 1878.710 234.360 1879.490 234.500 ;
        RECT 1878.710 234.300 1879.030 234.360 ;
        RECT 1879.170 234.300 1879.490 234.360 ;
        RECT 1878.710 145.080 1879.030 145.140 ;
        RECT 1879.170 145.080 1879.490 145.140 ;
        RECT 1878.710 144.940 1879.490 145.080 ;
        RECT 1878.710 144.880 1879.030 144.940 ;
        RECT 1879.170 144.880 1879.490 144.940 ;
        RECT 1879.170 137.940 1879.490 138.000 ;
        RECT 1878.975 137.800 1879.490 137.940 ;
        RECT 1879.170 137.740 1879.490 137.800 ;
        RECT 1879.170 104.280 1879.490 104.340 ;
        RECT 1878.975 104.140 1879.490 104.280 ;
        RECT 1879.170 104.080 1879.490 104.140 ;
        RECT 1879.170 14.180 1879.490 14.240 ;
        RECT 1784.500 14.040 1879.490 14.180 ;
        RECT 1780.730 13.500 1781.050 13.560 ;
        RECT 1784.500 13.500 1784.640 14.040 ;
        RECT 1879.170 13.980 1879.490 14.040 ;
        RECT 1780.730 13.360 1784.640 13.500 ;
        RECT 1780.730 13.300 1781.050 13.360 ;
      LAYER via ;
        RECT 1879.200 1607.900 1879.460 1608.160 ;
        RECT 1879.660 1606.880 1879.920 1607.140 ;
        RECT 1879.200 1449.120 1879.460 1449.380 ;
        RECT 1879.660 1449.120 1879.920 1449.380 ;
        RECT 1879.200 1400.500 1879.460 1400.760 ;
        RECT 1879.200 1352.560 1879.460 1352.820 ;
        RECT 1879.200 1303.940 1879.460 1304.200 ;
        RECT 1879.200 1256.000 1879.460 1256.260 ;
        RECT 1879.200 1207.040 1879.460 1207.300 ;
        RECT 1879.200 1159.100 1879.460 1159.360 ;
        RECT 1879.200 1110.480 1879.460 1110.740 ;
        RECT 1879.200 1062.540 1879.460 1062.800 ;
        RECT 1879.200 1013.920 1879.460 1014.180 ;
        RECT 1879.200 965.980 1879.460 966.240 ;
        RECT 1879.200 882.000 1879.460 882.260 ;
        RECT 1879.660 882.000 1879.920 882.260 ;
        RECT 1879.660 820.800 1879.920 821.060 ;
        RECT 1879.200 772.860 1879.460 773.120 ;
        RECT 1879.200 651.820 1879.460 652.080 ;
        RECT 1880.580 651.820 1880.840 652.080 ;
        RECT 1879.200 627.680 1879.460 627.940 ;
        RECT 1878.740 579.740 1879.000 580.000 ;
        RECT 1878.740 545.060 1879.000 545.320 ;
        RECT 1879.200 544.720 1879.460 544.980 ;
        RECT 1879.200 434.560 1879.460 434.820 ;
        RECT 1879.200 386.280 1879.460 386.540 ;
        RECT 1879.200 352.280 1879.460 352.540 ;
        RECT 1879.200 351.600 1879.460 351.860 ;
        RECT 1879.200 255.720 1879.460 255.980 ;
        RECT 1879.200 255.040 1879.460 255.300 ;
        RECT 1878.740 234.300 1879.000 234.560 ;
        RECT 1879.200 234.300 1879.460 234.560 ;
        RECT 1878.740 144.880 1879.000 145.140 ;
        RECT 1879.200 144.880 1879.460 145.140 ;
        RECT 1879.200 137.740 1879.460 138.000 ;
        RECT 1879.200 104.080 1879.460 104.340 ;
        RECT 1780.760 13.300 1781.020 13.560 ;
        RECT 1879.200 13.980 1879.460 14.240 ;
      LAYER met2 ;
        RECT 1882.345 1700.410 1882.625 1704.000 ;
        RECT 1880.180 1700.270 1882.625 1700.410 ;
        RECT 1880.180 1684.770 1880.320 1700.270 ;
        RECT 1882.345 1700.000 1882.625 1700.270 ;
        RECT 1879.260 1684.630 1880.320 1684.770 ;
        RECT 1879.260 1608.190 1879.400 1684.630 ;
        RECT 1879.200 1607.870 1879.460 1608.190 ;
        RECT 1879.660 1606.850 1879.920 1607.170 ;
        RECT 1879.720 1449.410 1879.860 1606.850 ;
        RECT 1879.200 1449.090 1879.460 1449.410 ;
        RECT 1879.660 1449.090 1879.920 1449.410 ;
        RECT 1879.260 1400.790 1879.400 1449.090 ;
        RECT 1879.200 1400.470 1879.460 1400.790 ;
        RECT 1879.200 1352.530 1879.460 1352.850 ;
        RECT 1879.260 1304.230 1879.400 1352.530 ;
        RECT 1879.200 1303.910 1879.460 1304.230 ;
        RECT 1879.200 1255.970 1879.460 1256.290 ;
        RECT 1879.260 1207.330 1879.400 1255.970 ;
        RECT 1879.200 1207.010 1879.460 1207.330 ;
        RECT 1879.200 1159.070 1879.460 1159.390 ;
        RECT 1879.260 1110.770 1879.400 1159.070 ;
        RECT 1879.200 1110.450 1879.460 1110.770 ;
        RECT 1879.200 1062.510 1879.460 1062.830 ;
        RECT 1879.260 1014.210 1879.400 1062.510 ;
        RECT 1879.200 1013.890 1879.460 1014.210 ;
        RECT 1879.200 965.950 1879.460 966.270 ;
        RECT 1879.260 882.290 1879.400 965.950 ;
        RECT 1879.200 881.970 1879.460 882.290 ;
        RECT 1879.660 881.970 1879.920 882.290 ;
        RECT 1879.720 821.090 1879.860 881.970 ;
        RECT 1879.660 820.770 1879.920 821.090 ;
        RECT 1879.200 772.830 1879.460 773.150 ;
        RECT 1879.260 738.890 1879.400 772.830 ;
        RECT 1878.800 738.750 1879.400 738.890 ;
        RECT 1878.800 738.210 1878.940 738.750 ;
        RECT 1878.800 738.070 1879.400 738.210 ;
        RECT 1879.260 652.110 1879.400 738.070 ;
        RECT 1879.200 651.790 1879.460 652.110 ;
        RECT 1880.580 651.790 1880.840 652.110 ;
        RECT 1880.640 628.165 1880.780 651.790 ;
        RECT 1879.190 627.795 1879.470 628.165 ;
        RECT 1880.570 627.795 1880.850 628.165 ;
        RECT 1879.200 627.650 1879.460 627.795 ;
        RECT 1878.740 579.710 1879.000 580.030 ;
        RECT 1878.800 545.350 1878.940 579.710 ;
        RECT 1878.740 545.030 1879.000 545.350 ;
        RECT 1879.200 544.690 1879.460 545.010 ;
        RECT 1879.260 434.850 1879.400 544.690 ;
        RECT 1879.200 434.530 1879.460 434.850 ;
        RECT 1879.200 386.250 1879.460 386.570 ;
        RECT 1879.260 352.570 1879.400 386.250 ;
        RECT 1879.200 352.250 1879.460 352.570 ;
        RECT 1879.200 351.570 1879.460 351.890 ;
        RECT 1879.260 256.010 1879.400 351.570 ;
        RECT 1879.200 255.690 1879.460 256.010 ;
        RECT 1879.200 255.010 1879.460 255.330 ;
        RECT 1879.260 234.590 1879.400 255.010 ;
        RECT 1878.740 234.270 1879.000 234.590 ;
        RECT 1879.200 234.270 1879.460 234.590 ;
        RECT 1878.800 145.170 1878.940 234.270 ;
        RECT 1878.740 144.850 1879.000 145.170 ;
        RECT 1879.200 144.850 1879.460 145.170 ;
        RECT 1879.260 138.030 1879.400 144.850 ;
        RECT 1879.200 137.710 1879.460 138.030 ;
        RECT 1879.200 104.050 1879.460 104.370 ;
        RECT 1879.260 14.270 1879.400 104.050 ;
        RECT 1879.200 13.950 1879.460 14.270 ;
        RECT 1780.760 13.270 1781.020 13.590 ;
        RECT 1780.820 2.400 1780.960 13.270 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
      LAYER via2 ;
        RECT 1879.190 627.840 1879.470 628.120 ;
        RECT 1880.570 627.840 1880.850 628.120 ;
      LAYER met3 ;
        RECT 1879.165 628.130 1879.495 628.145 ;
        RECT 1880.545 628.130 1880.875 628.145 ;
        RECT 1879.165 627.830 1880.875 628.130 ;
        RECT 1879.165 627.815 1879.495 627.830 ;
        RECT 1880.545 627.815 1880.875 627.830 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1885.685 1352.605 1885.855 1400.715 ;
        RECT 1885.685 1256.045 1885.855 1304.155 ;
        RECT 1885.225 572.645 1885.395 620.755 ;
        RECT 1885.685 386.325 1885.855 434.775 ;
        RECT 1885.685 338.045 1885.855 352.495 ;
      LAYER mcon ;
        RECT 1885.685 1400.545 1885.855 1400.715 ;
        RECT 1885.685 1303.985 1885.855 1304.155 ;
        RECT 1885.225 620.585 1885.395 620.755 ;
        RECT 1885.685 434.605 1885.855 434.775 ;
        RECT 1885.685 352.325 1885.855 352.495 ;
      LAYER met1 ;
        RECT 1885.610 1607.900 1885.930 1608.160 ;
        RECT 1885.700 1607.080 1885.840 1607.900 ;
        RECT 1886.070 1607.080 1886.390 1607.140 ;
        RECT 1885.700 1606.940 1886.390 1607.080 ;
        RECT 1886.070 1606.880 1886.390 1606.940 ;
        RECT 1885.610 1449.320 1885.930 1449.380 ;
        RECT 1886.070 1449.320 1886.390 1449.380 ;
        RECT 1885.610 1449.180 1886.390 1449.320 ;
        RECT 1885.610 1449.120 1885.930 1449.180 ;
        RECT 1886.070 1449.120 1886.390 1449.180 ;
        RECT 1885.610 1400.700 1885.930 1400.760 ;
        RECT 1885.415 1400.560 1885.930 1400.700 ;
        RECT 1885.610 1400.500 1885.930 1400.560 ;
        RECT 1885.610 1352.760 1885.930 1352.820 ;
        RECT 1885.415 1352.620 1885.930 1352.760 ;
        RECT 1885.610 1352.560 1885.930 1352.620 ;
        RECT 1885.610 1304.140 1885.930 1304.200 ;
        RECT 1885.415 1304.000 1885.930 1304.140 ;
        RECT 1885.610 1303.940 1885.930 1304.000 ;
        RECT 1885.610 1256.200 1885.930 1256.260 ;
        RECT 1885.415 1256.060 1885.930 1256.200 ;
        RECT 1885.610 1256.000 1885.930 1256.060 ;
        RECT 1884.690 1159.300 1885.010 1159.360 ;
        RECT 1885.610 1159.300 1885.930 1159.360 ;
        RECT 1884.690 1159.160 1885.930 1159.300 ;
        RECT 1884.690 1159.100 1885.010 1159.160 ;
        RECT 1885.610 1159.100 1885.930 1159.160 ;
        RECT 1884.690 1062.740 1885.010 1062.800 ;
        RECT 1885.610 1062.740 1885.930 1062.800 ;
        RECT 1884.690 1062.600 1885.930 1062.740 ;
        RECT 1884.690 1062.540 1885.010 1062.600 ;
        RECT 1885.610 1062.540 1885.930 1062.600 ;
        RECT 1884.690 966.180 1885.010 966.240 ;
        RECT 1885.610 966.180 1885.930 966.240 ;
        RECT 1884.690 966.040 1885.930 966.180 ;
        RECT 1884.690 965.980 1885.010 966.040 ;
        RECT 1885.610 965.980 1885.930 966.040 ;
        RECT 1884.690 869.620 1885.010 869.680 ;
        RECT 1885.150 869.620 1885.470 869.680 ;
        RECT 1884.690 869.480 1885.470 869.620 ;
        RECT 1884.690 869.420 1885.010 869.480 ;
        RECT 1885.150 869.420 1885.470 869.480 ;
        RECT 1885.610 628.220 1885.930 628.280 ;
        RECT 1886.070 628.220 1886.390 628.280 ;
        RECT 1885.610 628.080 1886.390 628.220 ;
        RECT 1885.610 628.020 1885.930 628.080 ;
        RECT 1886.070 628.020 1886.390 628.080 ;
        RECT 1885.165 620.740 1885.455 620.785 ;
        RECT 1885.610 620.740 1885.930 620.800 ;
        RECT 1885.165 620.600 1885.930 620.740 ;
        RECT 1885.165 620.555 1885.455 620.600 ;
        RECT 1885.610 620.540 1885.930 620.600 ;
        RECT 1885.150 572.800 1885.470 572.860 ;
        RECT 1884.955 572.660 1885.470 572.800 ;
        RECT 1885.150 572.600 1885.470 572.660 ;
        RECT 1885.150 545.060 1885.470 545.320 ;
        RECT 1885.240 544.920 1885.380 545.060 ;
        RECT 1885.610 544.920 1885.930 544.980 ;
        RECT 1885.240 544.780 1885.930 544.920 ;
        RECT 1885.610 544.720 1885.930 544.780 ;
        RECT 1885.610 497.120 1885.930 497.380 ;
        RECT 1885.700 496.700 1885.840 497.120 ;
        RECT 1885.610 496.440 1885.930 496.700 ;
        RECT 1885.610 434.760 1885.930 434.820 ;
        RECT 1885.415 434.620 1885.930 434.760 ;
        RECT 1885.610 434.560 1885.930 434.620 ;
        RECT 1885.610 386.480 1885.930 386.540 ;
        RECT 1885.415 386.340 1885.930 386.480 ;
        RECT 1885.610 386.280 1885.930 386.340 ;
        RECT 1885.610 352.480 1885.930 352.540 ;
        RECT 1885.415 352.340 1885.930 352.480 ;
        RECT 1885.610 352.280 1885.930 352.340 ;
        RECT 1885.610 338.200 1885.930 338.260 ;
        RECT 1885.415 338.060 1885.930 338.200 ;
        RECT 1885.610 338.000 1885.930 338.060 ;
        RECT 1885.150 234.500 1885.470 234.560 ;
        RECT 1885.610 234.500 1885.930 234.560 ;
        RECT 1885.150 234.360 1885.930 234.500 ;
        RECT 1885.150 234.300 1885.470 234.360 ;
        RECT 1885.610 234.300 1885.930 234.360 ;
        RECT 1885.610 158.820 1885.930 159.080 ;
        RECT 1885.700 158.400 1885.840 158.820 ;
        RECT 1885.610 158.140 1885.930 158.400 ;
        RECT 1885.610 110.540 1885.930 110.800 ;
        RECT 1885.700 110.120 1885.840 110.540 ;
        RECT 1885.610 109.860 1885.930 110.120 ;
        RECT 1798.670 19.960 1798.990 20.020 ;
        RECT 1885.610 19.960 1885.930 20.020 ;
        RECT 1798.670 19.820 1885.930 19.960 ;
        RECT 1798.670 19.760 1798.990 19.820 ;
        RECT 1885.610 19.760 1885.930 19.820 ;
      LAYER via ;
        RECT 1885.640 1607.900 1885.900 1608.160 ;
        RECT 1886.100 1606.880 1886.360 1607.140 ;
        RECT 1885.640 1449.120 1885.900 1449.380 ;
        RECT 1886.100 1449.120 1886.360 1449.380 ;
        RECT 1885.640 1400.500 1885.900 1400.760 ;
        RECT 1885.640 1352.560 1885.900 1352.820 ;
        RECT 1885.640 1303.940 1885.900 1304.200 ;
        RECT 1885.640 1256.000 1885.900 1256.260 ;
        RECT 1884.720 1159.100 1884.980 1159.360 ;
        RECT 1885.640 1159.100 1885.900 1159.360 ;
        RECT 1884.720 1062.540 1884.980 1062.800 ;
        RECT 1885.640 1062.540 1885.900 1062.800 ;
        RECT 1884.720 965.980 1884.980 966.240 ;
        RECT 1885.640 965.980 1885.900 966.240 ;
        RECT 1884.720 869.420 1884.980 869.680 ;
        RECT 1885.180 869.420 1885.440 869.680 ;
        RECT 1885.640 628.020 1885.900 628.280 ;
        RECT 1886.100 628.020 1886.360 628.280 ;
        RECT 1885.640 620.540 1885.900 620.800 ;
        RECT 1885.180 572.600 1885.440 572.860 ;
        RECT 1885.180 545.060 1885.440 545.320 ;
        RECT 1885.640 544.720 1885.900 544.980 ;
        RECT 1885.640 497.120 1885.900 497.380 ;
        RECT 1885.640 496.440 1885.900 496.700 ;
        RECT 1885.640 434.560 1885.900 434.820 ;
        RECT 1885.640 386.280 1885.900 386.540 ;
        RECT 1885.640 352.280 1885.900 352.540 ;
        RECT 1885.640 338.000 1885.900 338.260 ;
        RECT 1885.180 234.300 1885.440 234.560 ;
        RECT 1885.640 234.300 1885.900 234.560 ;
        RECT 1885.640 158.820 1885.900 159.080 ;
        RECT 1885.640 158.140 1885.900 158.400 ;
        RECT 1885.640 110.540 1885.900 110.800 ;
        RECT 1885.640 109.860 1885.900 110.120 ;
        RECT 1798.700 19.760 1798.960 20.020 ;
        RECT 1885.640 19.760 1885.900 20.020 ;
      LAYER met2 ;
        RECT 1889.245 1700.410 1889.525 1704.000 ;
        RECT 1887.540 1700.270 1889.525 1700.410 ;
        RECT 1887.540 1677.970 1887.680 1700.270 ;
        RECT 1889.245 1700.000 1889.525 1700.270 ;
        RECT 1885.700 1677.830 1887.680 1677.970 ;
        RECT 1885.700 1608.190 1885.840 1677.830 ;
        RECT 1885.640 1607.870 1885.900 1608.190 ;
        RECT 1886.100 1606.850 1886.360 1607.170 ;
        RECT 1886.160 1449.410 1886.300 1606.850 ;
        RECT 1885.640 1449.090 1885.900 1449.410 ;
        RECT 1886.100 1449.090 1886.360 1449.410 ;
        RECT 1885.700 1400.790 1885.840 1449.090 ;
        RECT 1885.640 1400.470 1885.900 1400.790 ;
        RECT 1885.640 1352.530 1885.900 1352.850 ;
        RECT 1885.700 1304.230 1885.840 1352.530 ;
        RECT 1885.640 1303.910 1885.900 1304.230 ;
        RECT 1885.640 1255.970 1885.900 1256.290 ;
        RECT 1885.700 1207.525 1885.840 1255.970 ;
        RECT 1884.710 1207.155 1884.990 1207.525 ;
        RECT 1885.630 1207.155 1885.910 1207.525 ;
        RECT 1884.780 1159.390 1884.920 1207.155 ;
        RECT 1884.720 1159.070 1884.980 1159.390 ;
        RECT 1885.640 1159.070 1885.900 1159.390 ;
        RECT 1885.700 1110.965 1885.840 1159.070 ;
        RECT 1884.710 1110.595 1884.990 1110.965 ;
        RECT 1885.630 1110.595 1885.910 1110.965 ;
        RECT 1884.780 1062.830 1884.920 1110.595 ;
        RECT 1884.720 1062.510 1884.980 1062.830 ;
        RECT 1885.640 1062.510 1885.900 1062.830 ;
        RECT 1885.700 1014.405 1885.840 1062.510 ;
        RECT 1884.710 1014.035 1884.990 1014.405 ;
        RECT 1885.630 1014.035 1885.910 1014.405 ;
        RECT 1884.780 966.270 1884.920 1014.035 ;
        RECT 1884.720 965.950 1884.980 966.270 ;
        RECT 1885.640 965.950 1885.900 966.270 ;
        RECT 1885.700 917.845 1885.840 965.950 ;
        RECT 1884.710 917.475 1884.990 917.845 ;
        RECT 1885.630 917.475 1885.910 917.845 ;
        RECT 1884.780 869.710 1884.920 917.475 ;
        RECT 1884.720 869.390 1884.980 869.710 ;
        RECT 1885.180 869.390 1885.440 869.710 ;
        RECT 1885.240 834.770 1885.380 869.390 ;
        RECT 1885.240 834.630 1885.840 834.770 ;
        RECT 1885.700 738.890 1885.840 834.630 ;
        RECT 1885.240 738.750 1885.840 738.890 ;
        RECT 1885.240 738.210 1885.380 738.750 ;
        RECT 1885.240 738.070 1885.840 738.210 ;
        RECT 1885.700 643.010 1885.840 738.070 ;
        RECT 1885.700 642.870 1886.300 643.010 ;
        RECT 1886.160 628.310 1886.300 642.870 ;
        RECT 1885.640 627.990 1885.900 628.310 ;
        RECT 1886.100 627.990 1886.360 628.310 ;
        RECT 1885.700 620.830 1885.840 627.990 ;
        RECT 1885.640 620.510 1885.900 620.830 ;
        RECT 1885.180 572.570 1885.440 572.890 ;
        RECT 1885.240 545.350 1885.380 572.570 ;
        RECT 1885.180 545.030 1885.440 545.350 ;
        RECT 1885.640 544.690 1885.900 545.010 ;
        RECT 1885.700 497.410 1885.840 544.690 ;
        RECT 1885.640 497.090 1885.900 497.410 ;
        RECT 1885.640 496.410 1885.900 496.730 ;
        RECT 1885.700 434.850 1885.840 496.410 ;
        RECT 1885.640 434.530 1885.900 434.850 ;
        RECT 1885.640 386.250 1885.900 386.570 ;
        RECT 1885.700 352.570 1885.840 386.250 ;
        RECT 1885.640 352.250 1885.900 352.570 ;
        RECT 1885.640 337.970 1885.900 338.290 ;
        RECT 1885.700 256.090 1885.840 337.970 ;
        RECT 1885.700 255.950 1886.300 256.090 ;
        RECT 1886.160 235.010 1886.300 255.950 ;
        RECT 1885.700 234.870 1886.300 235.010 ;
        RECT 1885.700 234.590 1885.840 234.870 ;
        RECT 1885.180 234.270 1885.440 234.590 ;
        RECT 1885.640 234.270 1885.900 234.590 ;
        RECT 1885.240 199.650 1885.380 234.270 ;
        RECT 1885.240 199.510 1885.840 199.650 ;
        RECT 1885.700 159.110 1885.840 199.510 ;
        RECT 1885.640 158.790 1885.900 159.110 ;
        RECT 1885.640 158.110 1885.900 158.430 ;
        RECT 1885.700 110.830 1885.840 158.110 ;
        RECT 1885.640 110.510 1885.900 110.830 ;
        RECT 1885.640 109.830 1885.900 110.150 ;
        RECT 1885.700 20.050 1885.840 109.830 ;
        RECT 1798.700 19.730 1798.960 20.050 ;
        RECT 1885.640 19.730 1885.900 20.050 ;
        RECT 1798.760 2.400 1798.900 19.730 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
      LAYER via2 ;
        RECT 1884.710 1207.200 1884.990 1207.480 ;
        RECT 1885.630 1207.200 1885.910 1207.480 ;
        RECT 1884.710 1110.640 1884.990 1110.920 ;
        RECT 1885.630 1110.640 1885.910 1110.920 ;
        RECT 1884.710 1014.080 1884.990 1014.360 ;
        RECT 1885.630 1014.080 1885.910 1014.360 ;
        RECT 1884.710 917.520 1884.990 917.800 ;
        RECT 1885.630 917.520 1885.910 917.800 ;
      LAYER met3 ;
        RECT 1884.685 1207.490 1885.015 1207.505 ;
        RECT 1885.605 1207.490 1885.935 1207.505 ;
        RECT 1884.685 1207.190 1885.935 1207.490 ;
        RECT 1884.685 1207.175 1885.015 1207.190 ;
        RECT 1885.605 1207.175 1885.935 1207.190 ;
        RECT 1884.685 1110.930 1885.015 1110.945 ;
        RECT 1885.605 1110.930 1885.935 1110.945 ;
        RECT 1884.685 1110.630 1885.935 1110.930 ;
        RECT 1884.685 1110.615 1885.015 1110.630 ;
        RECT 1885.605 1110.615 1885.935 1110.630 ;
        RECT 1884.685 1014.370 1885.015 1014.385 ;
        RECT 1885.605 1014.370 1885.935 1014.385 ;
        RECT 1884.685 1014.070 1885.935 1014.370 ;
        RECT 1884.685 1014.055 1885.015 1014.070 ;
        RECT 1885.605 1014.055 1885.935 1014.070 ;
        RECT 1884.685 917.810 1885.015 917.825 ;
        RECT 1885.605 917.810 1885.935 917.825 ;
        RECT 1884.685 917.510 1885.935 917.810 ;
        RECT 1884.685 917.495 1885.015 917.510 ;
        RECT 1885.605 917.495 1885.935 917.510 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1821.210 1690.040 1821.530 1690.100 ;
        RECT 1896.650 1690.040 1896.970 1690.100 ;
        RECT 1821.210 1689.900 1896.970 1690.040 ;
        RECT 1821.210 1689.840 1821.530 1689.900 ;
        RECT 1896.650 1689.840 1896.970 1689.900 ;
        RECT 1816.610 20.640 1816.930 20.700 ;
        RECT 1821.210 20.640 1821.530 20.700 ;
        RECT 1816.610 20.500 1821.530 20.640 ;
        RECT 1816.610 20.440 1816.930 20.500 ;
        RECT 1821.210 20.440 1821.530 20.500 ;
      LAYER via ;
        RECT 1821.240 1689.840 1821.500 1690.100 ;
        RECT 1896.680 1689.840 1896.940 1690.100 ;
        RECT 1816.640 20.440 1816.900 20.700 ;
        RECT 1821.240 20.440 1821.500 20.700 ;
      LAYER met2 ;
        RECT 1896.605 1700.000 1896.885 1704.000 ;
        RECT 1896.740 1690.130 1896.880 1700.000 ;
        RECT 1821.240 1689.810 1821.500 1690.130 ;
        RECT 1896.680 1689.810 1896.940 1690.130 ;
        RECT 1821.300 20.730 1821.440 1689.810 ;
        RECT 1816.640 20.410 1816.900 20.730 ;
        RECT 1821.240 20.410 1821.500 20.730 ;
        RECT 1816.700 2.400 1816.840 20.410 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1834.625 1642.285 1834.795 1689.375 ;
        RECT 1835.085 1594.005 1835.255 1641.775 ;
        RECT 1835.085 1497.445 1835.255 1545.555 ;
        RECT 1835.085 1400.885 1835.255 1448.995 ;
        RECT 1835.085 1304.325 1835.255 1352.435 ;
        RECT 1835.085 1207.425 1835.255 1255.535 ;
        RECT 1835.085 1110.865 1835.255 1158.975 ;
        RECT 1835.085 1014.305 1835.255 1062.415 ;
        RECT 1835.085 917.745 1835.255 965.855 ;
        RECT 1835.085 773.245 1835.255 821.015 ;
        RECT 1835.085 676.685 1835.255 724.455 ;
        RECT 1835.085 628.065 1835.255 676.175 ;
        RECT 1835.085 483.565 1835.255 531.335 ;
        RECT 1835.085 379.525 1835.255 427.635 ;
        RECT 1835.085 241.825 1835.255 331.075 ;
        RECT 1834.165 186.405 1834.335 234.515 ;
        RECT 1834.165 48.365 1834.335 137.955 ;
      LAYER mcon ;
        RECT 1834.625 1689.205 1834.795 1689.375 ;
        RECT 1835.085 1641.605 1835.255 1641.775 ;
        RECT 1835.085 1545.385 1835.255 1545.555 ;
        RECT 1835.085 1448.825 1835.255 1448.995 ;
        RECT 1835.085 1352.265 1835.255 1352.435 ;
        RECT 1835.085 1255.365 1835.255 1255.535 ;
        RECT 1835.085 1158.805 1835.255 1158.975 ;
        RECT 1835.085 1062.245 1835.255 1062.415 ;
        RECT 1835.085 965.685 1835.255 965.855 ;
        RECT 1835.085 820.845 1835.255 821.015 ;
        RECT 1835.085 724.285 1835.255 724.455 ;
        RECT 1835.085 676.005 1835.255 676.175 ;
        RECT 1835.085 531.165 1835.255 531.335 ;
        RECT 1835.085 427.465 1835.255 427.635 ;
        RECT 1835.085 330.905 1835.255 331.075 ;
        RECT 1834.165 234.345 1834.335 234.515 ;
        RECT 1834.165 137.785 1834.335 137.955 ;
      LAYER met1 ;
        RECT 1834.565 1689.360 1834.855 1689.405 ;
        RECT 1904.010 1689.360 1904.330 1689.420 ;
        RECT 1834.565 1689.220 1904.330 1689.360 ;
        RECT 1834.565 1689.175 1834.855 1689.220 ;
        RECT 1904.010 1689.160 1904.330 1689.220 ;
        RECT 1834.565 1642.440 1834.855 1642.485 ;
        RECT 1835.010 1642.440 1835.330 1642.500 ;
        RECT 1834.565 1642.300 1835.330 1642.440 ;
        RECT 1834.565 1642.255 1834.855 1642.300 ;
        RECT 1835.010 1642.240 1835.330 1642.300 ;
        RECT 1835.010 1641.760 1835.330 1641.820 ;
        RECT 1834.815 1641.620 1835.330 1641.760 ;
        RECT 1835.010 1641.560 1835.330 1641.620 ;
        RECT 1835.010 1594.160 1835.330 1594.220 ;
        RECT 1834.815 1594.020 1835.330 1594.160 ;
        RECT 1835.010 1593.960 1835.330 1594.020 ;
        RECT 1835.010 1545.540 1835.330 1545.600 ;
        RECT 1834.815 1545.400 1835.330 1545.540 ;
        RECT 1835.010 1545.340 1835.330 1545.400 ;
        RECT 1835.010 1497.600 1835.330 1497.660 ;
        RECT 1834.815 1497.460 1835.330 1497.600 ;
        RECT 1835.010 1497.400 1835.330 1497.460 ;
        RECT 1835.010 1448.980 1835.330 1449.040 ;
        RECT 1834.815 1448.840 1835.330 1448.980 ;
        RECT 1835.010 1448.780 1835.330 1448.840 ;
        RECT 1835.010 1401.040 1835.330 1401.100 ;
        RECT 1834.815 1400.900 1835.330 1401.040 ;
        RECT 1835.010 1400.840 1835.330 1400.900 ;
        RECT 1835.010 1352.420 1835.330 1352.480 ;
        RECT 1834.815 1352.280 1835.330 1352.420 ;
        RECT 1835.010 1352.220 1835.330 1352.280 ;
        RECT 1835.010 1304.480 1835.330 1304.540 ;
        RECT 1834.815 1304.340 1835.330 1304.480 ;
        RECT 1835.010 1304.280 1835.330 1304.340 ;
        RECT 1835.010 1257.020 1835.330 1257.280 ;
        RECT 1835.100 1256.260 1835.240 1257.020 ;
        RECT 1835.010 1256.000 1835.330 1256.260 ;
        RECT 1835.010 1255.520 1835.330 1255.580 ;
        RECT 1834.815 1255.380 1835.330 1255.520 ;
        RECT 1835.010 1255.320 1835.330 1255.380 ;
        RECT 1835.010 1207.580 1835.330 1207.640 ;
        RECT 1834.815 1207.440 1835.330 1207.580 ;
        RECT 1835.010 1207.380 1835.330 1207.440 ;
        RECT 1835.010 1158.960 1835.330 1159.020 ;
        RECT 1834.815 1158.820 1835.330 1158.960 ;
        RECT 1835.010 1158.760 1835.330 1158.820 ;
        RECT 1835.010 1111.020 1835.330 1111.080 ;
        RECT 1834.815 1110.880 1835.330 1111.020 ;
        RECT 1835.010 1110.820 1835.330 1110.880 ;
        RECT 1835.010 1062.400 1835.330 1062.460 ;
        RECT 1834.815 1062.260 1835.330 1062.400 ;
        RECT 1835.010 1062.200 1835.330 1062.260 ;
        RECT 1835.010 1014.460 1835.330 1014.520 ;
        RECT 1834.815 1014.320 1835.330 1014.460 ;
        RECT 1835.010 1014.260 1835.330 1014.320 ;
        RECT 1835.010 965.840 1835.330 965.900 ;
        RECT 1834.815 965.700 1835.330 965.840 ;
        RECT 1835.010 965.640 1835.330 965.700 ;
        RECT 1835.010 917.900 1835.330 917.960 ;
        RECT 1834.815 917.760 1835.330 917.900 ;
        RECT 1835.010 917.700 1835.330 917.760 ;
        RECT 1834.090 870.300 1834.410 870.360 ;
        RECT 1835.010 870.300 1835.330 870.360 ;
        RECT 1834.090 870.160 1835.330 870.300 ;
        RECT 1834.090 870.100 1834.410 870.160 ;
        RECT 1835.010 870.100 1835.330 870.160 ;
        RECT 1835.010 821.000 1835.330 821.060 ;
        RECT 1834.815 820.860 1835.330 821.000 ;
        RECT 1835.010 820.800 1835.330 820.860 ;
        RECT 1835.010 773.400 1835.330 773.460 ;
        RECT 1834.815 773.260 1835.330 773.400 ;
        RECT 1835.010 773.200 1835.330 773.260 ;
        RECT 1833.630 772.720 1833.950 772.780 ;
        RECT 1835.010 772.720 1835.330 772.780 ;
        RECT 1833.630 772.580 1835.330 772.720 ;
        RECT 1833.630 772.520 1833.950 772.580 ;
        RECT 1835.010 772.520 1835.330 772.580 ;
        RECT 1835.010 724.440 1835.330 724.500 ;
        RECT 1834.815 724.300 1835.330 724.440 ;
        RECT 1835.010 724.240 1835.330 724.300 ;
        RECT 1835.010 676.840 1835.330 676.900 ;
        RECT 1834.815 676.700 1835.330 676.840 ;
        RECT 1835.010 676.640 1835.330 676.700 ;
        RECT 1835.010 676.160 1835.330 676.220 ;
        RECT 1834.815 676.020 1835.330 676.160 ;
        RECT 1835.010 675.960 1835.330 676.020 ;
        RECT 1835.010 628.220 1835.330 628.280 ;
        RECT 1834.815 628.080 1835.330 628.220 ;
        RECT 1835.010 628.020 1835.330 628.080 ;
        RECT 1833.630 579.600 1833.950 579.660 ;
        RECT 1835.010 579.600 1835.330 579.660 ;
        RECT 1833.630 579.460 1835.330 579.600 ;
        RECT 1833.630 579.400 1833.950 579.460 ;
        RECT 1835.010 579.400 1835.330 579.460 ;
        RECT 1835.010 531.320 1835.330 531.380 ;
        RECT 1834.815 531.180 1835.330 531.320 ;
        RECT 1835.010 531.120 1835.330 531.180 ;
        RECT 1835.010 483.720 1835.330 483.780 ;
        RECT 1834.815 483.580 1835.330 483.720 ;
        RECT 1835.010 483.520 1835.330 483.580 ;
        RECT 1835.010 427.620 1835.330 427.680 ;
        RECT 1834.815 427.480 1835.330 427.620 ;
        RECT 1835.010 427.420 1835.330 427.480 ;
        RECT 1835.010 379.680 1835.330 379.740 ;
        RECT 1834.815 379.540 1835.330 379.680 ;
        RECT 1835.010 379.480 1835.330 379.540 ;
        RECT 1835.010 331.060 1835.330 331.120 ;
        RECT 1834.815 330.920 1835.330 331.060 ;
        RECT 1835.010 330.860 1835.330 330.920 ;
        RECT 1835.010 241.980 1835.330 242.040 ;
        RECT 1834.815 241.840 1835.330 241.980 ;
        RECT 1835.010 241.780 1835.330 241.840 ;
        RECT 1834.105 234.500 1834.395 234.545 ;
        RECT 1835.010 234.500 1835.330 234.560 ;
        RECT 1834.105 234.360 1835.330 234.500 ;
        RECT 1834.105 234.315 1834.395 234.360 ;
        RECT 1835.010 234.300 1835.330 234.360 ;
        RECT 1834.090 186.560 1834.410 186.620 ;
        RECT 1833.895 186.420 1834.410 186.560 ;
        RECT 1834.090 186.360 1834.410 186.420 ;
        RECT 1834.090 146.100 1834.410 146.160 ;
        RECT 1834.090 145.960 1835.240 146.100 ;
        RECT 1834.090 145.900 1834.410 145.960 ;
        RECT 1835.100 145.820 1835.240 145.960 ;
        RECT 1835.010 145.560 1835.330 145.820 ;
        RECT 1834.105 137.940 1834.395 137.985 ;
        RECT 1835.010 137.940 1835.330 138.000 ;
        RECT 1834.105 137.800 1835.330 137.940 ;
        RECT 1834.105 137.755 1834.395 137.800 ;
        RECT 1835.010 137.740 1835.330 137.800 ;
        RECT 1834.090 48.520 1834.410 48.580 ;
        RECT 1833.895 48.380 1834.410 48.520 ;
        RECT 1834.090 48.320 1834.410 48.380 ;
      LAYER via ;
        RECT 1904.040 1689.160 1904.300 1689.420 ;
        RECT 1835.040 1642.240 1835.300 1642.500 ;
        RECT 1835.040 1641.560 1835.300 1641.820 ;
        RECT 1835.040 1593.960 1835.300 1594.220 ;
        RECT 1835.040 1545.340 1835.300 1545.600 ;
        RECT 1835.040 1497.400 1835.300 1497.660 ;
        RECT 1835.040 1448.780 1835.300 1449.040 ;
        RECT 1835.040 1400.840 1835.300 1401.100 ;
        RECT 1835.040 1352.220 1835.300 1352.480 ;
        RECT 1835.040 1304.280 1835.300 1304.540 ;
        RECT 1835.040 1257.020 1835.300 1257.280 ;
        RECT 1835.040 1256.000 1835.300 1256.260 ;
        RECT 1835.040 1255.320 1835.300 1255.580 ;
        RECT 1835.040 1207.380 1835.300 1207.640 ;
        RECT 1835.040 1158.760 1835.300 1159.020 ;
        RECT 1835.040 1110.820 1835.300 1111.080 ;
        RECT 1835.040 1062.200 1835.300 1062.460 ;
        RECT 1835.040 1014.260 1835.300 1014.520 ;
        RECT 1835.040 965.640 1835.300 965.900 ;
        RECT 1835.040 917.700 1835.300 917.960 ;
        RECT 1834.120 870.100 1834.380 870.360 ;
        RECT 1835.040 870.100 1835.300 870.360 ;
        RECT 1835.040 820.800 1835.300 821.060 ;
        RECT 1835.040 773.200 1835.300 773.460 ;
        RECT 1833.660 772.520 1833.920 772.780 ;
        RECT 1835.040 772.520 1835.300 772.780 ;
        RECT 1835.040 724.240 1835.300 724.500 ;
        RECT 1835.040 676.640 1835.300 676.900 ;
        RECT 1835.040 675.960 1835.300 676.220 ;
        RECT 1835.040 628.020 1835.300 628.280 ;
        RECT 1833.660 579.400 1833.920 579.660 ;
        RECT 1835.040 579.400 1835.300 579.660 ;
        RECT 1835.040 531.120 1835.300 531.380 ;
        RECT 1835.040 483.520 1835.300 483.780 ;
        RECT 1835.040 427.420 1835.300 427.680 ;
        RECT 1835.040 379.480 1835.300 379.740 ;
        RECT 1835.040 330.860 1835.300 331.120 ;
        RECT 1835.040 241.780 1835.300 242.040 ;
        RECT 1835.040 234.300 1835.300 234.560 ;
        RECT 1834.120 186.360 1834.380 186.620 ;
        RECT 1834.120 145.900 1834.380 146.160 ;
        RECT 1835.040 145.560 1835.300 145.820 ;
        RECT 1835.040 137.740 1835.300 138.000 ;
        RECT 1834.120 48.320 1834.380 48.580 ;
      LAYER met2 ;
        RECT 1903.965 1700.000 1904.245 1704.000 ;
        RECT 1904.100 1689.450 1904.240 1700.000 ;
        RECT 1904.040 1689.130 1904.300 1689.450 ;
        RECT 1835.040 1642.210 1835.300 1642.530 ;
        RECT 1835.100 1641.850 1835.240 1642.210 ;
        RECT 1835.040 1641.530 1835.300 1641.850 ;
        RECT 1835.040 1593.930 1835.300 1594.250 ;
        RECT 1835.100 1545.630 1835.240 1593.930 ;
        RECT 1835.040 1545.310 1835.300 1545.630 ;
        RECT 1835.040 1497.370 1835.300 1497.690 ;
        RECT 1835.100 1449.070 1835.240 1497.370 ;
        RECT 1835.040 1448.750 1835.300 1449.070 ;
        RECT 1835.040 1400.810 1835.300 1401.130 ;
        RECT 1835.100 1352.510 1835.240 1400.810 ;
        RECT 1835.040 1352.190 1835.300 1352.510 ;
        RECT 1835.040 1304.250 1835.300 1304.570 ;
        RECT 1835.100 1257.310 1835.240 1304.250 ;
        RECT 1835.040 1256.990 1835.300 1257.310 ;
        RECT 1835.040 1255.970 1835.300 1256.290 ;
        RECT 1835.100 1255.610 1835.240 1255.970 ;
        RECT 1835.040 1255.290 1835.300 1255.610 ;
        RECT 1835.040 1207.350 1835.300 1207.670 ;
        RECT 1835.100 1159.050 1835.240 1207.350 ;
        RECT 1835.040 1158.730 1835.300 1159.050 ;
        RECT 1835.040 1110.790 1835.300 1111.110 ;
        RECT 1835.100 1062.490 1835.240 1110.790 ;
        RECT 1835.040 1062.170 1835.300 1062.490 ;
        RECT 1835.040 1014.230 1835.300 1014.550 ;
        RECT 1835.100 965.930 1835.240 1014.230 ;
        RECT 1835.040 965.610 1835.300 965.930 ;
        RECT 1835.040 917.845 1835.300 917.990 ;
        RECT 1834.110 917.475 1834.390 917.845 ;
        RECT 1835.030 917.475 1835.310 917.845 ;
        RECT 1834.180 870.390 1834.320 917.475 ;
        RECT 1834.120 870.070 1834.380 870.390 ;
        RECT 1835.040 870.070 1835.300 870.390 ;
        RECT 1835.100 869.565 1835.240 870.070 ;
        RECT 1835.030 869.195 1835.310 869.565 ;
        RECT 1835.030 820.915 1835.310 821.285 ;
        RECT 1835.040 820.770 1835.300 820.915 ;
        RECT 1835.040 773.170 1835.300 773.490 ;
        RECT 1835.100 772.810 1835.240 773.170 ;
        RECT 1833.660 772.490 1833.920 772.810 ;
        RECT 1835.040 772.490 1835.300 772.810 ;
        RECT 1833.720 724.725 1833.860 772.490 ;
        RECT 1833.650 724.355 1833.930 724.725 ;
        RECT 1835.030 724.355 1835.310 724.725 ;
        RECT 1835.040 724.210 1835.300 724.355 ;
        RECT 1835.040 676.610 1835.300 676.930 ;
        RECT 1835.100 676.250 1835.240 676.610 ;
        RECT 1835.040 675.930 1835.300 676.250 ;
        RECT 1835.040 627.990 1835.300 628.310 ;
        RECT 1835.100 579.690 1835.240 627.990 ;
        RECT 1833.660 579.370 1833.920 579.690 ;
        RECT 1835.040 579.370 1835.300 579.690 ;
        RECT 1833.720 531.605 1833.860 579.370 ;
        RECT 1833.650 531.235 1833.930 531.605 ;
        RECT 1835.030 531.235 1835.310 531.605 ;
        RECT 1835.040 531.090 1835.300 531.235 ;
        RECT 1835.040 483.490 1835.300 483.810 ;
        RECT 1835.100 436.405 1835.240 483.490 ;
        RECT 1835.030 436.035 1835.310 436.405 ;
        RECT 1835.030 435.355 1835.310 435.725 ;
        RECT 1835.100 427.710 1835.240 435.355 ;
        RECT 1835.040 427.390 1835.300 427.710 ;
        RECT 1835.040 379.450 1835.300 379.770 ;
        RECT 1835.100 331.150 1835.240 379.450 ;
        RECT 1835.040 330.830 1835.300 331.150 ;
        RECT 1835.040 241.750 1835.300 242.070 ;
        RECT 1835.100 234.590 1835.240 241.750 ;
        RECT 1835.040 234.270 1835.300 234.590 ;
        RECT 1834.120 186.330 1834.380 186.650 ;
        RECT 1834.180 146.190 1834.320 186.330 ;
        RECT 1834.120 145.870 1834.380 146.190 ;
        RECT 1835.040 145.530 1835.300 145.850 ;
        RECT 1835.100 138.030 1835.240 145.530 ;
        RECT 1835.040 137.710 1835.300 138.030 ;
        RECT 1834.120 48.290 1834.380 48.610 ;
        RECT 1834.180 48.010 1834.320 48.290 ;
        RECT 1833.720 47.870 1834.320 48.010 ;
        RECT 1833.720 22.170 1833.860 47.870 ;
        RECT 1833.720 22.030 1834.780 22.170 ;
        RECT 1834.640 2.400 1834.780 22.030 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
      LAYER via2 ;
        RECT 1834.110 917.520 1834.390 917.800 ;
        RECT 1835.030 917.520 1835.310 917.800 ;
        RECT 1835.030 869.240 1835.310 869.520 ;
        RECT 1835.030 820.960 1835.310 821.240 ;
        RECT 1833.650 724.400 1833.930 724.680 ;
        RECT 1835.030 724.400 1835.310 724.680 ;
        RECT 1833.650 531.280 1833.930 531.560 ;
        RECT 1835.030 531.280 1835.310 531.560 ;
        RECT 1835.030 436.080 1835.310 436.360 ;
        RECT 1835.030 435.400 1835.310 435.680 ;
      LAYER met3 ;
        RECT 1834.085 917.810 1834.415 917.825 ;
        RECT 1835.005 917.810 1835.335 917.825 ;
        RECT 1834.085 917.510 1835.335 917.810 ;
        RECT 1834.085 917.495 1834.415 917.510 ;
        RECT 1835.005 917.495 1835.335 917.510 ;
        RECT 1835.005 869.540 1835.335 869.545 ;
        RECT 1834.750 869.530 1835.335 869.540 ;
        RECT 1834.550 869.230 1835.335 869.530 ;
        RECT 1834.750 869.220 1835.335 869.230 ;
        RECT 1835.005 869.215 1835.335 869.220 ;
        RECT 1835.005 821.260 1835.335 821.265 ;
        RECT 1834.750 821.250 1835.335 821.260 ;
        RECT 1834.550 820.950 1835.335 821.250 ;
        RECT 1834.750 820.940 1835.335 820.950 ;
        RECT 1835.005 820.935 1835.335 820.940 ;
        RECT 1833.625 724.690 1833.955 724.705 ;
        RECT 1835.005 724.690 1835.335 724.705 ;
        RECT 1833.625 724.390 1835.335 724.690 ;
        RECT 1833.625 724.375 1833.955 724.390 ;
        RECT 1835.005 724.375 1835.335 724.390 ;
        RECT 1833.625 531.570 1833.955 531.585 ;
        RECT 1835.005 531.570 1835.335 531.585 ;
        RECT 1833.625 531.270 1835.335 531.570 ;
        RECT 1833.625 531.255 1833.955 531.270 ;
        RECT 1835.005 531.255 1835.335 531.270 ;
        RECT 1835.005 436.370 1835.335 436.385 ;
        RECT 1834.790 436.055 1835.335 436.370 ;
        RECT 1834.790 435.705 1835.090 436.055 ;
        RECT 1834.790 435.390 1835.335 435.705 ;
        RECT 1835.005 435.375 1835.335 435.390 ;
      LAYER via3 ;
        RECT 1834.780 869.220 1835.100 869.540 ;
        RECT 1834.780 820.940 1835.100 821.260 ;
      LAYER met4 ;
        RECT 1834.775 869.215 1835.105 869.545 ;
        RECT 1834.790 821.265 1835.090 869.215 ;
        RECT 1834.775 820.935 1835.105 821.265 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1855.710 1689.700 1856.030 1689.760 ;
        RECT 1911.370 1689.700 1911.690 1689.760 ;
        RECT 1855.710 1689.560 1911.690 1689.700 ;
        RECT 1855.710 1689.500 1856.030 1689.560 ;
        RECT 1911.370 1689.500 1911.690 1689.560 ;
        RECT 1852.030 20.640 1852.350 20.700 ;
        RECT 1855.710 20.640 1856.030 20.700 ;
        RECT 1852.030 20.500 1856.030 20.640 ;
        RECT 1852.030 20.440 1852.350 20.500 ;
        RECT 1855.710 20.440 1856.030 20.500 ;
      LAYER via ;
        RECT 1855.740 1689.500 1856.000 1689.760 ;
        RECT 1911.400 1689.500 1911.660 1689.760 ;
        RECT 1852.060 20.440 1852.320 20.700 ;
        RECT 1855.740 20.440 1856.000 20.700 ;
      LAYER met2 ;
        RECT 1911.325 1700.000 1911.605 1704.000 ;
        RECT 1911.460 1689.790 1911.600 1700.000 ;
        RECT 1855.740 1689.470 1856.000 1689.790 ;
        RECT 1911.400 1689.470 1911.660 1689.790 ;
        RECT 1855.800 20.730 1855.940 1689.470 ;
        RECT 1852.060 20.410 1852.320 20.730 ;
        RECT 1855.740 20.410 1856.000 20.730 ;
        RECT 1852.120 2.400 1852.260 20.410 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1876.410 1687.320 1876.730 1687.380 ;
        RECT 1918.730 1687.320 1919.050 1687.380 ;
        RECT 1876.410 1687.180 1919.050 1687.320 ;
        RECT 1876.410 1687.120 1876.730 1687.180 ;
        RECT 1918.730 1687.120 1919.050 1687.180 ;
        RECT 1869.970 18.940 1870.290 19.000 ;
        RECT 1876.410 18.940 1876.730 19.000 ;
        RECT 1869.970 18.800 1876.730 18.940 ;
        RECT 1869.970 18.740 1870.290 18.800 ;
        RECT 1876.410 18.740 1876.730 18.800 ;
      LAYER via ;
        RECT 1876.440 1687.120 1876.700 1687.380 ;
        RECT 1918.760 1687.120 1919.020 1687.380 ;
        RECT 1870.000 18.740 1870.260 19.000 ;
        RECT 1876.440 18.740 1876.700 19.000 ;
      LAYER met2 ;
        RECT 1918.685 1700.000 1918.965 1704.000 ;
        RECT 1918.820 1687.410 1918.960 1700.000 ;
        RECT 1876.440 1687.090 1876.700 1687.410 ;
        RECT 1918.760 1687.090 1919.020 1687.410 ;
        RECT 1876.500 19.030 1876.640 1687.090 ;
        RECT 1870.000 18.710 1870.260 19.030 ;
        RECT 1876.440 18.710 1876.700 19.030 ;
        RECT 1870.060 2.400 1870.200 18.710 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 746.190 36.280 746.510 36.340 ;
        RECT 1455.970 36.280 1456.290 36.340 ;
        RECT 746.190 36.140 1456.290 36.280 ;
        RECT 746.190 36.080 746.510 36.140 ;
        RECT 1455.970 36.080 1456.290 36.140 ;
      LAYER via ;
        RECT 746.220 36.080 746.480 36.340 ;
        RECT 1456.000 36.080 1456.260 36.340 ;
      LAYER met2 ;
        RECT 1455.925 1700.000 1456.205 1704.000 ;
        RECT 1456.060 36.370 1456.200 1700.000 ;
        RECT 746.220 36.050 746.480 36.370 ;
        RECT 1456.000 36.050 1456.260 36.370 ;
        RECT 746.280 2.400 746.420 36.050 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1890.210 1684.940 1890.530 1685.000 ;
        RECT 1926.090 1684.940 1926.410 1685.000 ;
        RECT 1890.210 1684.800 1926.410 1684.940 ;
        RECT 1890.210 1684.740 1890.530 1684.800 ;
        RECT 1926.090 1684.740 1926.410 1684.800 ;
        RECT 1887.910 20.640 1888.230 20.700 ;
        RECT 1890.210 20.640 1890.530 20.700 ;
        RECT 1887.910 20.500 1890.530 20.640 ;
        RECT 1887.910 20.440 1888.230 20.500 ;
        RECT 1890.210 20.440 1890.530 20.500 ;
      LAYER via ;
        RECT 1890.240 1684.740 1890.500 1685.000 ;
        RECT 1926.120 1684.740 1926.380 1685.000 ;
        RECT 1887.940 20.440 1888.200 20.700 ;
        RECT 1890.240 20.440 1890.500 20.700 ;
      LAYER met2 ;
        RECT 1926.045 1700.000 1926.325 1704.000 ;
        RECT 1926.180 1685.030 1926.320 1700.000 ;
        RECT 1890.240 1684.710 1890.500 1685.030 ;
        RECT 1926.120 1684.710 1926.380 1685.030 ;
        RECT 1890.300 20.730 1890.440 1684.710 ;
        RECT 1887.940 20.410 1888.200 20.730 ;
        RECT 1890.240 20.410 1890.500 20.730 ;
        RECT 1888.000 2.400 1888.140 20.410 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1910.910 1686.980 1911.230 1687.040 ;
        RECT 1933.450 1686.980 1933.770 1687.040 ;
        RECT 1910.910 1686.840 1933.770 1686.980 ;
        RECT 1910.910 1686.780 1911.230 1686.840 ;
        RECT 1933.450 1686.780 1933.770 1686.840 ;
        RECT 1905.850 17.580 1906.170 17.640 ;
        RECT 1910.910 17.580 1911.230 17.640 ;
        RECT 1905.850 17.440 1911.230 17.580 ;
        RECT 1905.850 17.380 1906.170 17.440 ;
        RECT 1910.910 17.380 1911.230 17.440 ;
      LAYER via ;
        RECT 1910.940 1686.780 1911.200 1687.040 ;
        RECT 1933.480 1686.780 1933.740 1687.040 ;
        RECT 1905.880 17.380 1906.140 17.640 ;
        RECT 1910.940 17.380 1911.200 17.640 ;
      LAYER met2 ;
        RECT 1933.405 1700.000 1933.685 1704.000 ;
        RECT 1933.540 1687.070 1933.680 1700.000 ;
        RECT 1910.940 1686.750 1911.200 1687.070 ;
        RECT 1933.480 1686.750 1933.740 1687.070 ;
        RECT 1911.000 17.670 1911.140 1686.750 ;
        RECT 1905.880 17.350 1906.140 17.670 ;
        RECT 1910.940 17.350 1911.200 17.670 ;
        RECT 1905.940 2.400 1906.080 17.350 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1924.710 1688.680 1925.030 1688.740 ;
        RECT 1940.810 1688.680 1941.130 1688.740 ;
        RECT 1924.710 1688.540 1941.130 1688.680 ;
        RECT 1924.710 1688.480 1925.030 1688.540 ;
        RECT 1940.810 1688.480 1941.130 1688.540 ;
        RECT 1923.330 2.960 1923.650 3.020 ;
        RECT 1924.710 2.960 1925.030 3.020 ;
        RECT 1923.330 2.820 1925.030 2.960 ;
        RECT 1923.330 2.760 1923.650 2.820 ;
        RECT 1924.710 2.760 1925.030 2.820 ;
      LAYER via ;
        RECT 1924.740 1688.480 1925.000 1688.740 ;
        RECT 1940.840 1688.480 1941.100 1688.740 ;
        RECT 1923.360 2.760 1923.620 3.020 ;
        RECT 1924.740 2.760 1925.000 3.020 ;
      LAYER met2 ;
        RECT 1940.765 1700.000 1941.045 1704.000 ;
        RECT 1940.900 1688.770 1941.040 1700.000 ;
        RECT 1924.740 1688.450 1925.000 1688.770 ;
        RECT 1940.840 1688.450 1941.100 1688.770 ;
        RECT 1924.800 3.050 1924.940 1688.450 ;
        RECT 1923.360 2.730 1923.620 3.050 ;
        RECT 1924.740 2.730 1925.000 3.050 ;
        RECT 1923.420 2.400 1923.560 2.730 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1941.270 17.580 1941.590 17.640 ;
        RECT 1945.410 17.580 1945.730 17.640 ;
        RECT 1941.270 17.440 1945.730 17.580 ;
        RECT 1941.270 17.380 1941.590 17.440 ;
        RECT 1945.410 17.380 1945.730 17.440 ;
      LAYER via ;
        RECT 1941.300 17.380 1941.560 17.640 ;
        RECT 1945.440 17.380 1945.700 17.640 ;
      LAYER met2 ;
        RECT 1948.125 1700.410 1948.405 1704.000 ;
        RECT 1946.420 1700.270 1948.405 1700.410 ;
        RECT 1946.420 1688.850 1946.560 1700.270 ;
        RECT 1948.125 1700.000 1948.405 1700.270 ;
        RECT 1945.500 1688.710 1946.560 1688.850 ;
        RECT 1945.500 17.670 1945.640 1688.710 ;
        RECT 1941.300 17.350 1941.560 17.670 ;
        RECT 1945.440 17.350 1945.700 17.670 ;
        RECT 1941.360 2.400 1941.500 17.350 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1954.150 20.640 1954.470 20.700 ;
        RECT 1959.210 20.640 1959.530 20.700 ;
        RECT 1954.150 20.500 1959.530 20.640 ;
        RECT 1954.150 20.440 1954.470 20.500 ;
        RECT 1959.210 20.440 1959.530 20.500 ;
      LAYER via ;
        RECT 1954.180 20.440 1954.440 20.700 ;
        RECT 1959.240 20.440 1959.500 20.700 ;
      LAYER met2 ;
        RECT 1955.485 1700.410 1955.765 1704.000 ;
        RECT 1954.240 1700.270 1955.765 1700.410 ;
        RECT 1954.240 20.730 1954.380 1700.270 ;
        RECT 1955.485 1700.000 1955.765 1700.270 ;
        RECT 1954.180 20.410 1954.440 20.730 ;
        RECT 1959.240 20.410 1959.500 20.730 ;
        RECT 1959.300 2.400 1959.440 20.410 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1962.890 1683.920 1963.210 1683.980 ;
        RECT 1966.110 1683.920 1966.430 1683.980 ;
        RECT 1962.890 1683.780 1966.430 1683.920 ;
        RECT 1962.890 1683.720 1963.210 1683.780 ;
        RECT 1966.110 1683.720 1966.430 1683.780 ;
        RECT 1966.110 20.640 1966.430 20.700 ;
        RECT 1977.150 20.640 1977.470 20.700 ;
        RECT 1966.110 20.500 1977.470 20.640 ;
        RECT 1966.110 20.440 1966.430 20.500 ;
        RECT 1977.150 20.440 1977.470 20.500 ;
      LAYER via ;
        RECT 1962.920 1683.720 1963.180 1683.980 ;
        RECT 1966.140 1683.720 1966.400 1683.980 ;
        RECT 1966.140 20.440 1966.400 20.700 ;
        RECT 1977.180 20.440 1977.440 20.700 ;
      LAYER met2 ;
        RECT 1962.845 1700.000 1963.125 1704.000 ;
        RECT 1962.980 1684.010 1963.120 1700.000 ;
        RECT 1962.920 1683.690 1963.180 1684.010 ;
        RECT 1966.140 1683.690 1966.400 1684.010 ;
        RECT 1966.200 20.730 1966.340 1683.690 ;
        RECT 1966.140 20.410 1966.400 20.730 ;
        RECT 1977.180 20.410 1977.440 20.730 ;
        RECT 1977.240 2.400 1977.380 20.410 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1970.250 1683.920 1970.570 1683.980 ;
        RECT 1973.010 1683.920 1973.330 1683.980 ;
        RECT 1970.250 1683.780 1973.330 1683.920 ;
        RECT 1970.250 1683.720 1970.570 1683.780 ;
        RECT 1973.010 1683.720 1973.330 1683.780 ;
        RECT 1973.010 17.580 1973.330 17.640 ;
        RECT 1995.090 17.580 1995.410 17.640 ;
        RECT 1973.010 17.440 1995.410 17.580 ;
        RECT 1973.010 17.380 1973.330 17.440 ;
        RECT 1995.090 17.380 1995.410 17.440 ;
      LAYER via ;
        RECT 1970.280 1683.720 1970.540 1683.980 ;
        RECT 1973.040 1683.720 1973.300 1683.980 ;
        RECT 1973.040 17.380 1973.300 17.640 ;
        RECT 1995.120 17.380 1995.380 17.640 ;
      LAYER met2 ;
        RECT 1970.205 1700.000 1970.485 1704.000 ;
        RECT 1970.340 1684.010 1970.480 1700.000 ;
        RECT 1970.280 1683.690 1970.540 1684.010 ;
        RECT 1973.040 1683.690 1973.300 1684.010 ;
        RECT 1973.100 17.670 1973.240 1683.690 ;
        RECT 1973.040 17.350 1973.300 17.670 ;
        RECT 1995.120 17.350 1995.380 17.670 ;
        RECT 1995.180 2.400 1995.320 17.350 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1979.910 14.860 1980.230 14.920 ;
        RECT 2012.570 14.860 2012.890 14.920 ;
        RECT 1979.910 14.720 2012.890 14.860 ;
        RECT 1979.910 14.660 1980.230 14.720 ;
        RECT 2012.570 14.660 2012.890 14.720 ;
      LAYER via ;
        RECT 1979.940 14.660 1980.200 14.920 ;
        RECT 2012.600 14.660 2012.860 14.920 ;
      LAYER met2 ;
        RECT 1977.565 1700.410 1977.845 1704.000 ;
        RECT 1977.565 1700.270 1980.140 1700.410 ;
        RECT 1977.565 1700.000 1977.845 1700.270 ;
        RECT 1980.000 14.950 1980.140 1700.270 ;
        RECT 1979.940 14.630 1980.200 14.950 ;
        RECT 2012.600 14.630 2012.860 14.950 ;
        RECT 2012.660 2.400 2012.800 14.630 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1984.970 1686.640 1985.290 1686.700 ;
        RECT 2029.590 1686.640 2029.910 1686.700 ;
        RECT 1984.970 1686.500 2029.910 1686.640 ;
        RECT 1984.970 1686.440 1985.290 1686.500 ;
        RECT 2029.590 1686.440 2029.910 1686.500 ;
        RECT 2029.590 2.960 2029.910 3.020 ;
        RECT 2030.510 2.960 2030.830 3.020 ;
        RECT 2029.590 2.820 2030.830 2.960 ;
        RECT 2029.590 2.760 2029.910 2.820 ;
        RECT 2030.510 2.760 2030.830 2.820 ;
      LAYER via ;
        RECT 1985.000 1686.440 1985.260 1686.700 ;
        RECT 2029.620 1686.440 2029.880 1686.700 ;
        RECT 2029.620 2.760 2029.880 3.020 ;
        RECT 2030.540 2.760 2030.800 3.020 ;
      LAYER met2 ;
        RECT 1984.925 1700.000 1985.205 1704.000 ;
        RECT 1985.060 1686.730 1985.200 1700.000 ;
        RECT 1985.000 1686.410 1985.260 1686.730 ;
        RECT 2029.620 1686.410 2029.880 1686.730 ;
        RECT 2029.680 3.050 2029.820 1686.410 ;
        RECT 2029.620 2.730 2029.880 3.050 ;
        RECT 2030.540 2.730 2030.800 3.050 ;
        RECT 2030.600 2.400 2030.740 2.730 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1992.330 1687.320 1992.650 1687.380 ;
        RECT 1992.330 1687.180 2011.880 1687.320 ;
        RECT 1992.330 1687.120 1992.650 1687.180 ;
        RECT 2011.740 1686.980 2011.880 1687.180 ;
        RECT 2043.390 1686.980 2043.710 1687.040 ;
        RECT 2011.740 1686.840 2043.710 1686.980 ;
        RECT 2043.390 1686.780 2043.710 1686.840 ;
      LAYER via ;
        RECT 1992.360 1687.120 1992.620 1687.380 ;
        RECT 2043.420 1686.780 2043.680 1687.040 ;
      LAYER met2 ;
        RECT 1992.285 1700.000 1992.565 1704.000 ;
        RECT 1992.420 1687.410 1992.560 1700.000 ;
        RECT 1992.360 1687.090 1992.620 1687.410 ;
        RECT 2043.420 1686.750 2043.680 1687.070 ;
        RECT 2043.480 12.650 2043.620 1686.750 ;
        RECT 2043.480 12.510 2048.680 12.650 ;
        RECT 2048.540 2.400 2048.680 12.510 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 763.670 35.940 763.990 36.000 ;
        RECT 1462.870 35.940 1463.190 36.000 ;
        RECT 763.670 35.800 1463.190 35.940 ;
        RECT 763.670 35.740 763.990 35.800 ;
        RECT 1462.870 35.740 1463.190 35.800 ;
      LAYER via ;
        RECT 763.700 35.740 763.960 36.000 ;
        RECT 1462.900 35.740 1463.160 36.000 ;
      LAYER met2 ;
        RECT 1463.285 1700.410 1463.565 1704.000 ;
        RECT 1462.960 1700.270 1463.565 1700.410 ;
        RECT 1462.960 36.030 1463.100 1700.270 ;
        RECT 1463.285 1700.000 1463.565 1700.270 ;
        RECT 763.700 35.710 763.960 36.030 ;
        RECT 1462.900 35.710 1463.160 36.030 ;
        RECT 763.760 2.400 763.900 35.710 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1999.690 1689.360 2000.010 1689.420 ;
        RECT 2064.090 1689.360 2064.410 1689.420 ;
        RECT 1999.690 1689.220 2064.410 1689.360 ;
        RECT 1999.690 1689.160 2000.010 1689.220 ;
        RECT 2064.090 1689.160 2064.410 1689.220 ;
      LAYER via ;
        RECT 1999.720 1689.160 1999.980 1689.420 ;
        RECT 2064.120 1689.160 2064.380 1689.420 ;
      LAYER met2 ;
        RECT 1999.645 1700.000 1999.925 1704.000 ;
        RECT 1999.780 1689.450 1999.920 1700.000 ;
        RECT 1999.720 1689.130 1999.980 1689.450 ;
        RECT 2064.120 1689.130 2064.380 1689.450 ;
        RECT 2064.180 16.730 2064.320 1689.130 ;
        RECT 2064.180 16.590 2066.620 16.730 ;
        RECT 2066.480 2.400 2066.620 16.590 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2007.050 1685.280 2007.370 1685.340 ;
        RECT 2024.990 1685.280 2025.310 1685.340 ;
        RECT 2007.050 1685.140 2025.310 1685.280 ;
        RECT 2007.050 1685.080 2007.370 1685.140 ;
        RECT 2024.990 1685.080 2025.310 1685.140 ;
        RECT 2024.990 19.620 2025.310 19.680 ;
        RECT 2084.330 19.620 2084.650 19.680 ;
        RECT 2024.990 19.480 2084.650 19.620 ;
        RECT 2024.990 19.420 2025.310 19.480 ;
        RECT 2084.330 19.420 2084.650 19.480 ;
      LAYER via ;
        RECT 2007.080 1685.080 2007.340 1685.340 ;
        RECT 2025.020 1685.080 2025.280 1685.340 ;
        RECT 2025.020 19.420 2025.280 19.680 ;
        RECT 2084.360 19.420 2084.620 19.680 ;
      LAYER met2 ;
        RECT 2007.005 1700.000 2007.285 1704.000 ;
        RECT 2007.140 1685.370 2007.280 1700.000 ;
        RECT 2007.080 1685.050 2007.340 1685.370 ;
        RECT 2025.020 1685.050 2025.280 1685.370 ;
        RECT 2025.080 19.710 2025.220 1685.050 ;
        RECT 2025.020 19.390 2025.280 19.710 ;
        RECT 2084.360 19.390 2084.620 19.710 ;
        RECT 2084.420 2.400 2084.560 19.390 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2014.410 17.920 2014.730 17.980 ;
        RECT 2101.810 17.920 2102.130 17.980 ;
        RECT 2014.410 17.780 2102.130 17.920 ;
        RECT 2014.410 17.720 2014.730 17.780 ;
        RECT 2101.810 17.720 2102.130 17.780 ;
      LAYER via ;
        RECT 2014.440 17.720 2014.700 17.980 ;
        RECT 2101.840 17.720 2102.100 17.980 ;
      LAYER met2 ;
        RECT 2014.365 1700.000 2014.645 1704.000 ;
        RECT 2014.500 18.010 2014.640 1700.000 ;
        RECT 2014.440 17.690 2014.700 18.010 ;
        RECT 2101.840 17.690 2102.100 18.010 ;
        RECT 2101.900 2.400 2102.040 17.690 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2062.340 1688.540 2068.000 1688.680 ;
        RECT 2021.770 1688.340 2022.090 1688.400 ;
        RECT 2062.340 1688.340 2062.480 1688.540 ;
        RECT 2021.770 1688.200 2062.480 1688.340 ;
        RECT 2067.860 1688.340 2068.000 1688.540 ;
        RECT 2100.890 1688.340 2101.210 1688.400 ;
        RECT 2067.860 1688.200 2101.210 1688.340 ;
        RECT 2021.770 1688.140 2022.090 1688.200 ;
        RECT 2100.890 1688.140 2101.210 1688.200 ;
        RECT 2100.890 19.960 2101.210 20.020 ;
        RECT 2119.750 19.960 2120.070 20.020 ;
        RECT 2100.890 19.820 2120.070 19.960 ;
        RECT 2100.890 19.760 2101.210 19.820 ;
        RECT 2119.750 19.760 2120.070 19.820 ;
      LAYER via ;
        RECT 2021.800 1688.140 2022.060 1688.400 ;
        RECT 2100.920 1688.140 2101.180 1688.400 ;
        RECT 2100.920 19.760 2101.180 20.020 ;
        RECT 2119.780 19.760 2120.040 20.020 ;
      LAYER met2 ;
        RECT 2021.725 1700.000 2022.005 1704.000 ;
        RECT 2021.860 1688.430 2022.000 1700.000 ;
        RECT 2021.800 1688.110 2022.060 1688.430 ;
        RECT 2100.920 1688.110 2101.180 1688.430 ;
        RECT 2100.980 20.050 2101.120 1688.110 ;
        RECT 2100.920 19.730 2101.180 20.050 ;
        RECT 2119.780 19.730 2120.040 20.050 ;
        RECT 2119.840 2.400 2119.980 19.730 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2029.130 1687.320 2029.450 1687.380 ;
        RECT 2132.170 1687.320 2132.490 1687.380 ;
        RECT 2029.130 1687.180 2132.490 1687.320 ;
        RECT 2029.130 1687.120 2029.450 1687.180 ;
        RECT 2132.170 1687.120 2132.490 1687.180 ;
      LAYER via ;
        RECT 2029.160 1687.120 2029.420 1687.380 ;
        RECT 2132.200 1687.120 2132.460 1687.380 ;
      LAYER met2 ;
        RECT 2029.085 1700.000 2029.365 1704.000 ;
        RECT 2029.220 1687.410 2029.360 1700.000 ;
        RECT 2029.160 1687.090 2029.420 1687.410 ;
        RECT 2132.200 1687.090 2132.460 1687.410 ;
        RECT 2132.260 16.730 2132.400 1687.090 ;
        RECT 2132.260 16.590 2137.920 16.730 ;
        RECT 2137.780 2.400 2137.920 16.590 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2130.405 1685.465 2130.575 1687.675 ;
      LAYER mcon ;
        RECT 2130.405 1687.505 2130.575 1687.675 ;
      LAYER met1 ;
        RECT 2036.490 1687.660 2036.810 1687.720 ;
        RECT 2130.345 1687.660 2130.635 1687.705 ;
        RECT 2036.490 1687.520 2130.635 1687.660 ;
        RECT 2036.490 1687.460 2036.810 1687.520 ;
        RECT 2130.345 1687.475 2130.635 1687.520 ;
        RECT 2130.345 1685.620 2130.635 1685.665 ;
        RECT 2135.390 1685.620 2135.710 1685.680 ;
        RECT 2130.345 1685.480 2135.710 1685.620 ;
        RECT 2130.345 1685.435 2130.635 1685.480 ;
        RECT 2135.390 1685.420 2135.710 1685.480 ;
        RECT 2135.390 18.260 2135.710 18.320 ;
        RECT 2155.630 18.260 2155.950 18.320 ;
        RECT 2135.390 18.120 2155.950 18.260 ;
        RECT 2135.390 18.060 2135.710 18.120 ;
        RECT 2155.630 18.060 2155.950 18.120 ;
      LAYER via ;
        RECT 2036.520 1687.460 2036.780 1687.720 ;
        RECT 2135.420 1685.420 2135.680 1685.680 ;
        RECT 2135.420 18.060 2135.680 18.320 ;
        RECT 2155.660 18.060 2155.920 18.320 ;
      LAYER met2 ;
        RECT 2036.445 1700.000 2036.725 1704.000 ;
        RECT 2036.580 1687.750 2036.720 1700.000 ;
        RECT 2036.520 1687.430 2036.780 1687.750 ;
        RECT 2135.420 1685.390 2135.680 1685.710 ;
        RECT 2135.480 18.350 2135.620 1685.390 ;
        RECT 2135.420 18.030 2135.680 18.350 ;
        RECT 2155.660 18.030 2155.920 18.350 ;
        RECT 2155.720 2.400 2155.860 18.030 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2043.850 1688.680 2044.170 1688.740 ;
        RECT 2048.910 1688.680 2049.230 1688.740 ;
        RECT 2043.850 1688.540 2049.230 1688.680 ;
        RECT 2043.850 1688.480 2044.170 1688.540 ;
        RECT 2048.910 1688.480 2049.230 1688.540 ;
        RECT 2048.910 16.900 2049.230 16.960 ;
        RECT 2048.910 16.760 2055.120 16.900 ;
        RECT 2048.910 16.700 2049.230 16.760 ;
        RECT 2054.980 16.560 2055.120 16.760 ;
        RECT 2054.980 16.420 2135.620 16.560 ;
        RECT 2135.480 15.880 2135.620 16.420 ;
        RECT 2173.110 15.880 2173.430 15.940 ;
        RECT 2135.480 15.740 2173.430 15.880 ;
        RECT 2173.110 15.680 2173.430 15.740 ;
      LAYER via ;
        RECT 2043.880 1688.480 2044.140 1688.740 ;
        RECT 2048.940 1688.480 2049.200 1688.740 ;
        RECT 2048.940 16.700 2049.200 16.960 ;
        RECT 2173.140 15.680 2173.400 15.940 ;
      LAYER met2 ;
        RECT 2043.805 1700.000 2044.085 1704.000 ;
        RECT 2043.940 1688.770 2044.080 1700.000 ;
        RECT 2043.880 1688.450 2044.140 1688.770 ;
        RECT 2048.940 1688.450 2049.200 1688.770 ;
        RECT 2049.000 16.990 2049.140 1688.450 ;
        RECT 2048.940 16.670 2049.200 16.990 ;
        RECT 2173.140 15.650 2173.400 15.970 ;
        RECT 2173.200 2.400 2173.340 15.650 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2051.210 1684.600 2051.530 1684.660 ;
        RECT 2055.810 1684.600 2056.130 1684.660 ;
        RECT 2051.210 1684.460 2056.130 1684.600 ;
        RECT 2051.210 1684.400 2051.530 1684.460 ;
        RECT 2055.810 1684.400 2056.130 1684.460 ;
        RECT 2055.810 16.900 2056.130 16.960 ;
        RECT 2191.050 16.900 2191.370 16.960 ;
        RECT 2055.810 16.760 2191.370 16.900 ;
        RECT 2055.810 16.700 2056.130 16.760 ;
        RECT 2191.050 16.700 2191.370 16.760 ;
      LAYER via ;
        RECT 2051.240 1684.400 2051.500 1684.660 ;
        RECT 2055.840 1684.400 2056.100 1684.660 ;
        RECT 2055.840 16.700 2056.100 16.960 ;
        RECT 2191.080 16.700 2191.340 16.960 ;
      LAYER met2 ;
        RECT 2051.165 1700.000 2051.445 1704.000 ;
        RECT 2051.300 1684.690 2051.440 1700.000 ;
        RECT 2051.240 1684.370 2051.500 1684.690 ;
        RECT 2055.840 1684.370 2056.100 1684.690 ;
        RECT 2055.900 16.990 2056.040 1684.370 ;
        RECT 2055.840 16.670 2056.100 16.990 ;
        RECT 2191.080 16.670 2191.340 16.990 ;
        RECT 2191.140 2.400 2191.280 16.670 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2158.005 1685.805 2158.175 1686.995 ;
      LAYER mcon ;
        RECT 2158.005 1686.825 2158.175 1686.995 ;
      LAYER met1 ;
        RECT 2058.570 1686.980 2058.890 1687.040 ;
        RECT 2157.945 1686.980 2158.235 1687.025 ;
        RECT 2058.570 1686.840 2158.235 1686.980 ;
        RECT 2058.570 1686.780 2058.890 1686.840 ;
        RECT 2157.945 1686.795 2158.235 1686.840 ;
        RECT 2157.945 1685.960 2158.235 1686.005 ;
        RECT 2170.350 1685.960 2170.670 1686.020 ;
        RECT 2157.945 1685.820 2170.670 1685.960 ;
        RECT 2157.945 1685.775 2158.235 1685.820 ;
        RECT 2170.350 1685.760 2170.670 1685.820 ;
        RECT 2170.350 16.560 2170.670 16.620 ;
        RECT 2208.990 16.560 2209.310 16.620 ;
        RECT 2170.350 16.420 2209.310 16.560 ;
        RECT 2170.350 16.360 2170.670 16.420 ;
        RECT 2208.990 16.360 2209.310 16.420 ;
      LAYER via ;
        RECT 2058.600 1686.780 2058.860 1687.040 ;
        RECT 2170.380 1685.760 2170.640 1686.020 ;
        RECT 2170.380 16.360 2170.640 16.620 ;
        RECT 2209.020 16.360 2209.280 16.620 ;
      LAYER met2 ;
        RECT 2058.525 1700.000 2058.805 1704.000 ;
        RECT 2058.660 1687.070 2058.800 1700.000 ;
        RECT 2058.600 1686.750 2058.860 1687.070 ;
        RECT 2170.380 1685.730 2170.640 1686.050 ;
        RECT 2170.440 16.650 2170.580 1685.730 ;
        RECT 2170.380 16.330 2170.640 16.650 ;
        RECT 2209.020 16.330 2209.280 16.650 ;
        RECT 2209.080 2.400 2209.220 16.330 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2069.610 18.940 2069.930 19.000 ;
        RECT 2226.930 18.940 2227.250 19.000 ;
        RECT 2069.610 18.800 2227.250 18.940 ;
        RECT 2069.610 18.740 2069.930 18.800 ;
        RECT 2226.930 18.740 2227.250 18.800 ;
      LAYER via ;
        RECT 2069.640 18.740 2069.900 19.000 ;
        RECT 2226.960 18.740 2227.220 19.000 ;
      LAYER met2 ;
        RECT 2065.885 1700.410 2066.165 1704.000 ;
        RECT 2065.885 1700.270 2068.000 1700.410 ;
        RECT 2065.885 1700.000 2066.165 1700.270 ;
        RECT 2067.860 1688.680 2068.000 1700.270 ;
        RECT 2067.860 1688.540 2069.840 1688.680 ;
        RECT 2069.700 19.030 2069.840 1688.540 ;
        RECT 2069.640 18.710 2069.900 19.030 ;
        RECT 2226.960 18.710 2227.220 19.030 ;
        RECT 2227.020 2.400 2227.160 18.710 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 781.610 35.600 781.930 35.660 ;
        RECT 1469.770 35.600 1470.090 35.660 ;
        RECT 781.610 35.460 1470.090 35.600 ;
        RECT 781.610 35.400 781.930 35.460 ;
        RECT 1469.770 35.400 1470.090 35.460 ;
      LAYER via ;
        RECT 781.640 35.400 781.900 35.660 ;
        RECT 1469.800 35.400 1470.060 35.660 ;
      LAYER met2 ;
        RECT 1470.645 1700.410 1470.925 1704.000 ;
        RECT 1469.860 1700.270 1470.925 1700.410 ;
        RECT 1469.860 35.690 1470.000 1700.270 ;
        RECT 1470.645 1700.000 1470.925 1700.270 ;
        RECT 781.640 35.370 781.900 35.690 ;
        RECT 1469.800 35.370 1470.060 35.690 ;
        RECT 781.700 2.400 781.840 35.370 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2169.505 16.065 2174.275 16.235 ;
        RECT 2180.085 14.365 2180.255 16.235 ;
      LAYER mcon ;
        RECT 2174.105 16.065 2174.275 16.235 ;
        RECT 2180.085 16.065 2180.255 16.235 ;
      LAYER met1 ;
        RECT 2073.290 1690.380 2073.610 1690.440 ;
        RECT 2149.190 1690.380 2149.510 1690.440 ;
        RECT 2073.290 1690.240 2149.510 1690.380 ;
        RECT 2073.290 1690.180 2073.610 1690.240 ;
        RECT 2149.190 1690.180 2149.510 1690.240 ;
        RECT 2150.570 16.220 2150.890 16.280 ;
        RECT 2169.445 16.220 2169.735 16.265 ;
        RECT 2150.570 16.080 2169.735 16.220 ;
        RECT 2150.570 16.020 2150.890 16.080 ;
        RECT 2169.445 16.035 2169.735 16.080 ;
        RECT 2174.045 16.220 2174.335 16.265 ;
        RECT 2180.025 16.220 2180.315 16.265 ;
        RECT 2174.045 16.080 2180.315 16.220 ;
        RECT 2174.045 16.035 2174.335 16.080 ;
        RECT 2180.025 16.035 2180.315 16.080 ;
        RECT 2180.025 14.520 2180.315 14.565 ;
        RECT 2244.870 14.520 2245.190 14.580 ;
        RECT 2180.025 14.380 2245.190 14.520 ;
        RECT 2180.025 14.335 2180.315 14.380 ;
        RECT 2244.870 14.320 2245.190 14.380 ;
      LAYER via ;
        RECT 2073.320 1690.180 2073.580 1690.440 ;
        RECT 2149.220 1690.180 2149.480 1690.440 ;
        RECT 2150.600 16.020 2150.860 16.280 ;
        RECT 2244.900 14.320 2245.160 14.580 ;
      LAYER met2 ;
        RECT 2073.245 1700.000 2073.525 1704.000 ;
        RECT 2073.380 1690.470 2073.520 1700.000 ;
        RECT 2073.320 1690.150 2073.580 1690.470 ;
        RECT 2149.220 1690.150 2149.480 1690.470 ;
        RECT 2149.280 38.490 2149.420 1690.150 ;
        RECT 2149.280 38.350 2150.800 38.490 ;
        RECT 2150.660 16.310 2150.800 38.350 ;
        RECT 2150.600 15.990 2150.860 16.310 ;
        RECT 2244.900 14.290 2245.160 14.610 ;
        RECT 2244.960 2.400 2245.100 14.290 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2140.525 15.045 2140.695 18.615 ;
      LAYER mcon ;
        RECT 2140.525 18.445 2140.695 18.615 ;
      LAYER met1 ;
        RECT 2140.465 18.600 2140.755 18.645 ;
        RECT 2262.350 18.600 2262.670 18.660 ;
        RECT 2140.465 18.460 2156.320 18.600 ;
        RECT 2140.465 18.415 2140.755 18.460 ;
        RECT 2156.180 18.260 2156.320 18.460 ;
        RECT 2232.080 18.460 2262.670 18.600 ;
        RECT 2232.080 18.260 2232.220 18.460 ;
        RECT 2262.350 18.400 2262.670 18.460 ;
        RECT 2156.180 18.120 2232.220 18.260 ;
        RECT 2083.410 15.200 2083.730 15.260 ;
        RECT 2140.465 15.200 2140.755 15.245 ;
        RECT 2083.410 15.060 2140.755 15.200 ;
        RECT 2083.410 15.000 2083.730 15.060 ;
        RECT 2140.465 15.015 2140.755 15.060 ;
      LAYER via ;
        RECT 2262.380 18.400 2262.640 18.660 ;
        RECT 2083.440 15.000 2083.700 15.260 ;
      LAYER met2 ;
        RECT 2080.605 1700.410 2080.885 1704.000 ;
        RECT 2080.605 1700.270 2082.720 1700.410 ;
        RECT 2080.605 1700.000 2080.885 1700.270 ;
        RECT 2082.580 1688.680 2082.720 1700.270 ;
        RECT 2082.580 1688.540 2083.640 1688.680 ;
        RECT 2083.500 15.290 2083.640 1688.540 ;
        RECT 2262.380 18.370 2262.640 18.690 ;
        RECT 2083.440 14.970 2083.700 15.290 ;
        RECT 2262.440 2.400 2262.580 18.370 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2088.010 1689.360 2088.330 1689.420 ;
        RECT 2277.990 1689.360 2278.310 1689.420 ;
        RECT 2088.010 1689.220 2278.310 1689.360 ;
        RECT 2088.010 1689.160 2088.330 1689.220 ;
        RECT 2277.990 1689.160 2278.310 1689.220 ;
      LAYER via ;
        RECT 2088.040 1689.160 2088.300 1689.420 ;
        RECT 2278.020 1689.160 2278.280 1689.420 ;
      LAYER met2 ;
        RECT 2087.965 1700.000 2088.245 1704.000 ;
        RECT 2088.100 1689.450 2088.240 1700.000 ;
        RECT 2088.040 1689.130 2088.300 1689.450 ;
        RECT 2278.020 1689.130 2278.280 1689.450 ;
        RECT 2278.080 10.610 2278.220 1689.130 ;
        RECT 2278.080 10.470 2280.060 10.610 ;
        RECT 2279.920 3.130 2280.060 10.470 ;
        RECT 2279.920 2.990 2280.520 3.130 ;
        RECT 2280.380 2.400 2280.520 2.990 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2156.625 386.325 2156.795 434.775 ;
        RECT 2156.625 338.045 2156.795 385.815 ;
      LAYER mcon ;
        RECT 2156.625 434.605 2156.795 434.775 ;
        RECT 2156.625 385.645 2156.795 385.815 ;
      LAYER met1 ;
        RECT 2157.470 1685.960 2157.790 1686.020 ;
        RECT 2129.960 1685.820 2157.790 1685.960 ;
        RECT 2095.370 1685.620 2095.690 1685.680 ;
        RECT 2129.960 1685.620 2130.100 1685.820 ;
        RECT 2157.470 1685.760 2157.790 1685.820 ;
        RECT 2095.370 1685.480 2130.100 1685.620 ;
        RECT 2095.370 1685.420 2095.690 1685.480 ;
        RECT 2157.010 1594.160 2157.330 1594.220 ;
        RECT 2157.470 1594.160 2157.790 1594.220 ;
        RECT 2157.010 1594.020 2157.790 1594.160 ;
        RECT 2157.010 1593.960 2157.330 1594.020 ;
        RECT 2157.470 1593.960 2157.790 1594.020 ;
        RECT 2157.010 1559.820 2157.330 1559.880 ;
        RECT 2157.470 1559.820 2157.790 1559.880 ;
        RECT 2157.010 1559.680 2157.790 1559.820 ;
        RECT 2157.010 1559.620 2157.330 1559.680 ;
        RECT 2157.470 1559.620 2157.790 1559.680 ;
        RECT 2156.550 1511.200 2156.870 1511.260 ;
        RECT 2157.470 1511.200 2157.790 1511.260 ;
        RECT 2156.550 1511.060 2157.790 1511.200 ;
        RECT 2156.550 1511.000 2156.870 1511.060 ;
        RECT 2157.470 1511.000 2157.790 1511.060 ;
        RECT 2156.550 1414.640 2156.870 1414.700 ;
        RECT 2157.470 1414.640 2157.790 1414.700 ;
        RECT 2156.550 1414.500 2157.790 1414.640 ;
        RECT 2156.550 1414.440 2156.870 1414.500 ;
        RECT 2157.470 1414.440 2157.790 1414.500 ;
        RECT 2156.550 1318.080 2156.870 1318.140 ;
        RECT 2157.470 1318.080 2157.790 1318.140 ;
        RECT 2156.550 1317.940 2157.790 1318.080 ;
        RECT 2156.550 1317.880 2156.870 1317.940 ;
        RECT 2157.470 1317.880 2157.790 1317.940 ;
        RECT 2156.550 1221.520 2156.870 1221.580 ;
        RECT 2157.470 1221.520 2157.790 1221.580 ;
        RECT 2156.550 1221.380 2157.790 1221.520 ;
        RECT 2156.550 1221.320 2156.870 1221.380 ;
        RECT 2157.470 1221.320 2157.790 1221.380 ;
        RECT 2156.550 1124.960 2156.870 1125.020 ;
        RECT 2157.470 1124.960 2157.790 1125.020 ;
        RECT 2156.550 1124.820 2157.790 1124.960 ;
        RECT 2156.550 1124.760 2156.870 1124.820 ;
        RECT 2157.470 1124.760 2157.790 1124.820 ;
        RECT 2156.550 1028.400 2156.870 1028.460 ;
        RECT 2157.470 1028.400 2157.790 1028.460 ;
        RECT 2156.550 1028.260 2157.790 1028.400 ;
        RECT 2156.550 1028.200 2156.870 1028.260 ;
        RECT 2157.470 1028.200 2157.790 1028.260 ;
        RECT 2156.550 931.840 2156.870 931.900 ;
        RECT 2157.470 931.840 2157.790 931.900 ;
        RECT 2156.550 931.700 2157.790 931.840 ;
        RECT 2156.550 931.640 2156.870 931.700 ;
        RECT 2157.470 931.640 2157.790 931.700 ;
        RECT 2156.550 835.280 2156.870 835.340 ;
        RECT 2157.470 835.280 2157.790 835.340 ;
        RECT 2156.550 835.140 2157.790 835.280 ;
        RECT 2156.550 835.080 2156.870 835.140 ;
        RECT 2157.470 835.080 2157.790 835.140 ;
        RECT 2156.550 448.700 2156.870 448.760 ;
        RECT 2157.470 448.700 2157.790 448.760 ;
        RECT 2156.550 448.560 2157.790 448.700 ;
        RECT 2156.550 448.500 2156.870 448.560 ;
        RECT 2157.470 448.500 2157.790 448.560 ;
        RECT 2156.550 434.760 2156.870 434.820 ;
        RECT 2156.355 434.620 2156.870 434.760 ;
        RECT 2156.550 434.560 2156.870 434.620 ;
        RECT 2156.550 386.480 2156.870 386.540 ;
        RECT 2156.355 386.340 2156.870 386.480 ;
        RECT 2156.550 386.280 2156.870 386.340 ;
        RECT 2156.550 385.800 2156.870 385.860 ;
        RECT 2156.355 385.660 2156.870 385.800 ;
        RECT 2156.550 385.600 2156.870 385.660 ;
        RECT 2156.565 338.200 2156.855 338.245 ;
        RECT 2157.010 338.200 2157.330 338.260 ;
        RECT 2156.565 338.060 2157.330 338.200 ;
        RECT 2156.565 338.015 2156.855 338.060 ;
        RECT 2157.010 338.000 2157.330 338.060 ;
        RECT 2298.230 14.860 2298.550 14.920 ;
        RECT 2162.160 14.720 2298.550 14.860 ;
        RECT 2156.550 14.520 2156.870 14.580 ;
        RECT 2162.160 14.520 2162.300 14.720 ;
        RECT 2298.230 14.660 2298.550 14.720 ;
        RECT 2156.550 14.380 2162.300 14.520 ;
        RECT 2156.550 14.320 2156.870 14.380 ;
      LAYER via ;
        RECT 2095.400 1685.420 2095.660 1685.680 ;
        RECT 2157.500 1685.760 2157.760 1686.020 ;
        RECT 2157.040 1593.960 2157.300 1594.220 ;
        RECT 2157.500 1593.960 2157.760 1594.220 ;
        RECT 2157.040 1559.620 2157.300 1559.880 ;
        RECT 2157.500 1559.620 2157.760 1559.880 ;
        RECT 2156.580 1511.000 2156.840 1511.260 ;
        RECT 2157.500 1511.000 2157.760 1511.260 ;
        RECT 2156.580 1414.440 2156.840 1414.700 ;
        RECT 2157.500 1414.440 2157.760 1414.700 ;
        RECT 2156.580 1317.880 2156.840 1318.140 ;
        RECT 2157.500 1317.880 2157.760 1318.140 ;
        RECT 2156.580 1221.320 2156.840 1221.580 ;
        RECT 2157.500 1221.320 2157.760 1221.580 ;
        RECT 2156.580 1124.760 2156.840 1125.020 ;
        RECT 2157.500 1124.760 2157.760 1125.020 ;
        RECT 2156.580 1028.200 2156.840 1028.460 ;
        RECT 2157.500 1028.200 2157.760 1028.460 ;
        RECT 2156.580 931.640 2156.840 931.900 ;
        RECT 2157.500 931.640 2157.760 931.900 ;
        RECT 2156.580 835.080 2156.840 835.340 ;
        RECT 2157.500 835.080 2157.760 835.340 ;
        RECT 2156.580 448.500 2156.840 448.760 ;
        RECT 2157.500 448.500 2157.760 448.760 ;
        RECT 2156.580 434.560 2156.840 434.820 ;
        RECT 2156.580 386.280 2156.840 386.540 ;
        RECT 2156.580 385.600 2156.840 385.860 ;
        RECT 2157.040 338.000 2157.300 338.260 ;
        RECT 2156.580 14.320 2156.840 14.580 ;
        RECT 2298.260 14.660 2298.520 14.920 ;
      LAYER met2 ;
        RECT 2095.325 1700.000 2095.605 1704.000 ;
        RECT 2095.460 1685.710 2095.600 1700.000 ;
        RECT 2157.500 1685.730 2157.760 1686.050 ;
        RECT 2095.400 1685.390 2095.660 1685.710 ;
        RECT 2157.560 1594.250 2157.700 1685.730 ;
        RECT 2157.040 1593.930 2157.300 1594.250 ;
        RECT 2157.500 1593.930 2157.760 1594.250 ;
        RECT 2157.100 1559.910 2157.240 1593.930 ;
        RECT 2157.040 1559.590 2157.300 1559.910 ;
        RECT 2157.500 1559.590 2157.760 1559.910 ;
        RECT 2157.560 1511.290 2157.700 1559.590 ;
        RECT 2156.580 1510.970 2156.840 1511.290 ;
        RECT 2157.500 1510.970 2157.760 1511.290 ;
        RECT 2156.640 1510.690 2156.780 1510.970 ;
        RECT 2156.640 1510.550 2157.240 1510.690 ;
        RECT 2157.100 1463.090 2157.240 1510.550 ;
        RECT 2157.100 1462.950 2157.700 1463.090 ;
        RECT 2157.560 1414.730 2157.700 1462.950 ;
        RECT 2156.580 1414.410 2156.840 1414.730 ;
        RECT 2157.500 1414.410 2157.760 1414.730 ;
        RECT 2156.640 1414.130 2156.780 1414.410 ;
        RECT 2156.640 1413.990 2157.240 1414.130 ;
        RECT 2157.100 1366.530 2157.240 1413.990 ;
        RECT 2157.100 1366.390 2157.700 1366.530 ;
        RECT 2157.560 1318.170 2157.700 1366.390 ;
        RECT 2156.580 1317.850 2156.840 1318.170 ;
        RECT 2157.500 1317.850 2157.760 1318.170 ;
        RECT 2156.640 1317.570 2156.780 1317.850 ;
        RECT 2156.640 1317.430 2157.240 1317.570 ;
        RECT 2157.100 1269.970 2157.240 1317.430 ;
        RECT 2157.100 1269.830 2157.700 1269.970 ;
        RECT 2157.560 1221.610 2157.700 1269.830 ;
        RECT 2156.580 1221.290 2156.840 1221.610 ;
        RECT 2157.500 1221.290 2157.760 1221.610 ;
        RECT 2156.640 1221.010 2156.780 1221.290 ;
        RECT 2156.640 1220.870 2157.240 1221.010 ;
        RECT 2157.100 1173.410 2157.240 1220.870 ;
        RECT 2157.100 1173.270 2157.700 1173.410 ;
        RECT 2157.560 1125.050 2157.700 1173.270 ;
        RECT 2156.580 1124.730 2156.840 1125.050 ;
        RECT 2157.500 1124.730 2157.760 1125.050 ;
        RECT 2156.640 1124.450 2156.780 1124.730 ;
        RECT 2156.640 1124.310 2157.240 1124.450 ;
        RECT 2157.100 1076.850 2157.240 1124.310 ;
        RECT 2157.100 1076.710 2157.700 1076.850 ;
        RECT 2157.560 1028.490 2157.700 1076.710 ;
        RECT 2156.580 1028.170 2156.840 1028.490 ;
        RECT 2157.500 1028.170 2157.760 1028.490 ;
        RECT 2156.640 1027.890 2156.780 1028.170 ;
        RECT 2156.640 1027.750 2157.240 1027.890 ;
        RECT 2157.100 980.290 2157.240 1027.750 ;
        RECT 2157.100 980.150 2157.700 980.290 ;
        RECT 2157.560 931.930 2157.700 980.150 ;
        RECT 2156.580 931.610 2156.840 931.930 ;
        RECT 2157.500 931.610 2157.760 931.930 ;
        RECT 2156.640 883.050 2156.780 931.610 ;
        RECT 2156.640 882.910 2157.700 883.050 ;
        RECT 2157.560 835.370 2157.700 882.910 ;
        RECT 2156.580 835.050 2156.840 835.370 ;
        RECT 2157.500 835.050 2157.760 835.370 ;
        RECT 2156.640 496.810 2156.780 835.050 ;
        RECT 2156.640 496.670 2157.700 496.810 ;
        RECT 2157.560 448.790 2157.700 496.670 ;
        RECT 2156.580 448.470 2156.840 448.790 ;
        RECT 2157.500 448.470 2157.760 448.790 ;
        RECT 2156.640 434.850 2156.780 448.470 ;
        RECT 2156.580 434.530 2156.840 434.850 ;
        RECT 2156.580 386.250 2156.840 386.570 ;
        RECT 2156.640 385.890 2156.780 386.250 ;
        RECT 2156.580 385.570 2156.840 385.890 ;
        RECT 2157.040 337.970 2157.300 338.290 ;
        RECT 2157.100 303.690 2157.240 337.970 ;
        RECT 2157.100 303.550 2157.700 303.690 ;
        RECT 2157.560 255.410 2157.700 303.550 ;
        RECT 2156.640 255.270 2157.700 255.410 ;
        RECT 2156.640 14.610 2156.780 255.270 ;
        RECT 2298.260 14.630 2298.520 14.950 ;
        RECT 2156.580 14.290 2156.840 14.610 ;
        RECT 2298.320 2.400 2298.460 14.630 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2111.545 1687.845 2111.715 1690.055 ;
        RECT 2201.705 1686.825 2201.875 1689.715 ;
        RECT 2209.525 1687.165 2209.695 1689.715 ;
        RECT 2255.525 1687.165 2255.695 1690.055 ;
        RECT 2273.465 1684.105 2273.635 1690.055 ;
        RECT 2301.065 1538.925 2301.235 1587.035 ;
        RECT 2300.145 1442.025 2300.315 1490.475 ;
        RECT 2300.605 1365.525 2300.775 1400.715 ;
        RECT 2300.145 1304.665 2300.315 1352.435 ;
        RECT 2300.145 1207.425 2300.315 1255.875 ;
        RECT 2300.605 882.385 2300.775 917.575 ;
        RECT 2300.145 241.485 2300.315 289.595 ;
        RECT 2300.145 206.805 2300.315 240.975 ;
        RECT 2300.605 158.525 2300.775 193.035 ;
      LAYER mcon ;
        RECT 2111.545 1689.885 2111.715 1690.055 ;
        RECT 2255.525 1689.885 2255.695 1690.055 ;
        RECT 2201.705 1689.545 2201.875 1689.715 ;
        RECT 2209.525 1689.545 2209.695 1689.715 ;
        RECT 2273.465 1689.885 2273.635 1690.055 ;
        RECT 2301.065 1586.865 2301.235 1587.035 ;
        RECT 2300.145 1490.305 2300.315 1490.475 ;
        RECT 2300.605 1400.545 2300.775 1400.715 ;
        RECT 2300.145 1352.265 2300.315 1352.435 ;
        RECT 2300.145 1255.705 2300.315 1255.875 ;
        RECT 2300.605 917.405 2300.775 917.575 ;
        RECT 2300.145 289.425 2300.315 289.595 ;
        RECT 2300.145 240.805 2300.315 240.975 ;
        RECT 2300.605 192.865 2300.775 193.035 ;
      LAYER met1 ;
        RECT 2102.730 1690.040 2103.050 1690.100 ;
        RECT 2111.485 1690.040 2111.775 1690.085 ;
        RECT 2102.730 1689.900 2111.775 1690.040 ;
        RECT 2102.730 1689.840 2103.050 1689.900 ;
        RECT 2111.485 1689.855 2111.775 1689.900 ;
        RECT 2255.465 1690.040 2255.755 1690.085 ;
        RECT 2273.405 1690.040 2273.695 1690.085 ;
        RECT 2255.465 1689.900 2273.695 1690.040 ;
        RECT 2255.465 1689.855 2255.755 1689.900 ;
        RECT 2273.405 1689.855 2273.695 1689.900 ;
        RECT 2201.645 1689.700 2201.935 1689.745 ;
        RECT 2209.465 1689.700 2209.755 1689.745 ;
        RECT 2201.645 1689.560 2209.755 1689.700 ;
        RECT 2201.645 1689.515 2201.935 1689.560 ;
        RECT 2209.465 1689.515 2209.755 1689.560 ;
        RECT 2111.485 1688.000 2111.775 1688.045 ;
        RECT 2111.485 1687.860 2132.860 1688.000 ;
        RECT 2111.485 1687.815 2111.775 1687.860 ;
        RECT 2132.720 1687.320 2132.860 1687.860 ;
        RECT 2218.740 1687.860 2243.260 1688.000 ;
        RECT 2218.740 1687.660 2218.880 1687.860 ;
        RECT 2212.300 1687.520 2218.880 1687.660 ;
        RECT 2209.465 1687.320 2209.755 1687.365 ;
        RECT 2212.300 1687.320 2212.440 1687.520 ;
        RECT 2132.720 1687.180 2163.220 1687.320 ;
        RECT 2163.080 1686.980 2163.220 1687.180 ;
        RECT 2209.465 1687.180 2212.440 1687.320 ;
        RECT 2243.120 1687.320 2243.260 1687.860 ;
        RECT 2255.465 1687.320 2255.755 1687.365 ;
        RECT 2243.120 1687.180 2255.755 1687.320 ;
        RECT 2209.465 1687.135 2209.755 1687.180 ;
        RECT 2255.465 1687.135 2255.755 1687.180 ;
        RECT 2201.645 1686.980 2201.935 1687.025 ;
        RECT 2163.080 1686.840 2201.935 1686.980 ;
        RECT 2201.645 1686.795 2201.935 1686.840 ;
        RECT 2273.405 1684.260 2273.695 1684.305 ;
        RECT 2298.230 1684.260 2298.550 1684.320 ;
        RECT 2273.405 1684.120 2298.550 1684.260 ;
        RECT 2273.405 1684.075 2273.695 1684.120 ;
        RECT 2298.230 1684.060 2298.550 1684.120 ;
        RECT 2298.230 1656.040 2298.550 1656.100 ;
        RECT 2300.530 1656.040 2300.850 1656.100 ;
        RECT 2298.230 1655.900 2300.850 1656.040 ;
        RECT 2298.230 1655.840 2298.550 1655.900 ;
        RECT 2300.530 1655.840 2300.850 1655.900 ;
        RECT 2300.990 1587.020 2301.310 1587.080 ;
        RECT 2300.795 1586.880 2301.310 1587.020 ;
        RECT 2300.990 1586.820 2301.310 1586.880 ;
        RECT 2300.990 1539.080 2301.310 1539.140 ;
        RECT 2300.795 1538.940 2301.310 1539.080 ;
        RECT 2300.990 1538.880 2301.310 1538.940 ;
        RECT 2300.070 1490.460 2300.390 1490.520 ;
        RECT 2299.875 1490.320 2300.390 1490.460 ;
        RECT 2300.070 1490.260 2300.390 1490.320 ;
        RECT 2300.085 1442.180 2300.375 1442.225 ;
        RECT 2300.530 1442.180 2300.850 1442.240 ;
        RECT 2300.085 1442.040 2300.850 1442.180 ;
        RECT 2300.085 1441.995 2300.375 1442.040 ;
        RECT 2300.530 1441.980 2300.850 1442.040 ;
        RECT 2300.530 1414.780 2300.850 1415.040 ;
        RECT 2300.620 1414.020 2300.760 1414.780 ;
        RECT 2300.530 1413.760 2300.850 1414.020 ;
        RECT 2300.530 1400.700 2300.850 1400.760 ;
        RECT 2300.335 1400.560 2300.850 1400.700 ;
        RECT 2300.530 1400.500 2300.850 1400.560 ;
        RECT 2300.530 1365.680 2300.850 1365.740 ;
        RECT 2300.335 1365.540 2300.850 1365.680 ;
        RECT 2300.530 1365.480 2300.850 1365.540 ;
        RECT 2300.085 1352.420 2300.375 1352.465 ;
        RECT 2300.530 1352.420 2300.850 1352.480 ;
        RECT 2300.085 1352.280 2300.850 1352.420 ;
        RECT 2300.085 1352.235 2300.375 1352.280 ;
        RECT 2300.530 1352.220 2300.850 1352.280 ;
        RECT 2300.070 1304.820 2300.390 1304.880 ;
        RECT 2299.875 1304.680 2300.390 1304.820 ;
        RECT 2300.070 1304.620 2300.390 1304.680 ;
        RECT 2300.070 1304.140 2300.390 1304.200 ;
        RECT 2300.990 1304.140 2301.310 1304.200 ;
        RECT 2300.070 1304.000 2301.310 1304.140 ;
        RECT 2300.070 1303.940 2300.390 1304.000 ;
        RECT 2300.990 1303.940 2301.310 1304.000 ;
        RECT 2300.085 1255.860 2300.375 1255.905 ;
        RECT 2300.530 1255.860 2300.850 1255.920 ;
        RECT 2300.085 1255.720 2300.850 1255.860 ;
        RECT 2300.085 1255.675 2300.375 1255.720 ;
        RECT 2300.530 1255.660 2300.850 1255.720 ;
        RECT 2300.070 1207.580 2300.390 1207.640 ;
        RECT 2299.875 1207.440 2300.390 1207.580 ;
        RECT 2300.070 1207.380 2300.390 1207.440 ;
        RECT 2300.530 1125.300 2300.850 1125.360 ;
        RECT 2300.160 1125.160 2300.850 1125.300 ;
        RECT 2300.160 1124.680 2300.300 1125.160 ;
        RECT 2300.530 1125.100 2300.850 1125.160 ;
        RECT 2300.070 1124.420 2300.390 1124.680 ;
        RECT 2299.150 1076.340 2299.470 1076.400 ;
        RECT 2300.070 1076.340 2300.390 1076.400 ;
        RECT 2299.150 1076.200 2300.390 1076.340 ;
        RECT 2299.150 1076.140 2299.470 1076.200 ;
        RECT 2300.070 1076.140 2300.390 1076.200 ;
        RECT 2300.530 1028.740 2300.850 1028.800 ;
        RECT 2300.160 1028.600 2300.850 1028.740 ;
        RECT 2300.160 1028.120 2300.300 1028.600 ;
        RECT 2300.530 1028.540 2300.850 1028.600 ;
        RECT 2300.070 1027.860 2300.390 1028.120 ;
        RECT 2300.070 979.920 2300.390 980.180 ;
        RECT 2300.160 979.440 2300.300 979.920 ;
        RECT 2300.530 979.440 2300.850 979.500 ;
        RECT 2300.160 979.300 2300.850 979.440 ;
        RECT 2300.530 979.240 2300.850 979.300 ;
        RECT 2300.070 931.840 2300.390 931.900 ;
        RECT 2300.070 931.700 2300.760 931.840 ;
        RECT 2300.070 931.640 2300.390 931.700 ;
        RECT 2300.620 931.560 2300.760 931.700 ;
        RECT 2300.530 931.300 2300.850 931.560 ;
        RECT 2300.530 917.560 2300.850 917.620 ;
        RECT 2300.335 917.420 2300.850 917.560 ;
        RECT 2300.530 917.360 2300.850 917.420 ;
        RECT 2300.530 882.540 2300.850 882.600 ;
        RECT 2300.335 882.400 2300.850 882.540 ;
        RECT 2300.530 882.340 2300.850 882.400 ;
        RECT 2300.990 787.340 2301.310 787.400 ;
        RECT 2300.160 787.200 2301.310 787.340 ;
        RECT 2300.160 786.720 2300.300 787.200 ;
        RECT 2300.990 787.140 2301.310 787.200 ;
        RECT 2300.070 786.460 2300.390 786.720 ;
        RECT 2299.610 724.440 2299.930 724.500 ;
        RECT 2300.990 724.440 2301.310 724.500 ;
        RECT 2299.610 724.300 2301.310 724.440 ;
        RECT 2299.610 724.240 2299.930 724.300 ;
        RECT 2300.990 724.240 2301.310 724.300 ;
        RECT 2299.610 531.320 2299.930 531.380 ;
        RECT 2300.530 531.320 2300.850 531.380 ;
        RECT 2299.610 531.180 2300.850 531.320 ;
        RECT 2299.610 531.120 2299.930 531.180 ;
        RECT 2300.530 531.120 2300.850 531.180 ;
        RECT 2299.610 337.860 2299.930 337.920 ;
        RECT 2300.990 337.860 2301.310 337.920 ;
        RECT 2299.610 337.720 2301.310 337.860 ;
        RECT 2299.610 337.660 2299.930 337.720 ;
        RECT 2300.990 337.660 2301.310 337.720 ;
        RECT 2300.085 289.580 2300.375 289.625 ;
        RECT 2300.530 289.580 2300.850 289.640 ;
        RECT 2300.085 289.440 2300.850 289.580 ;
        RECT 2300.085 289.395 2300.375 289.440 ;
        RECT 2300.530 289.380 2300.850 289.440 ;
        RECT 2300.070 241.640 2300.390 241.700 ;
        RECT 2299.875 241.500 2300.390 241.640 ;
        RECT 2300.070 241.440 2300.390 241.500 ;
        RECT 2300.070 240.960 2300.390 241.020 ;
        RECT 2299.875 240.820 2300.390 240.960 ;
        RECT 2300.070 240.760 2300.390 240.820 ;
        RECT 2300.085 206.960 2300.375 207.005 ;
        RECT 2300.990 206.960 2301.310 207.020 ;
        RECT 2300.085 206.820 2301.310 206.960 ;
        RECT 2300.085 206.775 2300.375 206.820 ;
        RECT 2300.990 206.760 2301.310 206.820 ;
        RECT 2300.545 193.020 2300.835 193.065 ;
        RECT 2300.990 193.020 2301.310 193.080 ;
        RECT 2300.545 192.880 2301.310 193.020 ;
        RECT 2300.545 192.835 2300.835 192.880 ;
        RECT 2300.990 192.820 2301.310 192.880 ;
        RECT 2300.530 158.680 2300.850 158.740 ;
        RECT 2300.335 158.540 2300.850 158.680 ;
        RECT 2300.530 158.480 2300.850 158.540 ;
        RECT 2300.530 110.060 2300.850 110.120 ;
        RECT 2301.910 110.060 2302.230 110.120 ;
        RECT 2300.530 109.920 2302.230 110.060 ;
        RECT 2300.530 109.860 2300.850 109.920 ;
        RECT 2301.910 109.860 2302.230 109.920 ;
        RECT 2301.910 18.940 2302.230 19.000 ;
        RECT 2316.170 18.940 2316.490 19.000 ;
        RECT 2301.910 18.800 2316.490 18.940 ;
        RECT 2301.910 18.740 2302.230 18.800 ;
        RECT 2316.170 18.740 2316.490 18.800 ;
      LAYER via ;
        RECT 2102.760 1689.840 2103.020 1690.100 ;
        RECT 2298.260 1684.060 2298.520 1684.320 ;
        RECT 2298.260 1655.840 2298.520 1656.100 ;
        RECT 2300.560 1655.840 2300.820 1656.100 ;
        RECT 2301.020 1586.820 2301.280 1587.080 ;
        RECT 2301.020 1538.880 2301.280 1539.140 ;
        RECT 2300.100 1490.260 2300.360 1490.520 ;
        RECT 2300.560 1441.980 2300.820 1442.240 ;
        RECT 2300.560 1414.780 2300.820 1415.040 ;
        RECT 2300.560 1413.760 2300.820 1414.020 ;
        RECT 2300.560 1400.500 2300.820 1400.760 ;
        RECT 2300.560 1365.480 2300.820 1365.740 ;
        RECT 2300.560 1352.220 2300.820 1352.480 ;
        RECT 2300.100 1304.620 2300.360 1304.880 ;
        RECT 2300.100 1303.940 2300.360 1304.200 ;
        RECT 2301.020 1303.940 2301.280 1304.200 ;
        RECT 2300.560 1255.660 2300.820 1255.920 ;
        RECT 2300.100 1207.380 2300.360 1207.640 ;
        RECT 2300.560 1125.100 2300.820 1125.360 ;
        RECT 2300.100 1124.420 2300.360 1124.680 ;
        RECT 2299.180 1076.140 2299.440 1076.400 ;
        RECT 2300.100 1076.140 2300.360 1076.400 ;
        RECT 2300.560 1028.540 2300.820 1028.800 ;
        RECT 2300.100 1027.860 2300.360 1028.120 ;
        RECT 2300.100 979.920 2300.360 980.180 ;
        RECT 2300.560 979.240 2300.820 979.500 ;
        RECT 2300.100 931.640 2300.360 931.900 ;
        RECT 2300.560 931.300 2300.820 931.560 ;
        RECT 2300.560 917.360 2300.820 917.620 ;
        RECT 2300.560 882.340 2300.820 882.600 ;
        RECT 2301.020 787.140 2301.280 787.400 ;
        RECT 2300.100 786.460 2300.360 786.720 ;
        RECT 2299.640 724.240 2299.900 724.500 ;
        RECT 2301.020 724.240 2301.280 724.500 ;
        RECT 2299.640 531.120 2299.900 531.380 ;
        RECT 2300.560 531.120 2300.820 531.380 ;
        RECT 2299.640 337.660 2299.900 337.920 ;
        RECT 2301.020 337.660 2301.280 337.920 ;
        RECT 2300.560 289.380 2300.820 289.640 ;
        RECT 2300.100 241.440 2300.360 241.700 ;
        RECT 2300.100 240.760 2300.360 241.020 ;
        RECT 2301.020 206.760 2301.280 207.020 ;
        RECT 2301.020 192.820 2301.280 193.080 ;
        RECT 2300.560 158.480 2300.820 158.740 ;
        RECT 2300.560 109.860 2300.820 110.120 ;
        RECT 2301.940 109.860 2302.200 110.120 ;
        RECT 2301.940 18.740 2302.200 19.000 ;
        RECT 2316.200 18.740 2316.460 19.000 ;
      LAYER met2 ;
        RECT 2102.685 1700.000 2102.965 1704.000 ;
        RECT 2102.820 1690.130 2102.960 1700.000 ;
        RECT 2102.760 1689.810 2103.020 1690.130 ;
        RECT 2298.260 1684.030 2298.520 1684.350 ;
        RECT 2298.320 1656.130 2298.460 1684.030 ;
        RECT 2298.260 1655.810 2298.520 1656.130 ;
        RECT 2300.560 1655.810 2300.820 1656.130 ;
        RECT 2300.620 1618.130 2300.760 1655.810 ;
        RECT 2300.160 1617.990 2300.760 1618.130 ;
        RECT 2300.160 1594.445 2300.300 1617.990 ;
        RECT 2300.090 1594.075 2300.370 1594.445 ;
        RECT 2301.010 1594.075 2301.290 1594.445 ;
        RECT 2301.080 1587.110 2301.220 1594.075 ;
        RECT 2301.020 1586.790 2301.280 1587.110 ;
        RECT 2301.020 1538.850 2301.280 1539.170 ;
        RECT 2301.080 1512.050 2301.220 1538.850 ;
        RECT 2300.620 1511.910 2301.220 1512.050 ;
        RECT 2300.620 1497.770 2300.760 1511.910 ;
        RECT 2300.160 1497.630 2300.760 1497.770 ;
        RECT 2300.160 1490.550 2300.300 1497.630 ;
        RECT 2300.100 1490.230 2300.360 1490.550 ;
        RECT 2300.560 1441.950 2300.820 1442.270 ;
        RECT 2300.620 1415.070 2300.760 1441.950 ;
        RECT 2300.560 1414.750 2300.820 1415.070 ;
        RECT 2300.560 1413.730 2300.820 1414.050 ;
        RECT 2300.620 1400.790 2300.760 1413.730 ;
        RECT 2300.560 1400.470 2300.820 1400.790 ;
        RECT 2300.560 1365.450 2300.820 1365.770 ;
        RECT 2300.620 1352.510 2300.760 1365.450 ;
        RECT 2300.560 1352.190 2300.820 1352.510 ;
        RECT 2300.100 1304.590 2300.360 1304.910 ;
        RECT 2300.160 1304.230 2300.300 1304.590 ;
        RECT 2300.100 1303.910 2300.360 1304.230 ;
        RECT 2301.020 1303.910 2301.280 1304.230 ;
        RECT 2301.080 1269.290 2301.220 1303.910 ;
        RECT 2300.620 1269.150 2301.220 1269.290 ;
        RECT 2300.620 1255.950 2300.760 1269.150 ;
        RECT 2300.560 1255.630 2300.820 1255.950 ;
        RECT 2300.100 1207.525 2300.360 1207.670 ;
        RECT 2300.090 1207.155 2300.370 1207.525 ;
        RECT 2300.550 1172.475 2300.830 1172.845 ;
        RECT 2300.620 1125.390 2300.760 1172.475 ;
        RECT 2300.560 1125.070 2300.820 1125.390 ;
        RECT 2300.100 1124.390 2300.360 1124.710 ;
        RECT 2300.160 1104.165 2300.300 1124.390 ;
        RECT 2299.170 1103.795 2299.450 1104.165 ;
        RECT 2300.090 1103.795 2300.370 1104.165 ;
        RECT 2299.240 1076.430 2299.380 1103.795 ;
        RECT 2299.180 1076.110 2299.440 1076.430 ;
        RECT 2300.100 1076.110 2300.360 1076.430 ;
        RECT 2300.160 1055.770 2300.300 1076.110 ;
        RECT 2300.160 1055.630 2300.760 1055.770 ;
        RECT 2300.620 1028.830 2300.760 1055.630 ;
        RECT 2300.560 1028.510 2300.820 1028.830 ;
        RECT 2300.100 1027.830 2300.360 1028.150 ;
        RECT 2300.160 980.210 2300.300 1027.830 ;
        RECT 2300.100 979.890 2300.360 980.210 ;
        RECT 2300.560 979.210 2300.820 979.530 ;
        RECT 2300.620 966.010 2300.760 979.210 ;
        RECT 2300.160 965.870 2300.760 966.010 ;
        RECT 2300.160 931.930 2300.300 965.870 ;
        RECT 2300.100 931.610 2300.360 931.930 ;
        RECT 2300.560 931.270 2300.820 931.590 ;
        RECT 2300.620 917.650 2300.760 931.270 ;
        RECT 2300.560 917.330 2300.820 917.650 ;
        RECT 2300.560 882.310 2300.820 882.630 ;
        RECT 2300.620 845.650 2300.760 882.310 ;
        RECT 2299.700 845.510 2300.760 845.650 ;
        RECT 2299.700 821.285 2299.840 845.510 ;
        RECT 2299.630 820.915 2299.910 821.285 ;
        RECT 2301.010 820.915 2301.290 821.285 ;
        RECT 2301.080 787.430 2301.220 820.915 ;
        RECT 2301.020 787.110 2301.280 787.430 ;
        RECT 2300.100 786.430 2300.360 786.750 ;
        RECT 2300.160 738.210 2300.300 786.430 ;
        RECT 2300.160 738.070 2301.220 738.210 ;
        RECT 2301.080 724.530 2301.220 738.070 ;
        RECT 2299.640 724.210 2299.900 724.530 ;
        RECT 2301.020 724.210 2301.280 724.530 ;
        RECT 2299.700 676.445 2299.840 724.210 ;
        RECT 2299.630 676.075 2299.910 676.445 ;
        RECT 2300.550 676.075 2300.830 676.445 ;
        RECT 2300.620 642.330 2300.760 676.075 ;
        RECT 2300.160 642.190 2300.760 642.330 ;
        RECT 2300.160 641.650 2300.300 642.190 ;
        RECT 2300.160 641.510 2300.760 641.650 ;
        RECT 2300.620 545.770 2300.760 641.510 ;
        RECT 2300.160 545.630 2300.760 545.770 ;
        RECT 2300.160 545.090 2300.300 545.630 ;
        RECT 2300.160 544.950 2300.760 545.090 ;
        RECT 2300.620 531.410 2300.760 544.950 ;
        RECT 2299.640 531.090 2299.900 531.410 ;
        RECT 2300.560 531.090 2300.820 531.410 ;
        RECT 2299.700 483.325 2299.840 531.090 ;
        RECT 2299.630 482.955 2299.910 483.325 ;
        RECT 2300.550 482.955 2300.830 483.325 ;
        RECT 2300.620 400.930 2300.760 482.955 ;
        RECT 2300.160 400.790 2300.760 400.930 ;
        RECT 2300.160 352.650 2300.300 400.790 ;
        RECT 2300.160 352.510 2300.760 352.650 ;
        RECT 2300.620 351.290 2300.760 352.510 ;
        RECT 2299.700 351.150 2300.760 351.290 ;
        RECT 2299.700 337.950 2299.840 351.150 ;
        RECT 2299.640 337.630 2299.900 337.950 ;
        RECT 2301.020 337.630 2301.280 337.950 ;
        RECT 2301.080 290.090 2301.220 337.630 ;
        RECT 2300.620 289.950 2301.220 290.090 ;
        RECT 2300.620 289.670 2300.760 289.950 ;
        RECT 2300.560 289.350 2300.820 289.670 ;
        RECT 2300.100 241.410 2300.360 241.730 ;
        RECT 2300.160 241.050 2300.300 241.410 ;
        RECT 2300.100 240.730 2300.360 241.050 ;
        RECT 2301.020 206.730 2301.280 207.050 ;
        RECT 2301.080 193.110 2301.220 206.730 ;
        RECT 2301.020 192.790 2301.280 193.110 ;
        RECT 2300.560 158.450 2300.820 158.770 ;
        RECT 2300.620 110.150 2300.760 158.450 ;
        RECT 2300.560 109.830 2300.820 110.150 ;
        RECT 2301.940 109.830 2302.200 110.150 ;
        RECT 2302.000 19.030 2302.140 109.830 ;
        RECT 2301.940 18.710 2302.200 19.030 ;
        RECT 2316.200 18.710 2316.460 19.030 ;
        RECT 2316.260 2.400 2316.400 18.710 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
      LAYER via2 ;
        RECT 2300.090 1594.120 2300.370 1594.400 ;
        RECT 2301.010 1594.120 2301.290 1594.400 ;
        RECT 2300.090 1207.200 2300.370 1207.480 ;
        RECT 2300.550 1172.520 2300.830 1172.800 ;
        RECT 2299.170 1103.840 2299.450 1104.120 ;
        RECT 2300.090 1103.840 2300.370 1104.120 ;
        RECT 2299.630 820.960 2299.910 821.240 ;
        RECT 2301.010 820.960 2301.290 821.240 ;
        RECT 2299.630 676.120 2299.910 676.400 ;
        RECT 2300.550 676.120 2300.830 676.400 ;
        RECT 2299.630 483.000 2299.910 483.280 ;
        RECT 2300.550 483.000 2300.830 483.280 ;
      LAYER met3 ;
        RECT 2300.065 1594.410 2300.395 1594.425 ;
        RECT 2300.985 1594.410 2301.315 1594.425 ;
        RECT 2300.065 1594.110 2301.315 1594.410 ;
        RECT 2300.065 1594.095 2300.395 1594.110 ;
        RECT 2300.985 1594.095 2301.315 1594.110 ;
        RECT 2300.065 1207.500 2300.395 1207.505 ;
        RECT 2300.065 1207.490 2300.650 1207.500 ;
        RECT 2300.065 1207.190 2300.850 1207.490 ;
        RECT 2300.065 1207.180 2300.650 1207.190 ;
        RECT 2300.065 1207.175 2300.395 1207.180 ;
        RECT 2300.525 1172.820 2300.855 1172.825 ;
        RECT 2300.270 1172.810 2300.855 1172.820 ;
        RECT 2300.070 1172.510 2300.855 1172.810 ;
        RECT 2300.270 1172.500 2300.855 1172.510 ;
        RECT 2300.525 1172.495 2300.855 1172.500 ;
        RECT 2299.145 1104.130 2299.475 1104.145 ;
        RECT 2300.065 1104.130 2300.395 1104.145 ;
        RECT 2299.145 1103.830 2300.395 1104.130 ;
        RECT 2299.145 1103.815 2299.475 1103.830 ;
        RECT 2300.065 1103.815 2300.395 1103.830 ;
        RECT 2299.605 821.250 2299.935 821.265 ;
        RECT 2300.985 821.250 2301.315 821.265 ;
        RECT 2299.605 820.950 2301.315 821.250 ;
        RECT 2299.605 820.935 2299.935 820.950 ;
        RECT 2300.985 820.935 2301.315 820.950 ;
        RECT 2299.605 676.410 2299.935 676.425 ;
        RECT 2300.525 676.410 2300.855 676.425 ;
        RECT 2299.605 676.110 2300.855 676.410 ;
        RECT 2299.605 676.095 2299.935 676.110 ;
        RECT 2300.525 676.095 2300.855 676.110 ;
        RECT 2299.605 483.290 2299.935 483.305 ;
        RECT 2300.525 483.290 2300.855 483.305 ;
        RECT 2299.605 482.990 2300.855 483.290 ;
        RECT 2299.605 482.975 2299.935 482.990 ;
        RECT 2300.525 482.975 2300.855 482.990 ;
      LAYER via3 ;
        RECT 2300.300 1207.180 2300.620 1207.500 ;
        RECT 2300.300 1172.500 2300.620 1172.820 ;
      LAYER met4 ;
        RECT 2300.295 1207.175 2300.625 1207.505 ;
        RECT 2300.310 1172.825 2300.610 1207.175 ;
        RECT 2300.295 1172.495 2300.625 1172.825 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2110.090 1689.700 2110.410 1689.760 ;
        RECT 2190.590 1689.700 2190.910 1689.760 ;
        RECT 2110.090 1689.560 2190.910 1689.700 ;
        RECT 2110.090 1689.500 2110.410 1689.560 ;
        RECT 2190.590 1689.500 2190.910 1689.560 ;
        RECT 2190.590 14.180 2190.910 14.240 ;
        RECT 2334.110 14.180 2334.430 14.240 ;
        RECT 2190.590 14.040 2334.430 14.180 ;
        RECT 2190.590 13.980 2190.910 14.040 ;
        RECT 2334.110 13.980 2334.430 14.040 ;
      LAYER via ;
        RECT 2110.120 1689.500 2110.380 1689.760 ;
        RECT 2190.620 1689.500 2190.880 1689.760 ;
        RECT 2190.620 13.980 2190.880 14.240 ;
        RECT 2334.140 13.980 2334.400 14.240 ;
      LAYER met2 ;
        RECT 2110.045 1700.000 2110.325 1704.000 ;
        RECT 2110.180 1689.790 2110.320 1700.000 ;
        RECT 2110.120 1689.470 2110.380 1689.790 ;
        RECT 2190.620 1689.470 2190.880 1689.790 ;
        RECT 2190.680 14.270 2190.820 1689.470 ;
        RECT 2190.620 13.950 2190.880 14.270 ;
        RECT 2334.140 13.950 2334.400 14.270 ;
        RECT 2334.200 2.400 2334.340 13.950 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2307.965 1684.105 2308.135 1686.315 ;
      LAYER mcon ;
        RECT 2307.965 1686.145 2308.135 1686.315 ;
      LAYER met1 ;
        RECT 2117.450 1686.300 2117.770 1686.360 ;
        RECT 2307.905 1686.300 2308.195 1686.345 ;
        RECT 2117.450 1686.160 2308.195 1686.300 ;
        RECT 2117.450 1686.100 2117.770 1686.160 ;
        RECT 2307.905 1686.115 2308.195 1686.160 ;
        RECT 2307.905 1684.260 2308.195 1684.305 ;
        RECT 2346.070 1684.260 2346.390 1684.320 ;
        RECT 2307.905 1684.120 2346.390 1684.260 ;
        RECT 2307.905 1684.075 2308.195 1684.120 ;
        RECT 2346.070 1684.060 2346.390 1684.120 ;
        RECT 2346.070 2.960 2346.390 3.020 ;
        RECT 2351.590 2.960 2351.910 3.020 ;
        RECT 2346.070 2.820 2351.910 2.960 ;
        RECT 2346.070 2.760 2346.390 2.820 ;
        RECT 2351.590 2.760 2351.910 2.820 ;
      LAYER via ;
        RECT 2117.480 1686.100 2117.740 1686.360 ;
        RECT 2346.100 1684.060 2346.360 1684.320 ;
        RECT 2346.100 2.760 2346.360 3.020 ;
        RECT 2351.620 2.760 2351.880 3.020 ;
      LAYER met2 ;
        RECT 2117.405 1700.000 2117.685 1704.000 ;
        RECT 2117.540 1686.390 2117.680 1700.000 ;
        RECT 2117.480 1686.070 2117.740 1686.390 ;
        RECT 2346.100 1684.030 2346.360 1684.350 ;
        RECT 2346.160 3.050 2346.300 1684.030 ;
        RECT 2346.100 2.730 2346.360 3.050 ;
        RECT 2351.620 2.730 2351.880 3.050 ;
        RECT 2351.680 2.400 2351.820 2.730 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2245.405 14.365 2245.575 19.975 ;
      LAYER mcon ;
        RECT 2245.405 19.805 2245.575 19.975 ;
      LAYER met1 ;
        RECT 2124.810 1689.020 2125.130 1689.080 ;
        RECT 2211.290 1689.020 2211.610 1689.080 ;
        RECT 2124.810 1688.880 2211.610 1689.020 ;
        RECT 2124.810 1688.820 2125.130 1688.880 ;
        RECT 2211.290 1688.820 2211.610 1688.880 ;
        RECT 2211.290 20.300 2211.610 20.360 ;
        RECT 2211.290 20.160 2233.600 20.300 ;
        RECT 2211.290 20.100 2211.610 20.160 ;
        RECT 2233.460 19.960 2233.600 20.160 ;
        RECT 2245.345 19.960 2245.635 20.005 ;
        RECT 2233.460 19.820 2245.635 19.960 ;
        RECT 2245.345 19.775 2245.635 19.820 ;
        RECT 2245.345 14.520 2245.635 14.565 ;
        RECT 2369.530 14.520 2369.850 14.580 ;
        RECT 2245.345 14.380 2369.850 14.520 ;
        RECT 2245.345 14.335 2245.635 14.380 ;
        RECT 2369.530 14.320 2369.850 14.380 ;
      LAYER via ;
        RECT 2124.840 1688.820 2125.100 1689.080 ;
        RECT 2211.320 1688.820 2211.580 1689.080 ;
        RECT 2211.320 20.100 2211.580 20.360 ;
        RECT 2369.560 14.320 2369.820 14.580 ;
      LAYER met2 ;
        RECT 2124.765 1700.000 2125.045 1704.000 ;
        RECT 2124.900 1689.110 2125.040 1700.000 ;
        RECT 2124.840 1688.790 2125.100 1689.110 ;
        RECT 2211.320 1688.790 2211.580 1689.110 ;
        RECT 2211.380 20.390 2211.520 1688.790 ;
        RECT 2211.320 20.070 2211.580 20.390 ;
        RECT 2369.560 14.290 2369.820 14.610 ;
        RECT 2369.620 2.400 2369.760 14.290 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2222.405 1684.785 2223.035 1684.955 ;
      LAYER mcon ;
        RECT 2222.865 1684.785 2223.035 1684.955 ;
      LAYER met1 ;
        RECT 2134.010 1684.940 2134.330 1685.000 ;
        RECT 2222.345 1684.940 2222.635 1684.985 ;
        RECT 2134.010 1684.800 2222.635 1684.940 ;
        RECT 2134.010 1684.740 2134.330 1684.800 ;
        RECT 2222.345 1684.755 2222.635 1684.800 ;
        RECT 2222.805 1684.940 2223.095 1684.985 ;
        RECT 2376.890 1684.940 2377.210 1685.000 ;
        RECT 2222.805 1684.800 2377.210 1684.940 ;
        RECT 2222.805 1684.755 2223.095 1684.800 ;
        RECT 2376.890 1684.740 2377.210 1684.800 ;
        RECT 2376.890 15.200 2377.210 15.260 ;
        RECT 2387.470 15.200 2387.790 15.260 ;
        RECT 2376.890 15.060 2387.790 15.200 ;
        RECT 2376.890 15.000 2377.210 15.060 ;
        RECT 2387.470 15.000 2387.790 15.060 ;
      LAYER via ;
        RECT 2134.040 1684.740 2134.300 1685.000 ;
        RECT 2376.920 1684.740 2377.180 1685.000 ;
        RECT 2376.920 15.000 2377.180 15.260 ;
        RECT 2387.500 15.000 2387.760 15.260 ;
      LAYER met2 ;
        RECT 2132.125 1700.410 2132.405 1704.000 ;
        RECT 2132.125 1700.270 2134.240 1700.410 ;
        RECT 2132.125 1700.000 2132.405 1700.270 ;
        RECT 2134.100 1685.030 2134.240 1700.270 ;
        RECT 2134.040 1684.710 2134.300 1685.030 ;
        RECT 2376.920 1684.710 2377.180 1685.030 ;
        RECT 2376.980 15.290 2377.120 1684.710 ;
        RECT 2376.920 14.970 2377.180 15.290 ;
        RECT 2387.500 14.970 2387.760 15.290 ;
        RECT 2387.560 2.400 2387.700 14.970 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 2209.985 1688.185 2210.155 1689.715 ;
        RECT 2307.965 14.705 2308.135 18.275 ;
      LAYER mcon ;
        RECT 2209.985 1689.545 2210.155 1689.715 ;
        RECT 2307.965 18.105 2308.135 18.275 ;
      LAYER met1 ;
        RECT 2209.925 1689.700 2210.215 1689.745 ;
        RECT 2245.790 1689.700 2246.110 1689.760 ;
        RECT 2209.925 1689.560 2246.110 1689.700 ;
        RECT 2209.925 1689.515 2210.215 1689.560 ;
        RECT 2245.790 1689.500 2246.110 1689.560 ;
        RECT 2139.530 1688.340 2139.850 1688.400 ;
        RECT 2209.925 1688.340 2210.215 1688.385 ;
        RECT 2139.530 1688.200 2210.215 1688.340 ;
        RECT 2139.530 1688.140 2139.850 1688.200 ;
        RECT 2209.925 1688.155 2210.215 1688.200 ;
        RECT 2245.790 18.260 2246.110 18.320 ;
        RECT 2307.905 18.260 2308.195 18.305 ;
        RECT 2245.790 18.120 2308.195 18.260 ;
        RECT 2245.790 18.060 2246.110 18.120 ;
        RECT 2307.905 18.075 2308.195 18.120 ;
        RECT 2307.905 14.860 2308.195 14.905 ;
        RECT 2405.410 14.860 2405.730 14.920 ;
        RECT 2307.905 14.720 2405.730 14.860 ;
        RECT 2307.905 14.675 2308.195 14.720 ;
        RECT 2405.410 14.660 2405.730 14.720 ;
      LAYER via ;
        RECT 2245.820 1689.500 2246.080 1689.760 ;
        RECT 2139.560 1688.140 2139.820 1688.400 ;
        RECT 2245.820 18.060 2246.080 18.320 ;
        RECT 2405.440 14.660 2405.700 14.920 ;
      LAYER met2 ;
        RECT 2139.485 1700.000 2139.765 1704.000 ;
        RECT 2139.620 1688.430 2139.760 1700.000 ;
        RECT 2245.820 1689.470 2246.080 1689.790 ;
        RECT 2139.560 1688.110 2139.820 1688.430 ;
        RECT 2245.880 18.350 2246.020 1689.470 ;
        RECT 2245.820 18.030 2246.080 18.350 ;
        RECT 2405.440 14.630 2405.700 14.950 ;
        RECT 2405.500 2.400 2405.640 14.630 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 799.550 35.260 799.870 35.320 ;
        RECT 1476.670 35.260 1476.990 35.320 ;
        RECT 799.550 35.120 1476.990 35.260 ;
        RECT 799.550 35.060 799.870 35.120 ;
        RECT 1476.670 35.060 1476.990 35.120 ;
      LAYER via ;
        RECT 799.580 35.060 799.840 35.320 ;
        RECT 1476.700 35.060 1476.960 35.320 ;
      LAYER met2 ;
        RECT 1478.005 1700.410 1478.285 1704.000 ;
        RECT 1476.760 1700.270 1478.285 1700.410 ;
        RECT 1476.760 35.350 1476.900 1700.270 ;
        RECT 1478.005 1700.000 1478.285 1700.270 ;
        RECT 799.580 35.030 799.840 35.350 ;
        RECT 1476.700 35.030 1476.960 35.350 ;
        RECT 799.640 2.400 799.780 35.030 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1414.525 1700.410 1414.805 1704.000 ;
        RECT 1414.525 1700.270 1415.720 1700.410 ;
        RECT 1414.525 1700.000 1414.805 1700.270 ;
        RECT 1415.580 37.925 1415.720 1700.270 ;
        RECT 645.010 37.555 645.290 37.925 ;
        RECT 1415.510 37.555 1415.790 37.925 ;
        RECT 645.080 2.400 645.220 37.555 ;
        RECT 644.870 -4.800 645.430 2.400 ;
      LAYER via2 ;
        RECT 645.010 37.600 645.290 37.880 ;
        RECT 1415.510 37.600 1415.790 37.880 ;
      LAYER met3 ;
        RECT 644.985 37.890 645.315 37.905 ;
        RECT 1415.485 37.890 1415.815 37.905 ;
        RECT 644.985 37.590 1415.815 37.890 ;
        RECT 644.985 37.575 645.315 37.590 ;
        RECT 1415.485 37.575 1415.815 37.590 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2175.945 1685.465 2176.115 1688.015 ;
        RECT 2222.405 1685.465 2223.495 1685.635 ;
      LAYER mcon ;
        RECT 2175.945 1687.845 2176.115 1688.015 ;
        RECT 2223.325 1685.465 2223.495 1685.635 ;
      LAYER met1 ;
        RECT 2150.570 1688.000 2150.890 1688.060 ;
        RECT 2175.885 1688.000 2176.175 1688.045 ;
        RECT 2150.570 1687.860 2176.175 1688.000 ;
        RECT 2150.570 1687.800 2150.890 1687.860 ;
        RECT 2175.885 1687.815 2176.175 1687.860 ;
        RECT 2175.885 1685.620 2176.175 1685.665 ;
        RECT 2222.345 1685.620 2222.635 1685.665 ;
        RECT 2175.885 1685.480 2222.635 1685.620 ;
        RECT 2175.885 1685.435 2176.175 1685.480 ;
        RECT 2222.345 1685.435 2222.635 1685.480 ;
        RECT 2223.265 1685.620 2223.555 1685.665 ;
        RECT 2428.870 1685.620 2429.190 1685.680 ;
        RECT 2223.265 1685.480 2429.190 1685.620 ;
        RECT 2223.265 1685.435 2223.555 1685.480 ;
        RECT 2428.870 1685.420 2429.190 1685.480 ;
      LAYER via ;
        RECT 2150.600 1687.800 2150.860 1688.060 ;
        RECT 2428.900 1685.420 2429.160 1685.680 ;
      LAYER met2 ;
        RECT 2149.145 1700.410 2149.425 1704.000 ;
        RECT 2149.145 1700.270 2150.800 1700.410 ;
        RECT 2149.145 1700.000 2149.425 1700.270 ;
        RECT 2150.660 1688.090 2150.800 1700.270 ;
        RECT 2150.600 1687.770 2150.860 1688.090 ;
        RECT 2428.900 1685.390 2429.160 1685.710 ;
        RECT 2428.960 2.400 2429.100 1685.390 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2156.550 1684.260 2156.870 1684.320 ;
        RECT 2169.890 1684.260 2170.210 1684.320 ;
        RECT 2156.550 1684.120 2170.210 1684.260 ;
        RECT 2156.550 1684.060 2156.870 1684.120 ;
        RECT 2169.890 1684.060 2170.210 1684.120 ;
        RECT 2169.890 16.220 2170.210 16.280 ;
        RECT 2169.890 16.080 2173.800 16.220 ;
        RECT 2169.890 16.020 2170.210 16.080 ;
        RECT 2173.660 15.880 2173.800 16.080 ;
        RECT 2446.810 15.880 2447.130 15.940 ;
        RECT 2173.660 15.740 2447.130 15.880 ;
        RECT 2446.810 15.680 2447.130 15.740 ;
      LAYER via ;
        RECT 2156.580 1684.060 2156.840 1684.320 ;
        RECT 2169.920 1684.060 2170.180 1684.320 ;
        RECT 2169.920 16.020 2170.180 16.280 ;
        RECT 2446.840 15.680 2447.100 15.940 ;
      LAYER met2 ;
        RECT 2156.505 1700.000 2156.785 1704.000 ;
        RECT 2156.640 1684.350 2156.780 1700.000 ;
        RECT 2156.580 1684.030 2156.840 1684.350 ;
        RECT 2169.920 1684.030 2170.180 1684.350 ;
        RECT 2169.980 16.310 2170.120 1684.030 ;
        RECT 2169.920 15.990 2170.180 16.310 ;
        RECT 2446.840 15.650 2447.100 15.970 ;
        RECT 2446.900 2.400 2447.040 15.650 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2221.945 1685.805 2223.035 1685.975 ;
      LAYER mcon ;
        RECT 2222.865 1685.805 2223.035 1685.975 ;
      LAYER met1 ;
        RECT 2221.885 1685.960 2222.175 1686.005 ;
        RECT 2175.500 1685.820 2222.175 1685.960 ;
        RECT 2163.910 1685.620 2164.230 1685.680 ;
        RECT 2175.500 1685.620 2175.640 1685.820 ;
        RECT 2221.885 1685.775 2222.175 1685.820 ;
        RECT 2222.805 1685.960 2223.095 1686.005 ;
        RECT 2463.370 1685.960 2463.690 1686.020 ;
        RECT 2222.805 1685.820 2463.690 1685.960 ;
        RECT 2222.805 1685.775 2223.095 1685.820 ;
        RECT 2463.370 1685.760 2463.690 1685.820 ;
        RECT 2163.910 1685.480 2175.640 1685.620 ;
        RECT 2163.910 1685.420 2164.230 1685.480 ;
      LAYER via ;
        RECT 2163.940 1685.420 2164.200 1685.680 ;
        RECT 2463.400 1685.760 2463.660 1686.020 ;
      LAYER met2 ;
        RECT 2163.865 1700.000 2164.145 1704.000 ;
        RECT 2164.000 1685.710 2164.140 1700.000 ;
        RECT 2463.400 1685.730 2463.660 1686.050 ;
        RECT 2163.940 1685.390 2164.200 1685.710 ;
        RECT 2463.460 17.410 2463.600 1685.730 ;
        RECT 2463.460 17.270 2464.980 17.410 ;
        RECT 2464.840 2.400 2464.980 17.270 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2171.270 1687.320 2171.590 1687.380 ;
        RECT 2197.490 1687.320 2197.810 1687.380 ;
        RECT 2171.270 1687.180 2197.810 1687.320 ;
        RECT 2171.270 1687.120 2171.590 1687.180 ;
        RECT 2197.490 1687.120 2197.810 1687.180 ;
        RECT 2197.490 16.220 2197.810 16.280 ;
        RECT 2482.690 16.220 2483.010 16.280 ;
        RECT 2197.490 16.080 2483.010 16.220 ;
        RECT 2197.490 16.020 2197.810 16.080 ;
        RECT 2482.690 16.020 2483.010 16.080 ;
      LAYER via ;
        RECT 2171.300 1687.120 2171.560 1687.380 ;
        RECT 2197.520 1687.120 2197.780 1687.380 ;
        RECT 2197.520 16.020 2197.780 16.280 ;
        RECT 2482.720 16.020 2482.980 16.280 ;
      LAYER met2 ;
        RECT 2171.225 1700.000 2171.505 1704.000 ;
        RECT 2171.360 1687.410 2171.500 1700.000 ;
        RECT 2171.300 1687.090 2171.560 1687.410 ;
        RECT 2197.520 1687.090 2197.780 1687.410 ;
        RECT 2197.580 16.310 2197.720 1687.090 ;
        RECT 2197.520 15.990 2197.780 16.310 ;
        RECT 2482.720 15.990 2482.980 16.310 ;
        RECT 2482.780 2.400 2482.920 15.990 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2178.630 1690.380 2178.950 1690.440 ;
        RECT 2497.870 1690.380 2498.190 1690.440 ;
        RECT 2178.630 1690.240 2498.190 1690.380 ;
        RECT 2178.630 1690.180 2178.950 1690.240 ;
        RECT 2497.870 1690.180 2498.190 1690.240 ;
      LAYER via ;
        RECT 2178.660 1690.180 2178.920 1690.440 ;
        RECT 2497.900 1690.180 2498.160 1690.440 ;
      LAYER met2 ;
        RECT 2178.585 1700.000 2178.865 1704.000 ;
        RECT 2178.720 1690.470 2178.860 1700.000 ;
        RECT 2178.660 1690.150 2178.920 1690.470 ;
        RECT 2497.900 1690.150 2498.160 1690.470 ;
        RECT 2497.960 17.410 2498.100 1690.150 ;
        RECT 2497.960 17.270 2500.860 17.410 ;
        RECT 2500.720 2.400 2500.860 17.270 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2185.990 1687.660 2186.310 1687.720 ;
        RECT 2211.750 1687.660 2212.070 1687.720 ;
        RECT 2185.990 1687.520 2212.070 1687.660 ;
        RECT 2185.990 1687.460 2186.310 1687.520 ;
        RECT 2211.750 1687.460 2212.070 1687.520 ;
        RECT 2211.750 16.560 2212.070 16.620 ;
        RECT 2518.110 16.560 2518.430 16.620 ;
        RECT 2211.750 16.420 2518.430 16.560 ;
        RECT 2211.750 16.360 2212.070 16.420 ;
        RECT 2518.110 16.360 2518.430 16.420 ;
      LAYER via ;
        RECT 2186.020 1687.460 2186.280 1687.720 ;
        RECT 2211.780 1687.460 2212.040 1687.720 ;
        RECT 2211.780 16.360 2212.040 16.620 ;
        RECT 2518.140 16.360 2518.400 16.620 ;
      LAYER met2 ;
        RECT 2185.945 1700.000 2186.225 1704.000 ;
        RECT 2186.080 1687.750 2186.220 1700.000 ;
        RECT 2186.020 1687.430 2186.280 1687.750 ;
        RECT 2211.780 1687.430 2212.040 1687.750 ;
        RECT 2211.840 16.650 2211.980 1687.430 ;
        RECT 2211.780 16.330 2212.040 16.650 ;
        RECT 2518.140 16.330 2518.400 16.650 ;
        RECT 2518.200 2.400 2518.340 16.330 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2201.245 1688.525 2201.415 1689.715 ;
      LAYER mcon ;
        RECT 2201.245 1689.545 2201.415 1689.715 ;
      LAYER met1 ;
        RECT 2193.350 1689.700 2193.670 1689.760 ;
        RECT 2201.185 1689.700 2201.475 1689.745 ;
        RECT 2193.350 1689.560 2201.475 1689.700 ;
        RECT 2193.350 1689.500 2193.670 1689.560 ;
        RECT 2201.185 1689.515 2201.475 1689.560 ;
        RECT 2201.185 1688.680 2201.475 1688.725 ;
        RECT 2532.370 1688.680 2532.690 1688.740 ;
        RECT 2201.185 1688.540 2532.690 1688.680 ;
        RECT 2201.185 1688.495 2201.475 1688.540 ;
        RECT 2532.370 1688.480 2532.690 1688.540 ;
      LAYER via ;
        RECT 2193.380 1689.500 2193.640 1689.760 ;
        RECT 2532.400 1688.480 2532.660 1688.740 ;
      LAYER met2 ;
        RECT 2193.305 1700.000 2193.585 1704.000 ;
        RECT 2193.440 1689.790 2193.580 1700.000 ;
        RECT 2193.380 1689.470 2193.640 1689.790 ;
        RECT 2532.400 1688.450 2532.660 1688.770 ;
        RECT 2532.460 17.410 2532.600 1688.450 ;
        RECT 2532.460 17.270 2536.280 17.410 ;
        RECT 2536.140 2.400 2536.280 17.270 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2200.785 1684.105 2200.955 1690.055 ;
        RECT 2234.825 1684.105 2234.995 1686.995 ;
      LAYER mcon ;
        RECT 2200.785 1689.885 2200.955 1690.055 ;
        RECT 2234.825 1686.825 2234.995 1686.995 ;
      LAYER met1 ;
        RECT 2200.710 1690.040 2201.030 1690.100 ;
        RECT 2200.515 1689.900 2201.030 1690.040 ;
        RECT 2200.710 1689.840 2201.030 1689.900 ;
        RECT 2234.765 1686.980 2235.055 1687.025 ;
        RECT 2553.070 1686.980 2553.390 1687.040 ;
        RECT 2234.765 1686.840 2553.390 1686.980 ;
        RECT 2234.765 1686.795 2235.055 1686.840 ;
        RECT 2553.070 1686.780 2553.390 1686.840 ;
        RECT 2200.725 1684.260 2201.015 1684.305 ;
        RECT 2234.765 1684.260 2235.055 1684.305 ;
        RECT 2200.725 1684.120 2235.055 1684.260 ;
        RECT 2200.725 1684.075 2201.015 1684.120 ;
        RECT 2234.765 1684.075 2235.055 1684.120 ;
      LAYER via ;
        RECT 2200.740 1689.840 2201.000 1690.100 ;
        RECT 2553.100 1686.780 2553.360 1687.040 ;
      LAYER met2 ;
        RECT 2200.665 1700.000 2200.945 1704.000 ;
        RECT 2200.800 1690.130 2200.940 1700.000 ;
        RECT 2200.740 1689.810 2201.000 1690.130 ;
        RECT 2553.100 1686.750 2553.360 1687.070 ;
        RECT 2553.160 17.410 2553.300 1686.750 ;
        RECT 2553.160 17.270 2554.220 17.410 ;
        RECT 2554.080 2.400 2554.220 17.270 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2208.070 1688.000 2208.390 1688.060 ;
        RECT 2218.190 1688.000 2218.510 1688.060 ;
        RECT 2208.070 1687.860 2218.510 1688.000 ;
        RECT 2208.070 1687.800 2208.390 1687.860 ;
        RECT 2218.190 1687.800 2218.510 1687.860 ;
        RECT 2218.190 16.900 2218.510 16.960 ;
        RECT 2218.190 16.760 2550.540 16.900 ;
        RECT 2218.190 16.700 2218.510 16.760 ;
        RECT 2550.400 16.560 2550.540 16.760 ;
        RECT 2571.930 16.560 2572.250 16.620 ;
        RECT 2550.400 16.420 2572.250 16.560 ;
        RECT 2571.930 16.360 2572.250 16.420 ;
      LAYER via ;
        RECT 2208.100 1687.800 2208.360 1688.060 ;
        RECT 2218.220 1687.800 2218.480 1688.060 ;
        RECT 2218.220 16.700 2218.480 16.960 ;
        RECT 2571.960 16.360 2572.220 16.620 ;
      LAYER met2 ;
        RECT 2208.025 1700.000 2208.305 1704.000 ;
        RECT 2208.160 1688.090 2208.300 1700.000 ;
        RECT 2208.100 1687.770 2208.360 1688.090 ;
        RECT 2218.220 1687.770 2218.480 1688.090 ;
        RECT 2218.280 16.990 2218.420 1687.770 ;
        RECT 2218.220 16.670 2218.480 16.990 ;
        RECT 2571.960 16.330 2572.220 16.650 ;
        RECT 2572.020 2.400 2572.160 16.330 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2242.645 1687.505 2243.735 1687.675 ;
        RECT 2242.645 1687.165 2242.815 1687.505 ;
      LAYER mcon ;
        RECT 2243.565 1687.505 2243.735 1687.675 ;
      LAYER met1 ;
        RECT 2243.505 1687.660 2243.795 1687.705 ;
        RECT 2570.090 1687.660 2570.410 1687.720 ;
        RECT 2243.505 1687.520 2570.410 1687.660 ;
        RECT 2243.505 1687.475 2243.795 1687.520 ;
        RECT 2570.090 1687.460 2570.410 1687.520 ;
        RECT 2215.430 1687.320 2215.750 1687.380 ;
        RECT 2242.585 1687.320 2242.875 1687.365 ;
        RECT 2215.430 1687.180 2242.875 1687.320 ;
        RECT 2215.430 1687.120 2215.750 1687.180 ;
        RECT 2242.585 1687.135 2242.875 1687.180 ;
        RECT 2570.090 16.900 2570.410 16.960 ;
        RECT 2589.410 16.900 2589.730 16.960 ;
        RECT 2570.090 16.760 2589.730 16.900 ;
        RECT 2570.090 16.700 2570.410 16.760 ;
        RECT 2589.410 16.700 2589.730 16.760 ;
      LAYER via ;
        RECT 2570.120 1687.460 2570.380 1687.720 ;
        RECT 2215.460 1687.120 2215.720 1687.380 ;
        RECT 2570.120 16.700 2570.380 16.960 ;
        RECT 2589.440 16.700 2589.700 16.960 ;
      LAYER met2 ;
        RECT 2215.385 1700.000 2215.665 1704.000 ;
        RECT 2215.520 1687.410 2215.660 1700.000 ;
        RECT 2570.120 1687.430 2570.380 1687.750 ;
        RECT 2215.460 1687.090 2215.720 1687.410 ;
        RECT 2570.180 16.990 2570.320 1687.430 ;
        RECT 2570.120 16.670 2570.380 16.990 ;
        RECT 2589.440 16.670 2589.700 16.990 ;
        RECT 2589.500 2.400 2589.640 16.670 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1485.025 1331.865 1485.195 1379.975 ;
        RECT 1484.105 1247.205 1484.275 1289.875 ;
        RECT 1484.565 613.445 1484.735 696.915 ;
      LAYER mcon ;
        RECT 1485.025 1379.805 1485.195 1379.975 ;
        RECT 1484.105 1289.705 1484.275 1289.875 ;
        RECT 1484.565 696.745 1484.735 696.915 ;
      LAYER met1 ;
        RECT 1484.030 1642.100 1484.350 1642.160 ;
        RECT 1484.950 1642.100 1485.270 1642.160 ;
        RECT 1484.030 1641.960 1485.270 1642.100 ;
        RECT 1484.030 1641.900 1484.350 1641.960 ;
        RECT 1484.950 1641.900 1485.270 1641.960 ;
        RECT 1484.490 1587.020 1484.810 1587.080 ;
        RECT 1484.950 1587.020 1485.270 1587.080 ;
        RECT 1484.490 1586.880 1485.270 1587.020 ;
        RECT 1484.490 1586.820 1484.810 1586.880 ;
        RECT 1484.950 1586.820 1485.270 1586.880 ;
        RECT 1484.030 1505.760 1484.350 1505.820 ;
        RECT 1484.950 1505.760 1485.270 1505.820 ;
        RECT 1484.030 1505.620 1485.270 1505.760 ;
        RECT 1484.030 1505.560 1484.350 1505.620 ;
        RECT 1484.950 1505.560 1485.270 1505.620 ;
        RECT 1484.030 1387.100 1484.350 1387.160 ;
        RECT 1484.490 1387.100 1484.810 1387.160 ;
        RECT 1484.030 1386.960 1484.810 1387.100 ;
        RECT 1484.030 1386.900 1484.350 1386.960 ;
        RECT 1484.490 1386.900 1484.810 1386.960 ;
        RECT 1484.965 1379.960 1485.255 1380.005 ;
        RECT 1485.410 1379.960 1485.730 1380.020 ;
        RECT 1484.965 1379.820 1485.730 1379.960 ;
        RECT 1484.965 1379.775 1485.255 1379.820 ;
        RECT 1485.410 1379.760 1485.730 1379.820 ;
        RECT 1484.950 1332.020 1485.270 1332.080 ;
        RECT 1484.755 1331.880 1485.270 1332.020 ;
        RECT 1484.950 1331.820 1485.270 1331.880 ;
        RECT 1484.030 1314.680 1484.350 1314.740 ;
        RECT 1484.950 1314.680 1485.270 1314.740 ;
        RECT 1484.030 1314.540 1485.270 1314.680 ;
        RECT 1484.030 1314.480 1484.350 1314.540 ;
        RECT 1484.950 1314.480 1485.270 1314.540 ;
        RECT 1484.045 1289.860 1484.335 1289.905 ;
        RECT 1484.950 1289.860 1485.270 1289.920 ;
        RECT 1484.045 1289.720 1485.270 1289.860 ;
        RECT 1484.045 1289.675 1484.335 1289.720 ;
        RECT 1484.950 1289.660 1485.270 1289.720 ;
        RECT 1484.030 1247.360 1484.350 1247.420 ;
        RECT 1483.835 1247.220 1484.350 1247.360 ;
        RECT 1484.030 1247.160 1484.350 1247.220 ;
        RECT 1484.030 1111.020 1484.350 1111.080 ;
        RECT 1484.490 1111.020 1484.810 1111.080 ;
        RECT 1484.030 1110.880 1484.810 1111.020 ;
        RECT 1484.030 1110.820 1484.350 1110.880 ;
        RECT 1484.490 1110.820 1484.810 1110.880 ;
        RECT 1484.030 1014.460 1484.350 1014.520 ;
        RECT 1484.490 1014.460 1484.810 1014.520 ;
        RECT 1484.030 1014.320 1484.810 1014.460 ;
        RECT 1484.030 1014.260 1484.350 1014.320 ;
        RECT 1484.490 1014.260 1484.810 1014.320 ;
        RECT 1484.490 932.180 1484.810 932.240 ;
        RECT 1484.120 932.040 1484.810 932.180 ;
        RECT 1484.120 931.560 1484.260 932.040 ;
        RECT 1484.490 931.980 1484.810 932.040 ;
        RECT 1484.030 931.300 1484.350 931.560 ;
        RECT 1484.030 893.760 1484.350 893.820 ;
        RECT 1484.950 893.760 1485.270 893.820 ;
        RECT 1484.030 893.620 1485.270 893.760 ;
        RECT 1484.030 893.560 1484.350 893.620 ;
        RECT 1484.950 893.560 1485.270 893.620 ;
        RECT 1484.490 807.400 1484.810 807.460 ;
        RECT 1484.950 807.400 1485.270 807.460 ;
        RECT 1484.490 807.260 1485.270 807.400 ;
        RECT 1484.490 807.200 1484.810 807.260 ;
        RECT 1484.950 807.200 1485.270 807.260 ;
        RECT 1483.110 751.980 1483.430 752.040 ;
        RECT 1484.490 751.980 1484.810 752.040 ;
        RECT 1483.110 751.840 1484.810 751.980 ;
        RECT 1483.110 751.780 1483.430 751.840 ;
        RECT 1484.490 751.780 1484.810 751.840 ;
        RECT 1484.030 703.700 1484.350 703.760 ;
        RECT 1484.950 703.700 1485.270 703.760 ;
        RECT 1484.030 703.560 1485.270 703.700 ;
        RECT 1484.030 703.500 1484.350 703.560 ;
        RECT 1484.950 703.500 1485.270 703.560 ;
        RECT 1484.505 696.900 1484.795 696.945 ;
        RECT 1484.950 696.900 1485.270 696.960 ;
        RECT 1484.505 696.760 1485.270 696.900 ;
        RECT 1484.505 696.715 1484.795 696.760 ;
        RECT 1484.950 696.700 1485.270 696.760 ;
        RECT 1484.505 613.600 1484.795 613.645 ;
        RECT 1484.950 613.600 1485.270 613.660 ;
        RECT 1484.505 613.460 1485.270 613.600 ;
        RECT 1484.505 613.415 1484.795 613.460 ;
        RECT 1484.950 613.400 1485.270 613.460 ;
        RECT 1484.950 564.100 1485.270 564.360 ;
        RECT 1485.040 563.680 1485.180 564.100 ;
        RECT 1484.950 563.420 1485.270 563.680 ;
        RECT 1484.490 517.720 1484.810 517.780 ;
        RECT 1484.950 517.720 1485.270 517.780 ;
        RECT 1484.490 517.580 1485.270 517.720 ;
        RECT 1484.490 517.520 1484.810 517.580 ;
        RECT 1484.950 517.520 1485.270 517.580 ;
        RECT 1484.490 475.900 1484.810 475.960 ;
        RECT 1484.950 475.900 1485.270 475.960 ;
        RECT 1484.490 475.760 1485.270 475.900 ;
        RECT 1484.490 475.700 1484.810 475.760 ;
        RECT 1484.950 475.700 1485.270 475.760 ;
        RECT 1484.950 386.820 1485.270 386.880 ;
        RECT 1484.120 386.680 1485.270 386.820 ;
        RECT 1484.120 386.200 1484.260 386.680 ;
        RECT 1484.950 386.620 1485.270 386.680 ;
        RECT 1484.030 385.940 1484.350 386.200 ;
        RECT 827.610 66.880 827.930 66.940 ;
        RECT 1484.490 66.880 1484.810 66.940 ;
        RECT 827.610 66.740 1484.810 66.880 ;
        RECT 827.610 66.680 827.930 66.740 ;
        RECT 1484.490 66.680 1484.810 66.740 ;
        RECT 823.470 2.960 823.790 3.020 ;
        RECT 827.610 2.960 827.930 3.020 ;
        RECT 823.470 2.820 827.930 2.960 ;
        RECT 823.470 2.760 823.790 2.820 ;
        RECT 827.610 2.760 827.930 2.820 ;
      LAYER via ;
        RECT 1484.060 1641.900 1484.320 1642.160 ;
        RECT 1484.980 1641.900 1485.240 1642.160 ;
        RECT 1484.520 1586.820 1484.780 1587.080 ;
        RECT 1484.980 1586.820 1485.240 1587.080 ;
        RECT 1484.060 1505.560 1484.320 1505.820 ;
        RECT 1484.980 1505.560 1485.240 1505.820 ;
        RECT 1484.060 1386.900 1484.320 1387.160 ;
        RECT 1484.520 1386.900 1484.780 1387.160 ;
        RECT 1485.440 1379.760 1485.700 1380.020 ;
        RECT 1484.980 1331.820 1485.240 1332.080 ;
        RECT 1484.060 1314.480 1484.320 1314.740 ;
        RECT 1484.980 1314.480 1485.240 1314.740 ;
        RECT 1484.980 1289.660 1485.240 1289.920 ;
        RECT 1484.060 1247.160 1484.320 1247.420 ;
        RECT 1484.060 1110.820 1484.320 1111.080 ;
        RECT 1484.520 1110.820 1484.780 1111.080 ;
        RECT 1484.060 1014.260 1484.320 1014.520 ;
        RECT 1484.520 1014.260 1484.780 1014.520 ;
        RECT 1484.520 931.980 1484.780 932.240 ;
        RECT 1484.060 931.300 1484.320 931.560 ;
        RECT 1484.060 893.560 1484.320 893.820 ;
        RECT 1484.980 893.560 1485.240 893.820 ;
        RECT 1484.520 807.200 1484.780 807.460 ;
        RECT 1484.980 807.200 1485.240 807.460 ;
        RECT 1483.140 751.780 1483.400 752.040 ;
        RECT 1484.520 751.780 1484.780 752.040 ;
        RECT 1484.060 703.500 1484.320 703.760 ;
        RECT 1484.980 703.500 1485.240 703.760 ;
        RECT 1484.980 696.700 1485.240 696.960 ;
        RECT 1484.980 613.400 1485.240 613.660 ;
        RECT 1484.980 564.100 1485.240 564.360 ;
        RECT 1484.980 563.420 1485.240 563.680 ;
        RECT 1484.520 517.520 1484.780 517.780 ;
        RECT 1484.980 517.520 1485.240 517.780 ;
        RECT 1484.520 475.700 1484.780 475.960 ;
        RECT 1484.980 475.700 1485.240 475.960 ;
        RECT 1484.980 386.620 1485.240 386.880 ;
        RECT 1484.060 385.940 1484.320 386.200 ;
        RECT 827.640 66.680 827.900 66.940 ;
        RECT 1484.520 66.680 1484.780 66.940 ;
        RECT 823.500 2.760 823.760 3.020 ;
        RECT 827.640 2.760 827.900 3.020 ;
      LAYER met2 ;
        RECT 1487.665 1700.410 1487.945 1704.000 ;
        RECT 1486.420 1700.270 1487.945 1700.410 ;
        RECT 1486.420 1660.970 1486.560 1700.270 ;
        RECT 1487.665 1700.000 1487.945 1700.270 ;
        RECT 1484.120 1660.830 1486.560 1660.970 ;
        RECT 1484.120 1642.190 1484.260 1660.830 ;
        RECT 1484.060 1641.870 1484.320 1642.190 ;
        RECT 1484.980 1641.870 1485.240 1642.190 ;
        RECT 1485.040 1617.450 1485.180 1641.870 ;
        RECT 1484.580 1617.310 1485.180 1617.450 ;
        RECT 1484.580 1587.110 1484.720 1617.310 ;
        RECT 1484.520 1586.790 1484.780 1587.110 ;
        RECT 1484.980 1586.790 1485.240 1587.110 ;
        RECT 1485.040 1505.850 1485.180 1586.790 ;
        RECT 1484.060 1505.530 1484.320 1505.850 ;
        RECT 1484.980 1505.530 1485.240 1505.850 ;
        RECT 1484.120 1448.130 1484.260 1505.530 ;
        RECT 1484.120 1447.990 1485.180 1448.130 ;
        RECT 1485.040 1435.210 1485.180 1447.990 ;
        RECT 1484.580 1435.070 1485.180 1435.210 ;
        RECT 1484.580 1387.190 1484.720 1435.070 ;
        RECT 1484.060 1387.045 1484.320 1387.190 ;
        RECT 1484.050 1386.675 1484.330 1387.045 ;
        RECT 1484.520 1386.870 1484.780 1387.190 ;
        RECT 1485.430 1386.675 1485.710 1387.045 ;
        RECT 1485.500 1380.050 1485.640 1386.675 ;
        RECT 1485.440 1379.730 1485.700 1380.050 ;
        RECT 1484.980 1331.790 1485.240 1332.110 ;
        RECT 1485.040 1314.770 1485.180 1331.790 ;
        RECT 1484.060 1314.450 1484.320 1314.770 ;
        RECT 1484.980 1314.450 1485.240 1314.770 ;
        RECT 1484.120 1290.485 1484.260 1314.450 ;
        RECT 1484.050 1290.115 1484.330 1290.485 ;
        RECT 1484.970 1290.115 1485.250 1290.485 ;
        RECT 1485.040 1289.950 1485.180 1290.115 ;
        RECT 1484.980 1289.630 1485.240 1289.950 ;
        RECT 1484.060 1247.130 1484.320 1247.450 ;
        RECT 1484.120 1207.410 1484.260 1247.130 ;
        RECT 1484.120 1207.270 1484.720 1207.410 ;
        RECT 1484.120 1111.110 1484.260 1111.265 ;
        RECT 1484.580 1111.110 1484.720 1207.270 ;
        RECT 1484.060 1110.850 1484.320 1111.110 ;
        RECT 1484.520 1110.850 1484.780 1111.110 ;
        RECT 1484.060 1110.790 1484.780 1110.850 ;
        RECT 1484.120 1110.710 1484.720 1110.790 ;
        RECT 1484.120 1014.550 1484.260 1014.705 ;
        RECT 1484.580 1014.550 1484.720 1110.710 ;
        RECT 1484.060 1014.290 1484.320 1014.550 ;
        RECT 1484.520 1014.290 1484.780 1014.550 ;
        RECT 1484.060 1014.230 1484.780 1014.290 ;
        RECT 1484.120 1014.150 1484.720 1014.230 ;
        RECT 1484.580 932.270 1484.720 1014.150 ;
        RECT 1484.520 931.950 1484.780 932.270 ;
        RECT 1484.060 931.270 1484.320 931.590 ;
        RECT 1484.120 893.850 1484.260 931.270 ;
        RECT 1484.060 893.530 1484.320 893.850 ;
        RECT 1484.980 893.530 1485.240 893.850 ;
        RECT 1485.040 807.490 1485.180 893.530 ;
        RECT 1484.520 807.170 1484.780 807.490 ;
        RECT 1484.980 807.170 1485.240 807.490 ;
        RECT 1484.580 752.070 1484.720 807.170 ;
        RECT 1483.140 751.750 1483.400 752.070 ;
        RECT 1484.520 751.750 1484.780 752.070 ;
        RECT 1483.200 704.325 1483.340 751.750 ;
        RECT 1483.130 703.955 1483.410 704.325 ;
        RECT 1484.050 703.955 1484.330 704.325 ;
        RECT 1484.120 703.790 1484.260 703.955 ;
        RECT 1484.060 703.470 1484.320 703.790 ;
        RECT 1484.980 703.470 1485.240 703.790 ;
        RECT 1485.040 696.990 1485.180 703.470 ;
        RECT 1484.980 696.670 1485.240 696.990 ;
        RECT 1484.980 613.370 1485.240 613.690 ;
        RECT 1485.040 564.390 1485.180 613.370 ;
        RECT 1484.980 564.070 1485.240 564.390 ;
        RECT 1484.980 563.390 1485.240 563.710 ;
        RECT 1485.040 517.810 1485.180 563.390 ;
        RECT 1484.520 517.490 1484.780 517.810 ;
        RECT 1484.980 517.490 1485.240 517.810 ;
        RECT 1484.580 475.990 1484.720 517.490 ;
        RECT 1484.520 475.670 1484.780 475.990 ;
        RECT 1484.980 475.670 1485.240 475.990 ;
        RECT 1485.040 386.910 1485.180 475.670 ;
        RECT 1484.980 386.590 1485.240 386.910 ;
        RECT 1484.060 385.910 1484.320 386.230 ;
        RECT 1484.120 234.330 1484.260 385.910 ;
        RECT 1484.120 234.190 1484.720 234.330 ;
        RECT 1484.580 66.970 1484.720 234.190 ;
        RECT 827.640 66.650 827.900 66.970 ;
        RECT 1484.520 66.650 1484.780 66.970 ;
        RECT 827.700 3.050 827.840 66.650 ;
        RECT 823.500 2.730 823.760 3.050 ;
        RECT 827.640 2.730 827.900 3.050 ;
        RECT 823.560 2.400 823.700 2.730 ;
        RECT 823.350 -4.800 823.910 2.400 ;
      LAYER via2 ;
        RECT 1484.050 1386.720 1484.330 1387.000 ;
        RECT 1485.430 1386.720 1485.710 1387.000 ;
        RECT 1484.050 1290.160 1484.330 1290.440 ;
        RECT 1484.970 1290.160 1485.250 1290.440 ;
        RECT 1483.130 704.000 1483.410 704.280 ;
        RECT 1484.050 704.000 1484.330 704.280 ;
      LAYER met3 ;
        RECT 1484.025 1387.010 1484.355 1387.025 ;
        RECT 1485.405 1387.010 1485.735 1387.025 ;
        RECT 1484.025 1386.710 1485.735 1387.010 ;
        RECT 1484.025 1386.695 1484.355 1386.710 ;
        RECT 1485.405 1386.695 1485.735 1386.710 ;
        RECT 1484.025 1290.450 1484.355 1290.465 ;
        RECT 1484.945 1290.450 1485.275 1290.465 ;
        RECT 1484.025 1290.150 1485.275 1290.450 ;
        RECT 1484.025 1290.135 1484.355 1290.150 ;
        RECT 1484.945 1290.135 1485.275 1290.150 ;
        RECT 1483.105 704.290 1483.435 704.305 ;
        RECT 1484.025 704.290 1484.355 704.305 ;
        RECT 1483.105 703.990 1484.355 704.290 ;
        RECT 1483.105 703.975 1483.435 703.990 ;
        RECT 1484.025 703.975 1484.355 703.990 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2222.790 1689.020 2223.110 1689.080 ;
        RECT 2228.310 1689.020 2228.630 1689.080 ;
        RECT 2222.790 1688.880 2228.630 1689.020 ;
        RECT 2222.790 1688.820 2223.110 1688.880 ;
        RECT 2228.310 1688.820 2228.630 1688.880 ;
        RECT 2228.310 20.640 2228.630 20.700 ;
        RECT 2607.350 20.640 2607.670 20.700 ;
        RECT 2228.310 20.500 2607.670 20.640 ;
        RECT 2228.310 20.440 2228.630 20.500 ;
        RECT 2607.350 20.440 2607.670 20.500 ;
      LAYER via ;
        RECT 2222.820 1688.820 2223.080 1689.080 ;
        RECT 2228.340 1688.820 2228.600 1689.080 ;
        RECT 2228.340 20.440 2228.600 20.700 ;
        RECT 2607.380 20.440 2607.640 20.700 ;
      LAYER met2 ;
        RECT 2222.745 1700.000 2223.025 1704.000 ;
        RECT 2222.880 1689.110 2223.020 1700.000 ;
        RECT 2222.820 1688.790 2223.080 1689.110 ;
        RECT 2228.340 1688.790 2228.600 1689.110 ;
        RECT 2228.400 20.730 2228.540 1688.790 ;
        RECT 2228.340 20.410 2228.600 20.730 ;
        RECT 2607.380 20.410 2607.640 20.730 ;
        RECT 2607.440 2.400 2607.580 20.410 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2266.105 1687.165 2266.275 1689.035 ;
      LAYER mcon ;
        RECT 2266.105 1688.865 2266.275 1689.035 ;
      LAYER met1 ;
        RECT 2230.150 1689.020 2230.470 1689.080 ;
        RECT 2266.045 1689.020 2266.335 1689.065 ;
        RECT 2230.150 1688.880 2266.335 1689.020 ;
        RECT 2230.150 1688.820 2230.470 1688.880 ;
        RECT 2266.045 1688.835 2266.335 1688.880 ;
        RECT 2266.045 1687.320 2266.335 1687.365 ;
        RECT 2583.890 1687.320 2584.210 1687.380 ;
        RECT 2266.045 1687.180 2584.210 1687.320 ;
        RECT 2266.045 1687.135 2266.335 1687.180 ;
        RECT 2583.890 1687.120 2584.210 1687.180 ;
        RECT 2583.430 34.580 2583.750 34.640 ;
        RECT 2584.350 34.580 2584.670 34.640 ;
        RECT 2583.430 34.440 2584.670 34.580 ;
        RECT 2583.430 34.380 2583.750 34.440 ;
        RECT 2584.350 34.380 2584.670 34.440 ;
        RECT 2625.290 16.900 2625.610 16.960 ;
        RECT 2589.960 16.760 2625.610 16.900 ;
        RECT 2584.350 16.560 2584.670 16.620 ;
        RECT 2589.960 16.560 2590.100 16.760 ;
        RECT 2625.290 16.700 2625.610 16.760 ;
        RECT 2584.350 16.420 2590.100 16.560 ;
        RECT 2584.350 16.360 2584.670 16.420 ;
      LAYER via ;
        RECT 2230.180 1688.820 2230.440 1689.080 ;
        RECT 2583.920 1687.120 2584.180 1687.380 ;
        RECT 2583.460 34.380 2583.720 34.640 ;
        RECT 2584.380 34.380 2584.640 34.640 ;
        RECT 2584.380 16.360 2584.640 16.620 ;
        RECT 2625.320 16.700 2625.580 16.960 ;
      LAYER met2 ;
        RECT 2230.105 1700.000 2230.385 1704.000 ;
        RECT 2230.240 1689.110 2230.380 1700.000 ;
        RECT 2230.180 1688.790 2230.440 1689.110 ;
        RECT 2583.920 1687.090 2584.180 1687.410 ;
        RECT 2583.980 58.890 2584.120 1687.090 ;
        RECT 2583.520 58.750 2584.120 58.890 ;
        RECT 2583.520 34.670 2583.660 58.750 ;
        RECT 2583.460 34.350 2583.720 34.670 ;
        RECT 2584.380 34.350 2584.640 34.670 ;
        RECT 2584.440 16.650 2584.580 34.350 ;
        RECT 2625.320 16.670 2625.580 16.990 ;
        RECT 2584.380 16.330 2584.640 16.650 ;
        RECT 2625.380 2.400 2625.520 16.670 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2237.510 1687.660 2237.830 1687.720 ;
        RECT 2242.110 1687.660 2242.430 1687.720 ;
        RECT 2237.510 1687.520 2242.430 1687.660 ;
        RECT 2237.510 1687.460 2237.830 1687.520 ;
        RECT 2242.110 1687.460 2242.430 1687.520 ;
        RECT 2242.110 20.300 2242.430 20.360 ;
        RECT 2643.230 20.300 2643.550 20.360 ;
        RECT 2242.110 20.160 2643.550 20.300 ;
        RECT 2242.110 20.100 2242.430 20.160 ;
        RECT 2643.230 20.100 2643.550 20.160 ;
      LAYER via ;
        RECT 2237.540 1687.460 2237.800 1687.720 ;
        RECT 2242.140 1687.460 2242.400 1687.720 ;
        RECT 2242.140 20.100 2242.400 20.360 ;
        RECT 2643.260 20.100 2643.520 20.360 ;
      LAYER met2 ;
        RECT 2237.465 1700.000 2237.745 1704.000 ;
        RECT 2237.600 1687.750 2237.740 1700.000 ;
        RECT 2237.540 1687.430 2237.800 1687.750 ;
        RECT 2242.140 1687.430 2242.400 1687.750 ;
        RECT 2242.200 20.390 2242.340 1687.430 ;
        RECT 2242.140 20.070 2242.400 20.390 ;
        RECT 2643.260 20.070 2643.520 20.390 ;
        RECT 2643.320 2.400 2643.460 20.070 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2244.870 1688.000 2245.190 1688.060 ;
        RECT 2590.790 1688.000 2591.110 1688.060 ;
        RECT 2244.870 1687.860 2591.110 1688.000 ;
        RECT 2244.870 1687.800 2245.190 1687.860 ;
        RECT 2590.790 1687.800 2591.110 1687.860 ;
        RECT 2590.790 14.180 2591.110 14.240 ;
        RECT 2661.170 14.180 2661.490 14.240 ;
        RECT 2590.790 14.040 2661.490 14.180 ;
        RECT 2590.790 13.980 2591.110 14.040 ;
        RECT 2661.170 13.980 2661.490 14.040 ;
      LAYER via ;
        RECT 2244.900 1687.800 2245.160 1688.060 ;
        RECT 2590.820 1687.800 2591.080 1688.060 ;
        RECT 2590.820 13.980 2591.080 14.240 ;
        RECT 2661.200 13.980 2661.460 14.240 ;
      LAYER met2 ;
        RECT 2244.825 1700.000 2245.105 1704.000 ;
        RECT 2244.960 1688.090 2245.100 1700.000 ;
        RECT 2244.900 1687.770 2245.160 1688.090 ;
        RECT 2590.820 1687.770 2591.080 1688.090 ;
        RECT 2590.880 14.270 2591.020 1687.770 ;
        RECT 2590.820 13.950 2591.080 14.270 ;
        RECT 2661.200 13.950 2661.460 14.270 ;
        RECT 2661.260 2.400 2661.400 13.950 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2252.230 1689.700 2252.550 1689.760 ;
        RECT 2255.910 1689.700 2256.230 1689.760 ;
        RECT 2252.230 1689.560 2256.230 1689.700 ;
        RECT 2252.230 1689.500 2252.550 1689.560 ;
        RECT 2255.910 1689.500 2256.230 1689.560 ;
        RECT 2255.910 19.960 2256.230 20.020 ;
        RECT 2678.650 19.960 2678.970 20.020 ;
        RECT 2255.910 19.820 2678.970 19.960 ;
        RECT 2255.910 19.760 2256.230 19.820 ;
        RECT 2678.650 19.760 2678.970 19.820 ;
      LAYER via ;
        RECT 2252.260 1689.500 2252.520 1689.760 ;
        RECT 2255.940 1689.500 2256.200 1689.760 ;
        RECT 2255.940 19.760 2256.200 20.020 ;
        RECT 2678.680 19.760 2678.940 20.020 ;
      LAYER met2 ;
        RECT 2252.185 1700.000 2252.465 1704.000 ;
        RECT 2252.320 1689.790 2252.460 1700.000 ;
        RECT 2252.260 1689.470 2252.520 1689.790 ;
        RECT 2255.940 1689.470 2256.200 1689.790 ;
        RECT 2256.000 20.050 2256.140 1689.470 ;
        RECT 2255.940 19.730 2256.200 20.050 ;
        RECT 2678.680 19.730 2678.940 20.050 ;
        RECT 2678.740 2.400 2678.880 19.730 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2307.965 1688.185 2308.135 1689.715 ;
      LAYER mcon ;
        RECT 2307.965 1689.545 2308.135 1689.715 ;
      LAYER met1 ;
        RECT 2259.130 1689.700 2259.450 1689.760 ;
        RECT 2307.905 1689.700 2308.195 1689.745 ;
        RECT 2259.130 1689.560 2308.195 1689.700 ;
        RECT 2259.130 1689.500 2259.450 1689.560 ;
        RECT 2307.905 1689.515 2308.195 1689.560 ;
        RECT 2307.905 1688.340 2308.195 1688.385 ;
        RECT 2604.590 1688.340 2604.910 1688.400 ;
        RECT 2307.905 1688.200 2604.910 1688.340 ;
        RECT 2307.905 1688.155 2308.195 1688.200 ;
        RECT 2604.590 1688.140 2604.910 1688.200 ;
        RECT 2604.590 14.520 2604.910 14.580 ;
        RECT 2696.590 14.520 2696.910 14.580 ;
        RECT 2604.590 14.380 2696.910 14.520 ;
        RECT 2604.590 14.320 2604.910 14.380 ;
        RECT 2696.590 14.320 2696.910 14.380 ;
      LAYER via ;
        RECT 2259.160 1689.500 2259.420 1689.760 ;
        RECT 2604.620 1688.140 2604.880 1688.400 ;
        RECT 2604.620 14.320 2604.880 14.580 ;
        RECT 2696.620 14.320 2696.880 14.580 ;
      LAYER met2 ;
        RECT 2259.085 1700.000 2259.365 1704.000 ;
        RECT 2259.220 1689.790 2259.360 1700.000 ;
        RECT 2259.160 1689.470 2259.420 1689.790 ;
        RECT 2604.620 1688.110 2604.880 1688.430 ;
        RECT 2604.680 14.610 2604.820 1688.110 ;
        RECT 2604.620 14.290 2604.880 14.610 ;
        RECT 2696.620 14.290 2696.880 14.610 ;
        RECT 2696.680 2.400 2696.820 14.290 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2266.490 1689.020 2266.810 1689.080 ;
        RECT 2269.710 1689.020 2270.030 1689.080 ;
        RECT 2266.490 1688.880 2270.030 1689.020 ;
        RECT 2266.490 1688.820 2266.810 1688.880 ;
        RECT 2269.710 1688.820 2270.030 1688.880 ;
        RECT 2269.710 19.620 2270.030 19.680 ;
        RECT 2714.530 19.620 2714.850 19.680 ;
        RECT 2269.710 19.480 2714.850 19.620 ;
        RECT 2269.710 19.420 2270.030 19.480 ;
        RECT 2714.530 19.420 2714.850 19.480 ;
      LAYER via ;
        RECT 2266.520 1688.820 2266.780 1689.080 ;
        RECT 2269.740 1688.820 2270.000 1689.080 ;
        RECT 2269.740 19.420 2270.000 19.680 ;
        RECT 2714.560 19.420 2714.820 19.680 ;
      LAYER met2 ;
        RECT 2266.445 1700.000 2266.725 1704.000 ;
        RECT 2266.580 1689.110 2266.720 1700.000 ;
        RECT 2266.520 1688.790 2266.780 1689.110 ;
        RECT 2269.740 1688.790 2270.000 1689.110 ;
        RECT 2269.800 19.710 2269.940 1688.790 ;
        RECT 2269.740 19.390 2270.000 19.710 ;
        RECT 2714.560 19.390 2714.820 19.710 ;
        RECT 2714.620 2.400 2714.760 19.390 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2345.685 1688.865 2345.855 1690.055 ;
      LAYER mcon ;
        RECT 2345.685 1689.885 2345.855 1690.055 ;
      LAYER met1 ;
        RECT 2273.850 1690.040 2274.170 1690.100 ;
        RECT 2345.625 1690.040 2345.915 1690.085 ;
        RECT 2273.850 1689.900 2345.915 1690.040 ;
        RECT 2273.850 1689.840 2274.170 1689.900 ;
        RECT 2345.625 1689.855 2345.915 1689.900 ;
        RECT 2345.625 1689.020 2345.915 1689.065 ;
        RECT 2605.050 1689.020 2605.370 1689.080 ;
        RECT 2345.625 1688.880 2605.370 1689.020 ;
        RECT 2345.625 1688.835 2345.915 1688.880 ;
        RECT 2605.050 1688.820 2605.370 1688.880 ;
        RECT 2605.050 14.860 2605.370 14.920 ;
        RECT 2732.470 14.860 2732.790 14.920 ;
        RECT 2605.050 14.720 2732.790 14.860 ;
        RECT 2605.050 14.660 2605.370 14.720 ;
        RECT 2732.470 14.660 2732.790 14.720 ;
      LAYER via ;
        RECT 2273.880 1689.840 2274.140 1690.100 ;
        RECT 2605.080 1688.820 2605.340 1689.080 ;
        RECT 2605.080 14.660 2605.340 14.920 ;
        RECT 2732.500 14.660 2732.760 14.920 ;
      LAYER met2 ;
        RECT 2273.805 1700.000 2274.085 1704.000 ;
        RECT 2273.940 1690.130 2274.080 1700.000 ;
        RECT 2273.880 1689.810 2274.140 1690.130 ;
        RECT 2605.080 1688.790 2605.340 1689.110 ;
        RECT 2605.140 14.950 2605.280 1688.790 ;
        RECT 2605.080 14.630 2605.340 14.950 ;
        RECT 2732.500 14.630 2732.760 14.950 ;
        RECT 2732.560 2.400 2732.700 14.630 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2330.965 19.125 2332.055 19.295 ;
        RECT 2301.065 17.425 2301.235 18.615 ;
        RECT 2330.965 17.425 2331.135 19.125 ;
      LAYER mcon ;
        RECT 2331.885 19.125 2332.055 19.295 ;
        RECT 2301.065 18.445 2301.235 18.615 ;
      LAYER met1 ;
        RECT 2331.825 19.280 2332.115 19.325 ;
        RECT 2750.410 19.280 2750.730 19.340 ;
        RECT 2331.825 19.140 2750.730 19.280 ;
        RECT 2331.825 19.095 2332.115 19.140 ;
        RECT 2750.410 19.080 2750.730 19.140 ;
        RECT 2283.510 18.600 2283.830 18.660 ;
        RECT 2301.005 18.600 2301.295 18.645 ;
        RECT 2283.510 18.460 2301.295 18.600 ;
        RECT 2283.510 18.400 2283.830 18.460 ;
        RECT 2301.005 18.415 2301.295 18.460 ;
        RECT 2301.005 17.580 2301.295 17.625 ;
        RECT 2330.905 17.580 2331.195 17.625 ;
        RECT 2301.005 17.440 2331.195 17.580 ;
        RECT 2301.005 17.395 2301.295 17.440 ;
        RECT 2330.905 17.395 2331.195 17.440 ;
      LAYER via ;
        RECT 2750.440 19.080 2750.700 19.340 ;
        RECT 2283.540 18.400 2283.800 18.660 ;
      LAYER met2 ;
        RECT 2281.165 1700.410 2281.445 1704.000 ;
        RECT 2281.165 1700.270 2283.740 1700.410 ;
        RECT 2281.165 1700.000 2281.445 1700.270 ;
        RECT 2283.600 18.690 2283.740 1700.270 ;
        RECT 2750.440 19.050 2750.700 19.370 ;
        RECT 2283.540 18.370 2283.800 18.690 ;
        RECT 2750.500 2.400 2750.640 19.050 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2307.505 1689.885 2308.595 1690.055 ;
        RECT 2307.505 1688.185 2307.675 1689.885 ;
        RECT 2308.425 1689.545 2308.595 1689.885 ;
        RECT 2317.165 1689.375 2317.335 1689.715 ;
        RECT 2317.165 1689.205 2318.255 1689.375 ;
      LAYER mcon ;
        RECT 2317.165 1689.545 2317.335 1689.715 ;
        RECT 2318.085 1689.205 2318.255 1689.375 ;
      LAYER met1 ;
        RECT 2308.365 1689.700 2308.655 1689.745 ;
        RECT 2317.105 1689.700 2317.395 1689.745 ;
        RECT 2308.365 1689.560 2317.395 1689.700 ;
        RECT 2308.365 1689.515 2308.655 1689.560 ;
        RECT 2317.105 1689.515 2317.395 1689.560 ;
        RECT 2318.025 1689.360 2318.315 1689.405 ;
        RECT 2618.390 1689.360 2618.710 1689.420 ;
        RECT 2318.025 1689.220 2618.710 1689.360 ;
        RECT 2318.025 1689.175 2318.315 1689.220 ;
        RECT 2618.390 1689.160 2618.710 1689.220 ;
        RECT 2290.870 1688.340 2291.190 1688.400 ;
        RECT 2307.445 1688.340 2307.735 1688.385 ;
        RECT 2290.870 1688.200 2307.735 1688.340 ;
        RECT 2290.870 1688.140 2291.190 1688.200 ;
        RECT 2307.445 1688.155 2307.735 1688.200 ;
        RECT 2618.390 15.200 2618.710 15.260 ;
        RECT 2767.890 15.200 2768.210 15.260 ;
        RECT 2618.390 15.060 2768.210 15.200 ;
        RECT 2618.390 15.000 2618.710 15.060 ;
        RECT 2767.890 15.000 2768.210 15.060 ;
      LAYER via ;
        RECT 2618.420 1689.160 2618.680 1689.420 ;
        RECT 2290.900 1688.140 2291.160 1688.400 ;
        RECT 2618.420 15.000 2618.680 15.260 ;
        RECT 2767.920 15.000 2768.180 15.260 ;
      LAYER met2 ;
        RECT 2288.525 1700.410 2288.805 1704.000 ;
        RECT 2288.525 1700.270 2290.640 1700.410 ;
        RECT 2288.525 1700.000 2288.805 1700.270 ;
        RECT 2290.500 1688.850 2290.640 1700.270 ;
        RECT 2618.420 1689.130 2618.680 1689.450 ;
        RECT 2290.500 1688.710 2291.100 1688.850 ;
        RECT 2290.960 1688.430 2291.100 1688.710 ;
        RECT 2290.900 1688.110 2291.160 1688.430 ;
        RECT 2618.480 15.290 2618.620 1689.130 ;
        RECT 2618.420 14.970 2618.680 15.290 ;
        RECT 2767.920 14.970 2768.180 15.290 ;
        RECT 2767.980 2.400 2768.120 14.970 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1491.390 1678.140 1491.710 1678.200 ;
        RECT 1493.230 1678.140 1493.550 1678.200 ;
        RECT 1491.390 1678.000 1493.550 1678.140 ;
        RECT 1491.390 1677.940 1491.710 1678.000 ;
        RECT 1493.230 1677.940 1493.550 1678.000 ;
        RECT 841.410 67.220 841.730 67.280 ;
        RECT 1491.390 67.220 1491.710 67.280 ;
        RECT 841.410 67.080 1491.710 67.220 ;
        RECT 841.410 67.020 841.730 67.080 ;
        RECT 1491.390 67.020 1491.710 67.080 ;
      LAYER via ;
        RECT 1491.420 1677.940 1491.680 1678.200 ;
        RECT 1493.260 1677.940 1493.520 1678.200 ;
        RECT 841.440 67.020 841.700 67.280 ;
        RECT 1491.420 67.020 1491.680 67.280 ;
      LAYER met2 ;
        RECT 1495.025 1700.410 1495.305 1704.000 ;
        RECT 1493.320 1700.270 1495.305 1700.410 ;
        RECT 1493.320 1678.230 1493.460 1700.270 ;
        RECT 1495.025 1700.000 1495.305 1700.270 ;
        RECT 1491.420 1677.910 1491.680 1678.230 ;
        RECT 1493.260 1677.910 1493.520 1678.230 ;
        RECT 1491.480 67.310 1491.620 1677.910 ;
        RECT 841.440 66.990 841.700 67.310 ;
        RECT 1491.420 66.990 1491.680 67.310 ;
        RECT 841.500 3.130 841.640 66.990 ;
        RECT 841.040 2.990 841.640 3.130 ;
        RECT 841.040 2.400 841.180 2.990 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2295.930 1684.600 2296.250 1684.660 ;
        RECT 2301.450 1684.600 2301.770 1684.660 ;
        RECT 2295.930 1684.460 2301.770 1684.600 ;
        RECT 2295.930 1684.400 2296.250 1684.460 ;
        RECT 2301.450 1684.400 2301.770 1684.460 ;
        RECT 2785.830 18.940 2786.150 19.000 ;
        RECT 2316.720 18.800 2786.150 18.940 ;
        RECT 2301.450 18.600 2301.770 18.660 ;
        RECT 2301.450 18.460 2308.580 18.600 ;
        RECT 2301.450 18.400 2301.770 18.460 ;
        RECT 2308.440 18.260 2308.580 18.460 ;
        RECT 2316.720 18.260 2316.860 18.800 ;
        RECT 2785.830 18.740 2786.150 18.800 ;
        RECT 2308.440 18.120 2316.860 18.260 ;
      LAYER via ;
        RECT 2295.960 1684.400 2296.220 1684.660 ;
        RECT 2301.480 1684.400 2301.740 1684.660 ;
        RECT 2301.480 18.400 2301.740 18.660 ;
        RECT 2785.860 18.740 2786.120 19.000 ;
      LAYER met2 ;
        RECT 2295.885 1700.000 2296.165 1704.000 ;
        RECT 2296.020 1684.690 2296.160 1700.000 ;
        RECT 2295.960 1684.370 2296.220 1684.690 ;
        RECT 2301.480 1684.370 2301.740 1684.690 ;
        RECT 2301.540 18.690 2301.680 1684.370 ;
        RECT 2785.860 18.710 2786.120 19.030 ;
        RECT 2301.480 18.370 2301.740 18.690 ;
        RECT 2785.920 2.400 2786.060 18.710 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2625.290 1689.700 2625.610 1689.760 ;
        RECT 2317.640 1689.560 2625.610 1689.700 ;
        RECT 2303.290 1689.360 2303.610 1689.420 ;
        RECT 2317.640 1689.360 2317.780 1689.560 ;
        RECT 2625.290 1689.500 2625.610 1689.560 ;
        RECT 2303.290 1689.220 2317.780 1689.360 ;
        RECT 2303.290 1689.160 2303.610 1689.220 ;
        RECT 2624.830 15.540 2625.150 15.600 ;
        RECT 2803.770 15.540 2804.090 15.600 ;
        RECT 2624.830 15.400 2804.090 15.540 ;
        RECT 2624.830 15.340 2625.150 15.400 ;
        RECT 2803.770 15.340 2804.090 15.400 ;
      LAYER via ;
        RECT 2303.320 1689.160 2303.580 1689.420 ;
        RECT 2625.320 1689.500 2625.580 1689.760 ;
        RECT 2624.860 15.340 2625.120 15.600 ;
        RECT 2803.800 15.340 2804.060 15.600 ;
      LAYER met2 ;
        RECT 2303.245 1700.000 2303.525 1704.000 ;
        RECT 2303.380 1689.450 2303.520 1700.000 ;
        RECT 2625.320 1689.470 2625.580 1689.790 ;
        RECT 2303.320 1689.130 2303.580 1689.450 ;
        RECT 2625.380 34.410 2625.520 1689.470 ;
        RECT 2624.920 34.270 2625.520 34.410 ;
        RECT 2624.920 15.630 2625.060 34.270 ;
        RECT 2624.860 15.310 2625.120 15.630 ;
        RECT 2803.800 15.310 2804.060 15.630 ;
        RECT 2803.860 2.400 2804.000 15.310 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2821.710 18.600 2822.030 18.660 ;
        RECT 2317.180 18.460 2822.030 18.600 ;
        RECT 2311.110 17.920 2311.430 17.980 ;
        RECT 2317.180 17.920 2317.320 18.460 ;
        RECT 2821.710 18.400 2822.030 18.460 ;
        RECT 2311.110 17.780 2317.320 17.920 ;
        RECT 2311.110 17.720 2311.430 17.780 ;
      LAYER via ;
        RECT 2311.140 17.720 2311.400 17.980 ;
        RECT 2821.740 18.400 2822.000 18.660 ;
      LAYER met2 ;
        RECT 2310.605 1700.410 2310.885 1704.000 ;
        RECT 2310.605 1700.270 2311.340 1700.410 ;
        RECT 2310.605 1700.000 2310.885 1700.270 ;
        RECT 2311.200 18.010 2311.340 1700.270 ;
        RECT 2821.740 18.370 2822.000 18.690 ;
        RECT 2311.140 17.690 2311.400 18.010 ;
        RECT 2821.800 2.400 2821.940 18.370 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2346.145 1686.145 2346.315 1690.055 ;
      LAYER mcon ;
        RECT 2346.145 1689.885 2346.315 1690.055 ;
      LAYER met1 ;
        RECT 2346.085 1690.040 2346.375 1690.085 ;
        RECT 2639.090 1690.040 2639.410 1690.100 ;
        RECT 2346.085 1689.900 2639.410 1690.040 ;
        RECT 2346.085 1689.855 2346.375 1689.900 ;
        RECT 2639.090 1689.840 2639.410 1689.900 ;
        RECT 2318.010 1686.300 2318.330 1686.360 ;
        RECT 2346.085 1686.300 2346.375 1686.345 ;
        RECT 2318.010 1686.160 2346.375 1686.300 ;
        RECT 2318.010 1686.100 2318.330 1686.160 ;
        RECT 2346.085 1686.115 2346.375 1686.160 ;
        RECT 2639.090 16.900 2639.410 16.960 ;
        RECT 2839.190 16.900 2839.510 16.960 ;
        RECT 2639.090 16.760 2839.510 16.900 ;
        RECT 2639.090 16.700 2639.410 16.760 ;
        RECT 2839.190 16.700 2839.510 16.760 ;
      LAYER via ;
        RECT 2639.120 1689.840 2639.380 1690.100 ;
        RECT 2318.040 1686.100 2318.300 1686.360 ;
        RECT 2639.120 16.700 2639.380 16.960 ;
        RECT 2839.220 16.700 2839.480 16.960 ;
      LAYER met2 ;
        RECT 2317.965 1700.000 2318.245 1704.000 ;
        RECT 2318.100 1686.390 2318.240 1700.000 ;
        RECT 2639.120 1689.810 2639.380 1690.130 ;
        RECT 2318.040 1686.070 2318.300 1686.390 ;
        RECT 2639.180 16.990 2639.320 1689.810 ;
        RECT 2639.120 16.670 2639.380 16.990 ;
        RECT 2839.220 16.670 2839.480 16.990 ;
        RECT 2839.280 2.400 2839.420 16.670 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2325.370 1684.600 2325.690 1684.660 ;
        RECT 2331.810 1684.600 2332.130 1684.660 ;
        RECT 2325.370 1684.460 2332.130 1684.600 ;
        RECT 2325.370 1684.400 2325.690 1684.460 ;
        RECT 2331.810 1684.400 2332.130 1684.460 ;
        RECT 2331.810 17.920 2332.130 17.980 ;
        RECT 2857.130 17.920 2857.450 17.980 ;
        RECT 2331.810 17.780 2857.450 17.920 ;
        RECT 2331.810 17.720 2332.130 17.780 ;
        RECT 2857.130 17.720 2857.450 17.780 ;
      LAYER via ;
        RECT 2325.400 1684.400 2325.660 1684.660 ;
        RECT 2331.840 1684.400 2332.100 1684.660 ;
        RECT 2331.840 17.720 2332.100 17.980 ;
        RECT 2857.160 17.720 2857.420 17.980 ;
      LAYER met2 ;
        RECT 2325.325 1700.000 2325.605 1704.000 ;
        RECT 2325.460 1684.690 2325.600 1700.000 ;
        RECT 2325.400 1684.370 2325.660 1684.690 ;
        RECT 2331.840 1684.370 2332.100 1684.690 ;
        RECT 2331.900 18.010 2332.040 1684.370 ;
        RECT 2331.840 17.690 2332.100 18.010 ;
        RECT 2857.160 17.690 2857.420 18.010 ;
        RECT 2857.220 2.400 2857.360 17.690 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2353.430 1686.640 2353.750 1686.700 ;
        RECT 2645.990 1686.640 2646.310 1686.700 ;
        RECT 2353.430 1686.500 2646.310 1686.640 ;
        RECT 2353.430 1686.440 2353.750 1686.500 ;
        RECT 2645.990 1686.440 2646.310 1686.500 ;
        RECT 2332.730 1684.600 2333.050 1684.660 ;
        RECT 2352.510 1684.600 2352.830 1684.660 ;
        RECT 2332.730 1684.460 2352.830 1684.600 ;
        RECT 2332.730 1684.400 2333.050 1684.460 ;
        RECT 2352.510 1684.400 2352.830 1684.460 ;
        RECT 2645.990 20.640 2646.310 20.700 ;
        RECT 2875.070 20.640 2875.390 20.700 ;
        RECT 2645.990 20.500 2875.390 20.640 ;
        RECT 2645.990 20.440 2646.310 20.500 ;
        RECT 2875.070 20.440 2875.390 20.500 ;
      LAYER via ;
        RECT 2353.460 1686.440 2353.720 1686.700 ;
        RECT 2646.020 1686.440 2646.280 1686.700 ;
        RECT 2332.760 1684.400 2333.020 1684.660 ;
        RECT 2352.540 1684.400 2352.800 1684.660 ;
        RECT 2646.020 20.440 2646.280 20.700 ;
        RECT 2875.100 20.440 2875.360 20.700 ;
      LAYER met2 ;
        RECT 2332.685 1700.000 2332.965 1704.000 ;
        RECT 2332.820 1684.690 2332.960 1700.000 ;
        RECT 2353.460 1686.410 2353.720 1686.730 ;
        RECT 2646.020 1686.410 2646.280 1686.730 ;
        RECT 2353.520 1686.245 2353.660 1686.410 ;
        RECT 2352.530 1685.875 2352.810 1686.245 ;
        RECT 2353.450 1685.875 2353.730 1686.245 ;
        RECT 2352.600 1684.690 2352.740 1685.875 ;
        RECT 2332.760 1684.370 2333.020 1684.690 ;
        RECT 2352.540 1684.370 2352.800 1684.690 ;
        RECT 2646.080 20.730 2646.220 1686.410 ;
        RECT 2646.020 20.410 2646.280 20.730 ;
        RECT 2875.100 20.410 2875.360 20.730 ;
        RECT 2875.160 2.400 2875.300 20.410 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
      LAYER via2 ;
        RECT 2352.530 1685.920 2352.810 1686.200 ;
        RECT 2353.450 1685.920 2353.730 1686.200 ;
      LAYER met3 ;
        RECT 2352.505 1686.210 2352.835 1686.225 ;
        RECT 2353.425 1686.210 2353.755 1686.225 ;
        RECT 2352.505 1685.910 2353.755 1686.210 ;
        RECT 2352.505 1685.895 2352.835 1685.910 ;
        RECT 2353.425 1685.895 2353.755 1685.910 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2340.090 1689.020 2340.410 1689.080 ;
        RECT 2345.150 1689.020 2345.470 1689.080 ;
        RECT 2340.090 1688.880 2345.470 1689.020 ;
        RECT 2340.090 1688.820 2340.410 1688.880 ;
        RECT 2345.150 1688.820 2345.470 1688.880 ;
        RECT 2345.150 17.240 2345.470 17.300 ;
        RECT 2893.010 17.240 2893.330 17.300 ;
        RECT 2345.150 17.100 2893.330 17.240 ;
        RECT 2345.150 17.040 2345.470 17.100 ;
        RECT 2893.010 17.040 2893.330 17.100 ;
      LAYER via ;
        RECT 2340.120 1688.820 2340.380 1689.080 ;
        RECT 2345.180 1688.820 2345.440 1689.080 ;
        RECT 2345.180 17.040 2345.440 17.300 ;
        RECT 2893.040 17.040 2893.300 17.300 ;
      LAYER met2 ;
        RECT 2340.045 1700.000 2340.325 1704.000 ;
        RECT 2340.180 1689.110 2340.320 1700.000 ;
        RECT 2340.120 1688.790 2340.380 1689.110 ;
        RECT 2345.180 1688.790 2345.440 1689.110 ;
        RECT 2345.240 17.330 2345.380 1688.790 ;
        RECT 2345.180 17.010 2345.440 17.330 ;
        RECT 2893.040 17.010 2893.300 17.330 ;
        RECT 2893.100 2.400 2893.240 17.010 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2347.450 1686.300 2347.770 1686.360 ;
        RECT 2652.890 1686.300 2653.210 1686.360 ;
        RECT 2347.450 1686.160 2653.210 1686.300 ;
        RECT 2347.450 1686.100 2347.770 1686.160 ;
        RECT 2652.890 1686.100 2653.210 1686.160 ;
        RECT 2652.890 20.300 2653.210 20.360 ;
        RECT 2910.950 20.300 2911.270 20.360 ;
        RECT 2652.890 20.160 2911.270 20.300 ;
        RECT 2652.890 20.100 2653.210 20.160 ;
        RECT 2910.950 20.100 2911.270 20.160 ;
      LAYER via ;
        RECT 2347.480 1686.100 2347.740 1686.360 ;
        RECT 2652.920 1686.100 2653.180 1686.360 ;
        RECT 2652.920 20.100 2653.180 20.360 ;
        RECT 2910.980 20.100 2911.240 20.360 ;
      LAYER met2 ;
        RECT 2347.405 1700.000 2347.685 1704.000 ;
        RECT 2347.540 1686.390 2347.680 1700.000 ;
        RECT 2347.480 1686.070 2347.740 1686.390 ;
        RECT 2652.920 1686.070 2653.180 1686.390 ;
        RECT 2652.980 20.390 2653.120 1686.070 ;
        RECT 2652.920 20.070 2653.180 20.390 ;
        RECT 2910.980 20.070 2911.240 20.390 ;
        RECT 2911.040 2.400 2911.180 20.070 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1499.285 855.525 1499.455 883.915 ;
        RECT 1498.825 620.925 1498.995 669.375 ;
        RECT 1498.825 179.605 1498.995 227.715 ;
      LAYER mcon ;
        RECT 1499.285 883.745 1499.455 883.915 ;
        RECT 1498.825 669.205 1498.995 669.375 ;
        RECT 1498.825 227.545 1498.995 227.715 ;
      LAYER met1 ;
        RECT 1498.750 1655.700 1499.070 1655.760 ;
        RECT 1501.510 1655.700 1501.830 1655.760 ;
        RECT 1498.750 1655.560 1501.830 1655.700 ;
        RECT 1498.750 1655.500 1499.070 1655.560 ;
        RECT 1501.510 1655.500 1501.830 1655.560 ;
        RECT 1498.750 1594.160 1499.070 1594.220 ;
        RECT 1499.210 1594.160 1499.530 1594.220 ;
        RECT 1498.750 1594.020 1499.530 1594.160 ;
        RECT 1498.750 1593.960 1499.070 1594.020 ;
        RECT 1499.210 1593.960 1499.530 1594.020 ;
        RECT 1499.210 1559.820 1499.530 1559.880 ;
        RECT 1498.840 1559.680 1499.530 1559.820 ;
        RECT 1498.840 1559.200 1498.980 1559.680 ;
        RECT 1499.210 1559.620 1499.530 1559.680 ;
        RECT 1498.750 1558.940 1499.070 1559.200 ;
        RECT 1498.750 1497.600 1499.070 1497.660 ;
        RECT 1499.210 1497.600 1499.530 1497.660 ;
        RECT 1498.750 1497.460 1499.530 1497.600 ;
        RECT 1498.750 1497.400 1499.070 1497.460 ;
        RECT 1499.210 1497.400 1499.530 1497.460 ;
        RECT 1499.210 1463.060 1499.530 1463.320 ;
        RECT 1499.300 1462.640 1499.440 1463.060 ;
        RECT 1499.210 1462.380 1499.530 1462.640 ;
        RECT 1499.210 1353.100 1499.530 1353.160 ;
        RECT 1498.840 1352.960 1499.530 1353.100 ;
        RECT 1498.840 1352.820 1498.980 1352.960 ;
        RECT 1499.210 1352.900 1499.530 1352.960 ;
        RECT 1498.750 1352.560 1499.070 1352.820 ;
        RECT 1498.750 1249.060 1499.070 1249.120 ;
        RECT 1499.670 1249.060 1499.990 1249.120 ;
        RECT 1498.750 1248.920 1499.990 1249.060 ;
        RECT 1498.750 1248.860 1499.070 1248.920 ;
        RECT 1499.670 1248.860 1499.990 1248.920 ;
        RECT 1498.750 1200.780 1499.070 1200.840 ;
        RECT 1499.670 1200.780 1499.990 1200.840 ;
        RECT 1498.750 1200.640 1499.990 1200.780 ;
        RECT 1498.750 1200.580 1499.070 1200.640 ;
        RECT 1499.670 1200.580 1499.990 1200.640 ;
        RECT 1498.750 1068.520 1499.070 1068.580 ;
        RECT 1499.670 1068.520 1499.990 1068.580 ;
        RECT 1498.750 1068.380 1499.990 1068.520 ;
        RECT 1498.750 1068.320 1499.070 1068.380 ;
        RECT 1499.670 1068.320 1499.990 1068.380 ;
        RECT 1498.750 1014.460 1499.070 1014.520 ;
        RECT 1499.210 1014.460 1499.530 1014.520 ;
        RECT 1498.750 1014.320 1499.530 1014.460 ;
        RECT 1498.750 1014.260 1499.070 1014.320 ;
        RECT 1499.210 1014.260 1499.530 1014.320 ;
        RECT 1499.210 980.460 1499.530 980.520 ;
        RECT 1498.840 980.320 1499.530 980.460 ;
        RECT 1498.840 979.840 1498.980 980.320 ;
        RECT 1499.210 980.260 1499.530 980.320 ;
        RECT 1498.750 979.580 1499.070 979.840 ;
        RECT 1498.750 917.900 1499.070 917.960 ;
        RECT 1499.210 917.900 1499.530 917.960 ;
        RECT 1498.750 917.760 1499.530 917.900 ;
        RECT 1498.750 917.700 1499.070 917.760 ;
        RECT 1499.210 917.700 1499.530 917.760 ;
        RECT 1499.210 883.900 1499.530 883.960 ;
        RECT 1499.015 883.760 1499.530 883.900 ;
        RECT 1499.210 883.700 1499.530 883.760 ;
        RECT 1498.750 855.680 1499.070 855.740 ;
        RECT 1499.225 855.680 1499.515 855.725 ;
        RECT 1498.750 855.540 1499.515 855.680 ;
        RECT 1498.750 855.480 1499.070 855.540 ;
        RECT 1499.225 855.495 1499.515 855.540 ;
        RECT 1498.750 783.260 1499.070 783.320 ;
        RECT 1499.670 783.260 1499.990 783.320 ;
        RECT 1498.750 783.120 1499.990 783.260 ;
        RECT 1498.750 783.060 1499.070 783.120 ;
        RECT 1499.670 783.060 1499.990 783.120 ;
        RECT 1498.750 687.040 1499.070 687.100 ;
        RECT 1499.670 687.040 1499.990 687.100 ;
        RECT 1498.750 686.900 1499.990 687.040 ;
        RECT 1498.750 686.840 1499.070 686.900 ;
        RECT 1499.670 686.840 1499.990 686.900 ;
        RECT 1498.750 669.360 1499.070 669.420 ;
        RECT 1498.555 669.220 1499.070 669.360 ;
        RECT 1498.750 669.160 1499.070 669.220 ;
        RECT 1498.765 621.080 1499.055 621.125 ;
        RECT 1499.210 621.080 1499.530 621.140 ;
        RECT 1498.765 620.940 1499.530 621.080 ;
        RECT 1498.765 620.895 1499.055 620.940 ;
        RECT 1499.210 620.880 1499.530 620.940 ;
        RECT 1498.290 524.520 1498.610 524.580 ;
        RECT 1498.750 524.520 1499.070 524.580 ;
        RECT 1498.290 524.380 1499.070 524.520 ;
        RECT 1498.290 524.320 1498.610 524.380 ;
        RECT 1498.750 524.320 1499.070 524.380 ;
        RECT 1498.750 476.580 1499.070 476.640 ;
        RECT 1498.750 476.440 1499.440 476.580 ;
        RECT 1498.750 476.380 1499.070 476.440 ;
        RECT 1499.300 476.300 1499.440 476.440 ;
        RECT 1499.210 476.040 1499.530 476.300 ;
        RECT 1499.210 386.620 1499.530 386.880 ;
        RECT 1499.300 386.200 1499.440 386.620 ;
        RECT 1499.210 385.940 1499.530 386.200 ;
        RECT 1498.750 338.200 1499.070 338.260 ;
        RECT 1499.210 338.200 1499.530 338.260 ;
        RECT 1498.750 338.060 1499.530 338.200 ;
        RECT 1498.750 338.000 1499.070 338.060 ;
        RECT 1499.210 338.000 1499.530 338.060 ;
        RECT 1498.750 241.440 1499.070 241.700 ;
        RECT 1498.840 240.960 1498.980 241.440 ;
        RECT 1499.210 240.960 1499.530 241.020 ;
        RECT 1498.840 240.820 1499.530 240.960 ;
        RECT 1499.210 240.760 1499.530 240.820 ;
        RECT 1498.765 227.700 1499.055 227.745 ;
        RECT 1499.210 227.700 1499.530 227.760 ;
        RECT 1498.765 227.560 1499.530 227.700 ;
        RECT 1498.765 227.515 1499.055 227.560 ;
        RECT 1499.210 227.500 1499.530 227.560 ;
        RECT 1498.750 179.760 1499.070 179.820 ;
        RECT 1498.555 179.620 1499.070 179.760 ;
        RECT 1498.750 179.560 1499.070 179.620 ;
        RECT 862.110 67.560 862.430 67.620 ;
        RECT 1498.750 67.560 1499.070 67.620 ;
        RECT 862.110 67.420 1499.070 67.560 ;
        RECT 862.110 67.360 862.430 67.420 ;
        RECT 1498.750 67.360 1499.070 67.420 ;
      LAYER via ;
        RECT 1498.780 1655.500 1499.040 1655.760 ;
        RECT 1501.540 1655.500 1501.800 1655.760 ;
        RECT 1498.780 1593.960 1499.040 1594.220 ;
        RECT 1499.240 1593.960 1499.500 1594.220 ;
        RECT 1499.240 1559.620 1499.500 1559.880 ;
        RECT 1498.780 1558.940 1499.040 1559.200 ;
        RECT 1498.780 1497.400 1499.040 1497.660 ;
        RECT 1499.240 1497.400 1499.500 1497.660 ;
        RECT 1499.240 1463.060 1499.500 1463.320 ;
        RECT 1499.240 1462.380 1499.500 1462.640 ;
        RECT 1499.240 1352.900 1499.500 1353.160 ;
        RECT 1498.780 1352.560 1499.040 1352.820 ;
        RECT 1498.780 1248.860 1499.040 1249.120 ;
        RECT 1499.700 1248.860 1499.960 1249.120 ;
        RECT 1498.780 1200.580 1499.040 1200.840 ;
        RECT 1499.700 1200.580 1499.960 1200.840 ;
        RECT 1498.780 1068.320 1499.040 1068.580 ;
        RECT 1499.700 1068.320 1499.960 1068.580 ;
        RECT 1498.780 1014.260 1499.040 1014.520 ;
        RECT 1499.240 1014.260 1499.500 1014.520 ;
        RECT 1499.240 980.260 1499.500 980.520 ;
        RECT 1498.780 979.580 1499.040 979.840 ;
        RECT 1498.780 917.700 1499.040 917.960 ;
        RECT 1499.240 917.700 1499.500 917.960 ;
        RECT 1499.240 883.700 1499.500 883.960 ;
        RECT 1498.780 855.480 1499.040 855.740 ;
        RECT 1498.780 783.060 1499.040 783.320 ;
        RECT 1499.700 783.060 1499.960 783.320 ;
        RECT 1498.780 686.840 1499.040 687.100 ;
        RECT 1499.700 686.840 1499.960 687.100 ;
        RECT 1498.780 669.160 1499.040 669.420 ;
        RECT 1499.240 620.880 1499.500 621.140 ;
        RECT 1498.320 524.320 1498.580 524.580 ;
        RECT 1498.780 524.320 1499.040 524.580 ;
        RECT 1498.780 476.380 1499.040 476.640 ;
        RECT 1499.240 476.040 1499.500 476.300 ;
        RECT 1499.240 386.620 1499.500 386.880 ;
        RECT 1499.240 385.940 1499.500 386.200 ;
        RECT 1498.780 338.000 1499.040 338.260 ;
        RECT 1499.240 338.000 1499.500 338.260 ;
        RECT 1498.780 241.440 1499.040 241.700 ;
        RECT 1499.240 240.760 1499.500 241.020 ;
        RECT 1499.240 227.500 1499.500 227.760 ;
        RECT 1498.780 179.560 1499.040 179.820 ;
        RECT 862.140 67.360 862.400 67.620 ;
        RECT 1498.780 67.360 1499.040 67.620 ;
      LAYER met2 ;
        RECT 1502.385 1700.410 1502.665 1704.000 ;
        RECT 1502.060 1700.270 1502.665 1700.410 ;
        RECT 1502.060 1695.650 1502.200 1700.270 ;
        RECT 1502.385 1700.000 1502.665 1700.270 ;
        RECT 1501.600 1695.510 1502.200 1695.650 ;
        RECT 1501.600 1655.790 1501.740 1695.510 ;
        RECT 1498.780 1655.470 1499.040 1655.790 ;
        RECT 1501.540 1655.470 1501.800 1655.790 ;
        RECT 1498.840 1594.250 1498.980 1655.470 ;
        RECT 1498.780 1593.930 1499.040 1594.250 ;
        RECT 1499.240 1593.930 1499.500 1594.250 ;
        RECT 1499.300 1559.910 1499.440 1593.930 ;
        RECT 1499.240 1559.590 1499.500 1559.910 ;
        RECT 1498.780 1558.910 1499.040 1559.230 ;
        RECT 1498.840 1497.690 1498.980 1558.910 ;
        RECT 1498.780 1497.370 1499.040 1497.690 ;
        RECT 1499.240 1497.370 1499.500 1497.690 ;
        RECT 1499.300 1463.350 1499.440 1497.370 ;
        RECT 1499.240 1463.030 1499.500 1463.350 ;
        RECT 1499.240 1462.350 1499.500 1462.670 ;
        RECT 1499.300 1353.190 1499.440 1462.350 ;
        RECT 1499.240 1352.870 1499.500 1353.190 ;
        RECT 1498.780 1352.530 1499.040 1352.850 ;
        RECT 1498.840 1334.570 1498.980 1352.530 ;
        RECT 1498.840 1334.430 1499.900 1334.570 ;
        RECT 1499.760 1317.570 1499.900 1334.430 ;
        RECT 1499.300 1317.430 1499.900 1317.570 ;
        RECT 1499.300 1273.370 1499.440 1317.430 ;
        RECT 1499.300 1273.230 1499.900 1273.370 ;
        RECT 1499.760 1249.150 1499.900 1273.230 ;
        RECT 1498.780 1248.830 1499.040 1249.150 ;
        RECT 1499.700 1248.830 1499.960 1249.150 ;
        RECT 1498.840 1200.870 1498.980 1248.830 ;
        RECT 1498.780 1200.550 1499.040 1200.870 ;
        RECT 1499.700 1200.550 1499.960 1200.870 ;
        RECT 1499.760 1159.810 1499.900 1200.550 ;
        RECT 1499.760 1159.670 1500.360 1159.810 ;
        RECT 1500.220 1158.450 1500.360 1159.670 ;
        RECT 1499.300 1158.310 1500.360 1158.450 ;
        RECT 1499.300 1104.050 1499.440 1158.310 ;
        RECT 1499.300 1103.910 1499.900 1104.050 ;
        RECT 1499.760 1068.610 1499.900 1103.910 ;
        RECT 1498.780 1068.290 1499.040 1068.610 ;
        RECT 1499.700 1068.290 1499.960 1068.610 ;
        RECT 1498.840 1014.550 1498.980 1068.290 ;
        RECT 1498.780 1014.230 1499.040 1014.550 ;
        RECT 1499.240 1014.230 1499.500 1014.550 ;
        RECT 1499.300 980.550 1499.440 1014.230 ;
        RECT 1499.240 980.230 1499.500 980.550 ;
        RECT 1498.780 979.550 1499.040 979.870 ;
        RECT 1498.840 917.990 1498.980 979.550 ;
        RECT 1498.780 917.670 1499.040 917.990 ;
        RECT 1499.240 917.670 1499.500 917.990 ;
        RECT 1499.300 883.990 1499.440 917.670 ;
        RECT 1499.240 883.670 1499.500 883.990 ;
        RECT 1498.780 855.450 1499.040 855.770 ;
        RECT 1498.840 783.350 1498.980 855.450 ;
        RECT 1498.780 783.030 1499.040 783.350 ;
        RECT 1499.700 783.030 1499.960 783.350 ;
        RECT 1499.760 687.130 1499.900 783.030 ;
        RECT 1498.780 686.810 1499.040 687.130 ;
        RECT 1499.700 686.810 1499.960 687.130 ;
        RECT 1498.840 669.450 1498.980 686.810 ;
        RECT 1498.780 669.130 1499.040 669.450 ;
        RECT 1499.240 620.850 1499.500 621.170 ;
        RECT 1499.300 579.770 1499.440 620.850 ;
        RECT 1498.380 579.630 1499.440 579.770 ;
        RECT 1498.380 524.610 1498.520 579.630 ;
        RECT 1498.320 524.290 1498.580 524.610 ;
        RECT 1498.780 524.290 1499.040 524.610 ;
        RECT 1498.840 476.670 1498.980 524.290 ;
        RECT 1498.780 476.350 1499.040 476.670 ;
        RECT 1499.240 476.010 1499.500 476.330 ;
        RECT 1499.300 386.910 1499.440 476.010 ;
        RECT 1499.240 386.590 1499.500 386.910 ;
        RECT 1499.240 385.910 1499.500 386.230 ;
        RECT 1499.300 338.290 1499.440 385.910 ;
        RECT 1498.780 337.970 1499.040 338.290 ;
        RECT 1499.240 337.970 1499.500 338.290 ;
        RECT 1498.840 241.730 1498.980 337.970 ;
        RECT 1498.780 241.410 1499.040 241.730 ;
        RECT 1499.240 240.730 1499.500 241.050 ;
        RECT 1499.300 227.790 1499.440 240.730 ;
        RECT 1499.240 227.470 1499.500 227.790 ;
        RECT 1498.780 179.530 1499.040 179.850 ;
        RECT 1498.840 145.250 1498.980 179.530 ;
        RECT 1498.380 145.110 1498.980 145.250 ;
        RECT 1498.380 144.570 1498.520 145.110 ;
        RECT 1498.380 144.430 1498.980 144.570 ;
        RECT 1498.840 67.650 1498.980 144.430 ;
        RECT 862.140 67.330 862.400 67.650 ;
        RECT 1498.780 67.330 1499.040 67.650 ;
        RECT 862.200 16.730 862.340 67.330 ;
        RECT 858.980 16.590 862.340 16.730 ;
        RECT 858.980 2.400 859.120 16.590 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1505.265 1587.205 1505.435 1635.315 ;
        RECT 1505.265 1462.425 1505.435 1490.475 ;
        RECT 1505.265 1242.105 1505.435 1249.415 ;
        RECT 1505.265 855.525 1505.435 903.975 ;
        RECT 1505.265 620.925 1505.435 669.375 ;
      LAYER mcon ;
        RECT 1505.265 1635.145 1505.435 1635.315 ;
        RECT 1505.265 1490.305 1505.435 1490.475 ;
        RECT 1505.265 1249.245 1505.435 1249.415 ;
        RECT 1505.265 903.805 1505.435 903.975 ;
        RECT 1505.265 669.205 1505.435 669.375 ;
      LAYER met1 ;
        RECT 1505.650 1642.440 1505.970 1642.500 ;
        RECT 1508.410 1642.440 1508.730 1642.500 ;
        RECT 1505.650 1642.300 1508.730 1642.440 ;
        RECT 1505.650 1642.240 1505.970 1642.300 ;
        RECT 1508.410 1642.240 1508.730 1642.300 ;
        RECT 1505.205 1635.300 1505.495 1635.345 ;
        RECT 1505.650 1635.300 1505.970 1635.360 ;
        RECT 1505.205 1635.160 1505.970 1635.300 ;
        RECT 1505.205 1635.115 1505.495 1635.160 ;
        RECT 1505.650 1635.100 1505.970 1635.160 ;
        RECT 1505.190 1587.360 1505.510 1587.420 ;
        RECT 1504.995 1587.220 1505.510 1587.360 ;
        RECT 1505.190 1587.160 1505.510 1587.220 ;
        RECT 1505.190 1490.460 1505.510 1490.520 ;
        RECT 1504.995 1490.320 1505.510 1490.460 ;
        RECT 1505.190 1490.260 1505.510 1490.320 ;
        RECT 1505.190 1462.580 1505.510 1462.640 ;
        RECT 1504.995 1462.440 1505.510 1462.580 ;
        RECT 1505.190 1462.380 1505.510 1462.440 ;
        RECT 1505.190 1366.160 1505.510 1366.420 ;
        RECT 1505.280 1366.020 1505.420 1366.160 ;
        RECT 1505.650 1366.020 1505.970 1366.080 ;
        RECT 1505.280 1365.880 1505.970 1366.020 ;
        RECT 1505.650 1365.820 1505.970 1365.880 ;
        RECT 1505.205 1249.400 1505.495 1249.445 ;
        RECT 1505.650 1249.400 1505.970 1249.460 ;
        RECT 1505.205 1249.260 1505.970 1249.400 ;
        RECT 1505.205 1249.215 1505.495 1249.260 ;
        RECT 1505.650 1249.200 1505.970 1249.260 ;
        RECT 1505.190 1242.260 1505.510 1242.320 ;
        RECT 1504.995 1242.120 1505.510 1242.260 ;
        RECT 1505.190 1242.060 1505.510 1242.120 ;
        RECT 1505.190 1200.780 1505.510 1200.840 ;
        RECT 1505.650 1200.780 1505.970 1200.840 ;
        RECT 1505.190 1200.640 1505.970 1200.780 ;
        RECT 1505.190 1200.580 1505.510 1200.640 ;
        RECT 1505.650 1200.580 1505.970 1200.640 ;
        RECT 1505.650 1159.100 1505.970 1159.360 ;
        RECT 1505.740 1158.960 1505.880 1159.100 ;
        RECT 1506.110 1158.960 1506.430 1159.020 ;
        RECT 1505.740 1158.820 1506.430 1158.960 ;
        RECT 1506.110 1158.760 1506.430 1158.820 ;
        RECT 1505.190 1111.020 1505.510 1111.080 ;
        RECT 1506.110 1111.020 1506.430 1111.080 ;
        RECT 1505.190 1110.880 1506.430 1111.020 ;
        RECT 1505.190 1110.820 1505.510 1110.880 ;
        RECT 1506.110 1110.820 1506.430 1110.880 ;
        RECT 1505.190 1076.480 1505.510 1076.740 ;
        RECT 1505.280 1076.000 1505.420 1076.480 ;
        RECT 1505.650 1076.000 1505.970 1076.060 ;
        RECT 1505.280 1075.860 1505.970 1076.000 ;
        RECT 1505.650 1075.800 1505.970 1075.860 ;
        RECT 1505.190 1014.460 1505.510 1014.520 ;
        RECT 1505.650 1014.460 1505.970 1014.520 ;
        RECT 1505.190 1014.320 1505.970 1014.460 ;
        RECT 1505.190 1014.260 1505.510 1014.320 ;
        RECT 1505.650 1014.260 1505.970 1014.320 ;
        RECT 1505.190 979.920 1505.510 980.180 ;
        RECT 1505.280 979.440 1505.420 979.920 ;
        RECT 1505.650 979.440 1505.970 979.500 ;
        RECT 1505.280 979.300 1505.970 979.440 ;
        RECT 1505.650 979.240 1505.970 979.300 ;
        RECT 1505.190 917.900 1505.510 917.960 ;
        RECT 1505.650 917.900 1505.970 917.960 ;
        RECT 1505.190 917.760 1505.970 917.900 ;
        RECT 1505.190 917.700 1505.510 917.760 ;
        RECT 1505.650 917.700 1505.970 917.760 ;
        RECT 1505.190 903.960 1505.510 904.020 ;
        RECT 1504.995 903.820 1505.510 903.960 ;
        RECT 1505.190 903.760 1505.510 903.820 ;
        RECT 1505.190 855.680 1505.510 855.740 ;
        RECT 1504.995 855.540 1505.510 855.680 ;
        RECT 1505.190 855.480 1505.510 855.540 ;
        RECT 1505.190 669.360 1505.510 669.420 ;
        RECT 1504.995 669.220 1505.510 669.360 ;
        RECT 1505.190 669.160 1505.510 669.220 ;
        RECT 1505.205 621.080 1505.495 621.125 ;
        RECT 1505.650 621.080 1505.970 621.140 ;
        RECT 1505.205 620.940 1505.970 621.080 ;
        RECT 1505.205 620.895 1505.495 620.940 ;
        RECT 1505.650 620.880 1505.970 620.940 ;
        RECT 1505.650 566.340 1505.970 566.400 ;
        RECT 1505.280 566.200 1505.970 566.340 ;
        RECT 1505.280 566.060 1505.420 566.200 ;
        RECT 1505.650 566.140 1505.970 566.200 ;
        RECT 1505.190 565.800 1505.510 566.060 ;
        RECT 1505.190 338.200 1505.510 338.260 ;
        RECT 1506.110 338.200 1506.430 338.260 ;
        RECT 1505.190 338.060 1506.430 338.200 ;
        RECT 1505.190 338.000 1505.510 338.060 ;
        RECT 1506.110 338.000 1506.430 338.060 ;
        RECT 1505.190 241.440 1505.510 241.700 ;
        RECT 1505.280 240.960 1505.420 241.440 ;
        RECT 1505.650 240.960 1505.970 241.020 ;
        RECT 1505.280 240.820 1505.970 240.960 ;
        RECT 1505.650 240.760 1505.970 240.820 ;
        RECT 1505.650 145.080 1505.970 145.140 ;
        RECT 1506.110 145.080 1506.430 145.140 ;
        RECT 1505.650 144.940 1506.430 145.080 ;
        RECT 1505.650 144.880 1505.970 144.940 ;
        RECT 1506.110 144.880 1506.430 144.940 ;
        RECT 882.810 67.900 883.130 67.960 ;
        RECT 1505.190 67.900 1505.510 67.960 ;
        RECT 882.810 67.760 1505.510 67.900 ;
        RECT 882.810 67.700 883.130 67.760 ;
        RECT 1505.190 67.700 1505.510 67.760 ;
        RECT 876.830 20.980 877.150 21.040 ;
        RECT 882.810 20.980 883.130 21.040 ;
        RECT 876.830 20.840 883.130 20.980 ;
        RECT 876.830 20.780 877.150 20.840 ;
        RECT 882.810 20.780 883.130 20.840 ;
      LAYER via ;
        RECT 1505.680 1642.240 1505.940 1642.500 ;
        RECT 1508.440 1642.240 1508.700 1642.500 ;
        RECT 1505.680 1635.100 1505.940 1635.360 ;
        RECT 1505.220 1587.160 1505.480 1587.420 ;
        RECT 1505.220 1490.260 1505.480 1490.520 ;
        RECT 1505.220 1462.380 1505.480 1462.640 ;
        RECT 1505.220 1366.160 1505.480 1366.420 ;
        RECT 1505.680 1365.820 1505.940 1366.080 ;
        RECT 1505.680 1249.200 1505.940 1249.460 ;
        RECT 1505.220 1242.060 1505.480 1242.320 ;
        RECT 1505.220 1200.580 1505.480 1200.840 ;
        RECT 1505.680 1200.580 1505.940 1200.840 ;
        RECT 1505.680 1159.100 1505.940 1159.360 ;
        RECT 1506.140 1158.760 1506.400 1159.020 ;
        RECT 1505.220 1110.820 1505.480 1111.080 ;
        RECT 1506.140 1110.820 1506.400 1111.080 ;
        RECT 1505.220 1076.480 1505.480 1076.740 ;
        RECT 1505.680 1075.800 1505.940 1076.060 ;
        RECT 1505.220 1014.260 1505.480 1014.520 ;
        RECT 1505.680 1014.260 1505.940 1014.520 ;
        RECT 1505.220 979.920 1505.480 980.180 ;
        RECT 1505.680 979.240 1505.940 979.500 ;
        RECT 1505.220 917.700 1505.480 917.960 ;
        RECT 1505.680 917.700 1505.940 917.960 ;
        RECT 1505.220 903.760 1505.480 904.020 ;
        RECT 1505.220 855.480 1505.480 855.740 ;
        RECT 1505.220 669.160 1505.480 669.420 ;
        RECT 1505.680 620.880 1505.940 621.140 ;
        RECT 1505.680 566.140 1505.940 566.400 ;
        RECT 1505.220 565.800 1505.480 566.060 ;
        RECT 1505.220 338.000 1505.480 338.260 ;
        RECT 1506.140 338.000 1506.400 338.260 ;
        RECT 1505.220 241.440 1505.480 241.700 ;
        RECT 1505.680 240.760 1505.940 241.020 ;
        RECT 1505.680 144.880 1505.940 145.140 ;
        RECT 1506.140 144.880 1506.400 145.140 ;
        RECT 882.840 67.700 883.100 67.960 ;
        RECT 1505.220 67.700 1505.480 67.960 ;
        RECT 876.860 20.780 877.120 21.040 ;
        RECT 882.840 20.780 883.100 21.040 ;
      LAYER met2 ;
        RECT 1509.745 1700.410 1510.025 1704.000 ;
        RECT 1508.500 1700.270 1510.025 1700.410 ;
        RECT 1508.500 1642.530 1508.640 1700.270 ;
        RECT 1509.745 1700.000 1510.025 1700.270 ;
        RECT 1505.680 1642.210 1505.940 1642.530 ;
        RECT 1508.440 1642.210 1508.700 1642.530 ;
        RECT 1505.740 1635.390 1505.880 1642.210 ;
        RECT 1505.680 1635.070 1505.940 1635.390 ;
        RECT 1505.220 1587.130 1505.480 1587.450 ;
        RECT 1505.280 1539.930 1505.420 1587.130 ;
        RECT 1505.280 1539.790 1505.880 1539.930 ;
        RECT 1505.740 1539.250 1505.880 1539.790 ;
        RECT 1505.280 1539.110 1505.880 1539.250 ;
        RECT 1505.280 1490.550 1505.420 1539.110 ;
        RECT 1505.220 1490.230 1505.480 1490.550 ;
        RECT 1505.220 1462.350 1505.480 1462.670 ;
        RECT 1505.280 1366.450 1505.420 1462.350 ;
        RECT 1505.220 1366.130 1505.480 1366.450 ;
        RECT 1505.680 1365.790 1505.940 1366.110 ;
        RECT 1505.740 1345.450 1505.880 1365.790 ;
        RECT 1505.740 1345.310 1506.800 1345.450 ;
        RECT 1506.660 1303.290 1506.800 1345.310 ;
        RECT 1506.200 1303.150 1506.800 1303.290 ;
        RECT 1506.200 1297.170 1506.340 1303.150 ;
        RECT 1505.740 1297.030 1506.340 1297.170 ;
        RECT 1505.740 1249.490 1505.880 1297.030 ;
        RECT 1505.680 1249.170 1505.940 1249.490 ;
        RECT 1505.220 1242.030 1505.480 1242.350 ;
        RECT 1505.280 1200.870 1505.420 1242.030 ;
        RECT 1505.220 1200.550 1505.480 1200.870 ;
        RECT 1505.680 1200.550 1505.940 1200.870 ;
        RECT 1505.740 1159.390 1505.880 1200.550 ;
        RECT 1505.680 1159.070 1505.940 1159.390 ;
        RECT 1506.140 1158.730 1506.400 1159.050 ;
        RECT 1506.200 1111.110 1506.340 1158.730 ;
        RECT 1505.220 1110.790 1505.480 1111.110 ;
        RECT 1506.140 1110.790 1506.400 1111.110 ;
        RECT 1505.280 1076.770 1505.420 1110.790 ;
        RECT 1505.220 1076.450 1505.480 1076.770 ;
        RECT 1505.680 1075.770 1505.940 1076.090 ;
        RECT 1505.740 1014.550 1505.880 1075.770 ;
        RECT 1505.220 1014.230 1505.480 1014.550 ;
        RECT 1505.680 1014.230 1505.940 1014.550 ;
        RECT 1505.280 980.210 1505.420 1014.230 ;
        RECT 1505.220 979.890 1505.480 980.210 ;
        RECT 1505.680 979.210 1505.940 979.530 ;
        RECT 1505.740 917.990 1505.880 979.210 ;
        RECT 1505.220 917.670 1505.480 917.990 ;
        RECT 1505.680 917.670 1505.940 917.990 ;
        RECT 1505.280 904.050 1505.420 917.670 ;
        RECT 1505.220 903.730 1505.480 904.050 ;
        RECT 1505.220 855.450 1505.480 855.770 ;
        RECT 1505.280 772.890 1505.420 855.450 ;
        RECT 1505.280 772.750 1505.880 772.890 ;
        RECT 1505.740 676.330 1505.880 772.750 ;
        RECT 1505.280 676.190 1505.880 676.330 ;
        RECT 1505.280 669.450 1505.420 676.190 ;
        RECT 1505.220 669.130 1505.480 669.450 ;
        RECT 1505.680 620.850 1505.940 621.170 ;
        RECT 1505.740 566.430 1505.880 620.850 ;
        RECT 1505.680 566.110 1505.940 566.430 ;
        RECT 1505.220 565.770 1505.480 566.090 ;
        RECT 1505.280 500.210 1505.420 565.770 ;
        RECT 1505.280 500.070 1506.340 500.210 ;
        RECT 1506.200 338.290 1506.340 500.070 ;
        RECT 1505.220 337.970 1505.480 338.290 ;
        RECT 1506.140 337.970 1506.400 338.290 ;
        RECT 1505.280 241.730 1505.420 337.970 ;
        RECT 1505.220 241.410 1505.480 241.730 ;
        RECT 1505.680 240.730 1505.940 241.050 ;
        RECT 1505.740 227.530 1505.880 240.730 ;
        RECT 1505.740 227.390 1506.340 227.530 ;
        RECT 1506.200 145.170 1506.340 227.390 ;
        RECT 1505.680 144.850 1505.940 145.170 ;
        RECT 1506.140 144.850 1506.400 145.170 ;
        RECT 1505.740 111.250 1505.880 144.850 ;
        RECT 1505.740 111.110 1506.340 111.250 ;
        RECT 1506.200 109.890 1506.340 111.110 ;
        RECT 1505.280 109.750 1506.340 109.890 ;
        RECT 1505.280 67.990 1505.420 109.750 ;
        RECT 882.840 67.670 883.100 67.990 ;
        RECT 1505.220 67.670 1505.480 67.990 ;
        RECT 882.900 21.070 883.040 67.670 ;
        RECT 876.860 20.750 877.120 21.070 ;
        RECT 882.840 20.750 883.100 21.070 ;
        RECT 876.920 2.400 877.060 20.750 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1512.550 1673.720 1512.870 1673.780 ;
        RECT 1515.310 1673.720 1515.630 1673.780 ;
        RECT 1512.550 1673.580 1515.630 1673.720 ;
        RECT 1512.550 1673.520 1512.870 1673.580 ;
        RECT 1515.310 1673.520 1515.630 1673.580 ;
        RECT 1512.550 1594.160 1512.870 1594.220 ;
        RECT 1513.010 1594.160 1513.330 1594.220 ;
        RECT 1512.550 1594.020 1513.330 1594.160 ;
        RECT 1512.550 1593.960 1512.870 1594.020 ;
        RECT 1513.010 1593.960 1513.330 1594.020 ;
        RECT 1513.010 1559.820 1513.330 1559.880 ;
        RECT 1512.640 1559.680 1513.330 1559.820 ;
        RECT 1512.640 1559.200 1512.780 1559.680 ;
        RECT 1513.010 1559.620 1513.330 1559.680 ;
        RECT 1512.550 1558.940 1512.870 1559.200 ;
        RECT 1512.550 1497.600 1512.870 1497.660 ;
        RECT 1513.010 1497.600 1513.330 1497.660 ;
        RECT 1512.550 1497.460 1513.330 1497.600 ;
        RECT 1512.550 1497.400 1512.870 1497.460 ;
        RECT 1513.010 1497.400 1513.330 1497.460 ;
        RECT 1512.550 1352.760 1512.870 1352.820 ;
        RECT 1513.470 1352.760 1513.790 1352.820 ;
        RECT 1512.550 1352.620 1513.790 1352.760 ;
        RECT 1512.550 1352.560 1512.870 1352.620 ;
        RECT 1513.470 1352.560 1513.790 1352.620 ;
        RECT 1512.550 1249.060 1512.870 1249.120 ;
        RECT 1513.010 1249.060 1513.330 1249.120 ;
        RECT 1512.550 1248.920 1513.330 1249.060 ;
        RECT 1512.550 1248.860 1512.870 1248.920 ;
        RECT 1513.010 1248.860 1513.330 1248.920 ;
        RECT 1512.550 1200.780 1512.870 1200.840 ;
        RECT 1513.470 1200.780 1513.790 1200.840 ;
        RECT 1512.550 1200.640 1513.790 1200.780 ;
        RECT 1512.550 1200.580 1512.870 1200.640 ;
        RECT 1513.470 1200.580 1513.790 1200.640 ;
        RECT 1513.470 1159.640 1513.790 1159.700 ;
        RECT 1513.100 1159.500 1513.790 1159.640 ;
        RECT 1513.100 1159.020 1513.240 1159.500 ;
        RECT 1513.470 1159.440 1513.790 1159.500 ;
        RECT 1513.010 1158.760 1513.330 1159.020 ;
        RECT 1512.550 1014.460 1512.870 1014.520 ;
        RECT 1513.010 1014.460 1513.330 1014.520 ;
        RECT 1512.550 1014.320 1513.330 1014.460 ;
        RECT 1512.550 1014.260 1512.870 1014.320 ;
        RECT 1513.010 1014.260 1513.330 1014.320 ;
        RECT 1513.010 980.460 1513.330 980.520 ;
        RECT 1512.640 980.320 1513.330 980.460 ;
        RECT 1512.640 979.840 1512.780 980.320 ;
        RECT 1513.010 980.260 1513.330 980.320 ;
        RECT 1512.550 979.580 1512.870 979.840 ;
        RECT 1512.550 917.900 1512.870 917.960 ;
        RECT 1513.010 917.900 1513.330 917.960 ;
        RECT 1512.550 917.760 1513.330 917.900 ;
        RECT 1512.550 917.700 1512.870 917.760 ;
        RECT 1513.010 917.700 1513.330 917.760 ;
        RECT 1513.010 883.700 1513.330 883.960 ;
        RECT 1513.100 883.280 1513.240 883.700 ;
        RECT 1513.010 883.020 1513.330 883.280 ;
        RECT 1512.550 692.820 1512.870 692.880 ;
        RECT 1513.470 692.820 1513.790 692.880 ;
        RECT 1512.550 692.680 1513.790 692.820 ;
        RECT 1512.550 692.620 1512.870 692.680 ;
        RECT 1513.470 692.620 1513.790 692.680 ;
        RECT 1512.550 386.480 1512.870 386.540 ;
        RECT 1513.010 386.480 1513.330 386.540 ;
        RECT 1512.550 386.340 1513.330 386.480 ;
        RECT 1512.550 386.280 1512.870 386.340 ;
        RECT 1513.010 386.280 1513.330 386.340 ;
        RECT 1512.550 331.060 1512.870 331.120 ;
        RECT 1513.470 331.060 1513.790 331.120 ;
        RECT 1512.550 330.920 1513.790 331.060 ;
        RECT 1512.550 330.860 1512.870 330.920 ;
        RECT 1513.470 330.860 1513.790 330.920 ;
        RECT 1512.550 137.940 1512.870 138.000 ;
        RECT 1513.010 137.940 1513.330 138.000 ;
        RECT 1512.550 137.800 1513.330 137.940 ;
        RECT 1512.550 137.740 1512.870 137.800 ;
        RECT 1513.010 137.740 1513.330 137.800 ;
        RECT 896.610 68.240 896.930 68.300 ;
        RECT 1512.550 68.240 1512.870 68.300 ;
        RECT 896.610 68.100 1512.870 68.240 ;
        RECT 896.610 68.040 896.930 68.100 ;
        RECT 1512.550 68.040 1512.870 68.100 ;
      LAYER via ;
        RECT 1512.580 1673.520 1512.840 1673.780 ;
        RECT 1515.340 1673.520 1515.600 1673.780 ;
        RECT 1512.580 1593.960 1512.840 1594.220 ;
        RECT 1513.040 1593.960 1513.300 1594.220 ;
        RECT 1513.040 1559.620 1513.300 1559.880 ;
        RECT 1512.580 1558.940 1512.840 1559.200 ;
        RECT 1512.580 1497.400 1512.840 1497.660 ;
        RECT 1513.040 1497.400 1513.300 1497.660 ;
        RECT 1512.580 1352.560 1512.840 1352.820 ;
        RECT 1513.500 1352.560 1513.760 1352.820 ;
        RECT 1512.580 1248.860 1512.840 1249.120 ;
        RECT 1513.040 1248.860 1513.300 1249.120 ;
        RECT 1512.580 1200.580 1512.840 1200.840 ;
        RECT 1513.500 1200.580 1513.760 1200.840 ;
        RECT 1513.500 1159.440 1513.760 1159.700 ;
        RECT 1513.040 1158.760 1513.300 1159.020 ;
        RECT 1512.580 1014.260 1512.840 1014.520 ;
        RECT 1513.040 1014.260 1513.300 1014.520 ;
        RECT 1513.040 980.260 1513.300 980.520 ;
        RECT 1512.580 979.580 1512.840 979.840 ;
        RECT 1512.580 917.700 1512.840 917.960 ;
        RECT 1513.040 917.700 1513.300 917.960 ;
        RECT 1513.040 883.700 1513.300 883.960 ;
        RECT 1513.040 883.020 1513.300 883.280 ;
        RECT 1512.580 692.620 1512.840 692.880 ;
        RECT 1513.500 692.620 1513.760 692.880 ;
        RECT 1512.580 386.280 1512.840 386.540 ;
        RECT 1513.040 386.280 1513.300 386.540 ;
        RECT 1512.580 330.860 1512.840 331.120 ;
        RECT 1513.500 330.860 1513.760 331.120 ;
        RECT 1512.580 137.740 1512.840 138.000 ;
        RECT 1513.040 137.740 1513.300 138.000 ;
        RECT 896.640 68.040 896.900 68.300 ;
        RECT 1512.580 68.040 1512.840 68.300 ;
      LAYER met2 ;
        RECT 1517.105 1700.410 1517.385 1704.000 ;
        RECT 1515.400 1700.270 1517.385 1700.410 ;
        RECT 1515.400 1673.810 1515.540 1700.270 ;
        RECT 1517.105 1700.000 1517.385 1700.270 ;
        RECT 1512.580 1673.490 1512.840 1673.810 ;
        RECT 1515.340 1673.490 1515.600 1673.810 ;
        RECT 1512.640 1594.250 1512.780 1673.490 ;
        RECT 1512.580 1593.930 1512.840 1594.250 ;
        RECT 1513.040 1593.930 1513.300 1594.250 ;
        RECT 1513.100 1559.910 1513.240 1593.930 ;
        RECT 1513.040 1559.590 1513.300 1559.910 ;
        RECT 1512.580 1558.910 1512.840 1559.230 ;
        RECT 1512.640 1497.690 1512.780 1558.910 ;
        RECT 1512.580 1497.370 1512.840 1497.690 ;
        RECT 1513.040 1497.370 1513.300 1497.690 ;
        RECT 1513.100 1466.490 1513.240 1497.370 ;
        RECT 1512.640 1466.350 1513.240 1466.490 ;
        RECT 1512.640 1425.010 1512.780 1466.350 ;
        RECT 1512.640 1424.870 1513.700 1425.010 ;
        RECT 1513.560 1352.850 1513.700 1424.870 ;
        RECT 1512.580 1352.530 1512.840 1352.850 ;
        RECT 1513.500 1352.530 1513.760 1352.850 ;
        RECT 1512.640 1321.650 1512.780 1352.530 ;
        RECT 1512.640 1321.510 1513.700 1321.650 ;
        RECT 1513.560 1317.570 1513.700 1321.510 ;
        RECT 1513.100 1317.430 1513.700 1317.570 ;
        RECT 1513.100 1249.150 1513.240 1317.430 ;
        RECT 1512.580 1248.830 1512.840 1249.150 ;
        RECT 1513.040 1248.830 1513.300 1249.150 ;
        RECT 1512.640 1200.870 1512.780 1248.830 ;
        RECT 1512.580 1200.550 1512.840 1200.870 ;
        RECT 1513.500 1200.550 1513.760 1200.870 ;
        RECT 1513.560 1159.730 1513.700 1200.550 ;
        RECT 1513.500 1159.410 1513.760 1159.730 ;
        RECT 1513.040 1158.730 1513.300 1159.050 ;
        RECT 1513.100 1104.165 1513.240 1158.730 ;
        RECT 1513.030 1103.795 1513.310 1104.165 ;
        RECT 1512.570 1103.115 1512.850 1103.485 ;
        RECT 1512.640 1014.550 1512.780 1103.115 ;
        RECT 1512.580 1014.230 1512.840 1014.550 ;
        RECT 1513.040 1014.230 1513.300 1014.550 ;
        RECT 1513.100 980.550 1513.240 1014.230 ;
        RECT 1513.040 980.230 1513.300 980.550 ;
        RECT 1512.580 979.550 1512.840 979.870 ;
        RECT 1512.640 917.990 1512.780 979.550 ;
        RECT 1512.580 917.670 1512.840 917.990 ;
        RECT 1513.040 917.670 1513.300 917.990 ;
        RECT 1513.100 883.990 1513.240 917.670 ;
        RECT 1513.040 883.670 1513.300 883.990 ;
        RECT 1513.040 882.990 1513.300 883.310 ;
        RECT 1513.100 772.890 1513.240 882.990 ;
        RECT 1512.640 772.750 1513.240 772.890 ;
        RECT 1512.640 749.090 1512.780 772.750 ;
        RECT 1512.640 748.950 1513.700 749.090 ;
        RECT 1513.560 692.910 1513.700 748.950 ;
        RECT 1512.580 692.590 1512.840 692.910 ;
        RECT 1513.500 692.590 1513.760 692.910 ;
        RECT 1512.640 641.650 1512.780 692.590 ;
        RECT 1512.640 641.510 1513.240 641.650 ;
        RECT 1513.100 497.490 1513.240 641.510 ;
        RECT 1512.640 497.350 1513.240 497.490 ;
        RECT 1512.640 447.850 1512.780 497.350 ;
        RECT 1512.640 447.710 1513.240 447.850 ;
        RECT 1513.100 386.570 1513.240 447.710 ;
        RECT 1512.580 386.250 1512.840 386.570 ;
        RECT 1513.040 386.250 1513.300 386.570 ;
        RECT 1512.640 331.150 1512.780 386.250 ;
        RECT 1512.580 330.830 1512.840 331.150 ;
        RECT 1513.500 330.830 1513.760 331.150 ;
        RECT 1513.560 193.360 1513.700 330.830 ;
        RECT 1512.640 193.220 1513.700 193.360 ;
        RECT 1512.640 192.850 1512.780 193.220 ;
        RECT 1512.640 192.710 1513.240 192.850 ;
        RECT 1513.100 138.030 1513.240 192.710 ;
        RECT 1512.580 137.710 1512.840 138.030 ;
        RECT 1513.040 137.710 1513.300 138.030 ;
        RECT 1512.640 68.330 1512.780 137.710 ;
        RECT 896.640 68.010 896.900 68.330 ;
        RECT 1512.580 68.010 1512.840 68.330 ;
        RECT 896.700 16.730 896.840 68.010 ;
        RECT 894.860 16.590 896.840 16.730 ;
        RECT 894.860 2.400 895.000 16.590 ;
        RECT 894.650 -4.800 895.210 2.400 ;
      LAYER via2 ;
        RECT 1513.030 1103.840 1513.310 1104.120 ;
        RECT 1512.570 1103.160 1512.850 1103.440 ;
      LAYER met3 ;
        RECT 1513.005 1104.130 1513.335 1104.145 ;
        RECT 1512.790 1103.815 1513.335 1104.130 ;
        RECT 1512.790 1103.465 1513.090 1103.815 ;
        RECT 1512.545 1103.150 1513.090 1103.465 ;
        RECT 1512.545 1103.135 1512.875 1103.150 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1519.525 565.845 1519.695 613.955 ;
        RECT 1519.525 269.025 1519.695 317.475 ;
        RECT 1519.985 124.185 1520.155 131.495 ;
      LAYER mcon ;
        RECT 1519.525 613.785 1519.695 613.955 ;
        RECT 1519.525 317.305 1519.695 317.475 ;
        RECT 1519.985 131.325 1520.155 131.495 ;
      LAYER met1 ;
        RECT 1519.450 1656.040 1519.770 1656.100 ;
        RECT 1523.130 1656.040 1523.450 1656.100 ;
        RECT 1519.450 1655.900 1523.450 1656.040 ;
        RECT 1519.450 1655.840 1519.770 1655.900 ;
        RECT 1523.130 1655.840 1523.450 1655.900 ;
        RECT 1519.450 613.940 1519.770 614.000 ;
        RECT 1519.255 613.800 1519.770 613.940 ;
        RECT 1519.450 613.740 1519.770 613.800 ;
        RECT 1519.450 566.000 1519.770 566.060 ;
        RECT 1519.255 565.860 1519.770 566.000 ;
        RECT 1519.450 565.800 1519.770 565.860 ;
        RECT 1519.450 373.360 1519.770 373.620 ;
        RECT 1519.540 372.940 1519.680 373.360 ;
        RECT 1519.450 372.680 1519.770 372.940 ;
        RECT 1519.450 317.460 1519.770 317.520 ;
        RECT 1519.255 317.320 1519.770 317.460 ;
        RECT 1519.450 317.260 1519.770 317.320 ;
        RECT 1519.465 269.180 1519.755 269.225 ;
        RECT 1519.910 269.180 1520.230 269.240 ;
        RECT 1519.465 269.040 1520.230 269.180 ;
        RECT 1519.465 268.995 1519.755 269.040 ;
        RECT 1519.910 268.980 1520.230 269.040 ;
        RECT 1518.990 212.060 1519.310 212.120 ;
        RECT 1520.370 212.060 1520.690 212.120 ;
        RECT 1518.990 211.920 1520.690 212.060 ;
        RECT 1518.990 211.860 1519.310 211.920 ;
        RECT 1520.370 211.860 1520.690 211.920 ;
        RECT 1519.910 131.480 1520.230 131.540 ;
        RECT 1519.715 131.340 1520.230 131.480 ;
        RECT 1519.910 131.280 1520.230 131.340 ;
        RECT 1519.910 124.340 1520.230 124.400 ;
        RECT 1519.715 124.200 1520.230 124.340 ;
        RECT 1519.910 124.140 1520.230 124.200 ;
        RECT 917.310 68.920 917.630 68.980 ;
        RECT 1519.910 68.920 1520.230 68.980 ;
        RECT 917.310 68.780 1520.230 68.920 ;
        RECT 917.310 68.720 917.630 68.780 ;
        RECT 1519.910 68.720 1520.230 68.780 ;
        RECT 912.710 2.960 913.030 3.020 ;
        RECT 917.310 2.960 917.630 3.020 ;
        RECT 912.710 2.820 917.630 2.960 ;
        RECT 912.710 2.760 913.030 2.820 ;
        RECT 917.310 2.760 917.630 2.820 ;
      LAYER via ;
        RECT 1519.480 1655.840 1519.740 1656.100 ;
        RECT 1523.160 1655.840 1523.420 1656.100 ;
        RECT 1519.480 613.740 1519.740 614.000 ;
        RECT 1519.480 565.800 1519.740 566.060 ;
        RECT 1519.480 373.360 1519.740 373.620 ;
        RECT 1519.480 372.680 1519.740 372.940 ;
        RECT 1519.480 317.260 1519.740 317.520 ;
        RECT 1519.940 268.980 1520.200 269.240 ;
        RECT 1519.020 211.860 1519.280 212.120 ;
        RECT 1520.400 211.860 1520.660 212.120 ;
        RECT 1519.940 131.280 1520.200 131.540 ;
        RECT 1519.940 124.140 1520.200 124.400 ;
        RECT 917.340 68.720 917.600 68.980 ;
        RECT 1519.940 68.720 1520.200 68.980 ;
        RECT 912.740 2.760 913.000 3.020 ;
        RECT 917.340 2.760 917.600 3.020 ;
      LAYER met2 ;
        RECT 1524.465 1700.410 1524.745 1704.000 ;
        RECT 1523.220 1700.270 1524.745 1700.410 ;
        RECT 1523.220 1656.130 1523.360 1700.270 ;
        RECT 1524.465 1700.000 1524.745 1700.270 ;
        RECT 1519.480 1655.810 1519.740 1656.130 ;
        RECT 1523.160 1655.810 1523.420 1656.130 ;
        RECT 1519.540 1559.650 1519.680 1655.810 ;
        RECT 1519.080 1559.510 1519.680 1559.650 ;
        RECT 1519.080 1558.970 1519.220 1559.510 ;
        RECT 1519.080 1558.830 1519.680 1558.970 ;
        RECT 1519.540 1463.090 1519.680 1558.830 ;
        RECT 1519.080 1462.950 1519.680 1463.090 ;
        RECT 1519.080 1462.410 1519.220 1462.950 ;
        RECT 1519.080 1462.270 1519.680 1462.410 ;
        RECT 1519.540 1076.850 1519.680 1462.270 ;
        RECT 1519.080 1076.710 1519.680 1076.850 ;
        RECT 1519.080 1076.170 1519.220 1076.710 ;
        RECT 1519.080 1076.030 1519.680 1076.170 ;
        RECT 1519.540 980.290 1519.680 1076.030 ;
        RECT 1519.080 980.150 1519.680 980.290 ;
        RECT 1519.080 979.610 1519.220 980.150 ;
        RECT 1519.080 979.470 1519.680 979.610 ;
        RECT 1519.540 883.730 1519.680 979.470 ;
        RECT 1519.080 883.590 1519.680 883.730 ;
        RECT 1519.080 883.050 1519.220 883.590 ;
        RECT 1519.080 882.910 1519.680 883.050 ;
        RECT 1519.540 724.610 1519.680 882.910 ;
        RECT 1519.540 724.470 1520.140 724.610 ;
        RECT 1520.000 662.730 1520.140 724.470 ;
        RECT 1519.540 662.590 1520.140 662.730 ;
        RECT 1519.540 614.030 1519.680 662.590 ;
        RECT 1519.480 613.710 1519.740 614.030 ;
        RECT 1519.480 565.770 1519.740 566.090 ;
        RECT 1519.540 428.810 1519.680 565.770 ;
        RECT 1519.080 428.670 1519.680 428.810 ;
        RECT 1519.080 428.130 1519.220 428.670 ;
        RECT 1519.080 427.990 1519.680 428.130 ;
        RECT 1519.540 373.650 1519.680 427.990 ;
        RECT 1519.480 373.330 1519.740 373.650 ;
        RECT 1519.480 372.650 1519.740 372.970 ;
        RECT 1519.540 317.550 1519.680 372.650 ;
        RECT 1519.480 317.230 1519.740 317.550 ;
        RECT 1519.940 268.950 1520.200 269.270 ;
        RECT 1520.000 229.005 1520.140 268.950 ;
        RECT 1519.930 228.635 1520.210 229.005 ;
        RECT 1519.010 227.955 1519.290 228.325 ;
        RECT 1519.080 212.150 1519.220 227.955 ;
        RECT 1519.020 211.830 1519.280 212.150 ;
        RECT 1520.400 211.830 1520.660 212.150 ;
        RECT 1520.460 172.450 1520.600 211.830 ;
        RECT 1520.000 172.310 1520.600 172.450 ;
        RECT 1520.000 131.570 1520.140 172.310 ;
        RECT 1519.940 131.250 1520.200 131.570 ;
        RECT 1519.940 124.110 1520.200 124.430 ;
        RECT 1520.000 69.010 1520.140 124.110 ;
        RECT 917.340 68.690 917.600 69.010 ;
        RECT 1519.940 68.690 1520.200 69.010 ;
        RECT 917.400 3.050 917.540 68.690 ;
        RECT 912.740 2.730 913.000 3.050 ;
        RECT 917.340 2.730 917.600 3.050 ;
        RECT 912.800 2.400 912.940 2.730 ;
        RECT 912.590 -4.800 913.150 2.400 ;
      LAYER via2 ;
        RECT 1519.930 228.680 1520.210 228.960 ;
        RECT 1519.010 228.000 1519.290 228.280 ;
      LAYER met3 ;
        RECT 1519.905 228.970 1520.235 228.985 ;
        RECT 1518.310 228.670 1520.235 228.970 ;
        RECT 1518.310 228.290 1518.610 228.670 ;
        RECT 1519.905 228.655 1520.235 228.670 ;
        RECT 1518.985 228.290 1519.315 228.305 ;
        RECT 1518.310 227.990 1519.315 228.290 ;
        RECT 1518.985 227.975 1519.315 227.990 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 931.110 68.580 931.430 68.640 ;
        RECT 1532.790 68.580 1533.110 68.640 ;
        RECT 931.110 68.440 1533.110 68.580 ;
        RECT 931.110 68.380 931.430 68.440 ;
        RECT 1532.790 68.380 1533.110 68.440 ;
      LAYER via ;
        RECT 931.140 68.380 931.400 68.640 ;
        RECT 1532.820 68.380 1533.080 68.640 ;
      LAYER met2 ;
        RECT 1531.825 1700.000 1532.105 1704.000 ;
        RECT 1531.960 1667.090 1532.100 1700.000 ;
        RECT 1531.960 1666.950 1533.020 1667.090 ;
        RECT 1532.880 68.670 1533.020 1666.950 ;
        RECT 931.140 68.350 931.400 68.670 ;
        RECT 1532.820 68.350 1533.080 68.670 ;
        RECT 931.200 3.130 931.340 68.350 ;
        RECT 930.280 2.990 931.340 3.130 ;
        RECT 930.280 2.400 930.420 2.990 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 951.810 65.180 952.130 65.240 ;
        RECT 1539.690 65.180 1540.010 65.240 ;
        RECT 951.810 65.040 1540.010 65.180 ;
        RECT 951.810 64.980 952.130 65.040 ;
        RECT 1539.690 64.980 1540.010 65.040 ;
        RECT 948.130 2.960 948.450 3.020 ;
        RECT 951.810 2.960 952.130 3.020 ;
        RECT 948.130 2.820 952.130 2.960 ;
        RECT 948.130 2.760 948.450 2.820 ;
        RECT 951.810 2.760 952.130 2.820 ;
      LAYER via ;
        RECT 951.840 64.980 952.100 65.240 ;
        RECT 1539.720 64.980 1539.980 65.240 ;
        RECT 948.160 2.760 948.420 3.020 ;
        RECT 951.840 2.760 952.100 3.020 ;
      LAYER met2 ;
        RECT 1539.185 1700.410 1539.465 1704.000 ;
        RECT 1539.185 1700.270 1539.920 1700.410 ;
        RECT 1539.185 1700.000 1539.465 1700.270 ;
        RECT 1539.780 65.270 1539.920 1700.270 ;
        RECT 951.840 64.950 952.100 65.270 ;
        RECT 1539.720 64.950 1539.980 65.270 ;
        RECT 951.900 3.050 952.040 64.950 ;
        RECT 948.160 2.730 948.420 3.050 ;
        RECT 951.840 2.730 952.100 3.050 ;
        RECT 948.220 2.400 948.360 2.730 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 966.070 47.160 966.390 47.220 ;
        RECT 1546.130 47.160 1546.450 47.220 ;
        RECT 966.070 47.020 1546.450 47.160 ;
        RECT 966.070 46.960 966.390 47.020 ;
        RECT 1546.130 46.960 1546.450 47.020 ;
      LAYER via ;
        RECT 966.100 46.960 966.360 47.220 ;
        RECT 1546.160 46.960 1546.420 47.220 ;
      LAYER met2 ;
        RECT 1546.545 1700.410 1546.825 1704.000 ;
        RECT 1546.220 1700.270 1546.825 1700.410 ;
        RECT 1546.220 47.250 1546.360 1700.270 ;
        RECT 1546.545 1700.000 1546.825 1700.270 ;
        RECT 966.100 46.930 966.360 47.250 ;
        RECT 1546.160 46.930 1546.420 47.250 ;
        RECT 966.160 2.400 966.300 46.930 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 984.010 47.500 984.330 47.560 ;
        RECT 1553.030 47.500 1553.350 47.560 ;
        RECT 984.010 47.360 1553.350 47.500 ;
        RECT 984.010 47.300 984.330 47.360 ;
        RECT 1553.030 47.300 1553.350 47.360 ;
      LAYER via ;
        RECT 984.040 47.300 984.300 47.560 ;
        RECT 1553.060 47.300 1553.320 47.560 ;
      LAYER met2 ;
        RECT 1553.905 1700.410 1554.185 1704.000 ;
        RECT 1553.120 1700.270 1554.185 1700.410 ;
        RECT 1553.120 47.590 1553.260 1700.270 ;
        RECT 1553.905 1700.000 1554.185 1700.270 ;
        RECT 984.040 47.270 984.300 47.590 ;
        RECT 1553.060 47.270 1553.320 47.590 ;
        RECT 984.100 2.400 984.240 47.270 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1421.885 1700.410 1422.165 1704.000 ;
        RECT 1421.885 1700.270 1423.080 1700.410 ;
        RECT 1421.885 1700.000 1422.165 1700.270 ;
        RECT 1422.940 1676.100 1423.080 1700.270 ;
        RECT 1422.480 1675.960 1423.080 1676.100 ;
        RECT 1422.480 44.725 1422.620 1675.960 ;
        RECT 662.950 44.355 663.230 44.725 ;
        RECT 1422.410 44.355 1422.690 44.725 ;
        RECT 663.020 2.400 663.160 44.355 ;
        RECT 662.810 -4.800 663.370 2.400 ;
      LAYER via2 ;
        RECT 662.950 44.400 663.230 44.680 ;
        RECT 1422.410 44.400 1422.690 44.680 ;
      LAYER met3 ;
        RECT 662.925 44.690 663.255 44.705 ;
        RECT 1422.385 44.690 1422.715 44.705 ;
        RECT 662.925 44.390 1422.715 44.690 ;
        RECT 662.925 44.375 663.255 44.390 ;
        RECT 1422.385 44.375 1422.715 44.390 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1001.950 47.840 1002.270 47.900 ;
        RECT 1559.930 47.840 1560.250 47.900 ;
        RECT 1001.950 47.700 1560.250 47.840 ;
        RECT 1001.950 47.640 1002.270 47.700 ;
        RECT 1559.930 47.640 1560.250 47.700 ;
      LAYER via ;
        RECT 1001.980 47.640 1002.240 47.900 ;
        RECT 1559.960 47.640 1560.220 47.900 ;
      LAYER met2 ;
        RECT 1561.265 1700.410 1561.545 1704.000 ;
        RECT 1560.020 1700.270 1561.545 1700.410 ;
        RECT 1560.020 47.930 1560.160 1700.270 ;
        RECT 1561.265 1700.000 1561.545 1700.270 ;
        RECT 1001.980 47.610 1002.240 47.930 ;
        RECT 1559.960 47.610 1560.220 47.930 ;
        RECT 1002.040 2.400 1002.180 47.610 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1019.430 48.180 1019.750 48.240 ;
        RECT 1566.830 48.180 1567.150 48.240 ;
        RECT 1019.430 48.040 1567.150 48.180 ;
        RECT 1019.430 47.980 1019.750 48.040 ;
        RECT 1566.830 47.980 1567.150 48.040 ;
      LAYER via ;
        RECT 1019.460 47.980 1019.720 48.240 ;
        RECT 1566.860 47.980 1567.120 48.240 ;
      LAYER met2 ;
        RECT 1568.625 1700.410 1568.905 1704.000 ;
        RECT 1566.920 1700.270 1568.905 1700.410 ;
        RECT 1566.920 48.270 1567.060 1700.270 ;
        RECT 1568.625 1700.000 1568.905 1700.270 ;
        RECT 1019.460 47.950 1019.720 48.270 ;
        RECT 1566.860 47.950 1567.120 48.270 ;
        RECT 1019.520 2.400 1019.660 47.950 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1037.370 44.440 1037.690 44.500 ;
        RECT 1574.650 44.440 1574.970 44.500 ;
        RECT 1037.370 44.300 1574.970 44.440 ;
        RECT 1037.370 44.240 1037.690 44.300 ;
        RECT 1574.650 44.240 1574.970 44.300 ;
      LAYER via ;
        RECT 1037.400 44.240 1037.660 44.500 ;
        RECT 1574.680 44.240 1574.940 44.500 ;
      LAYER met2 ;
        RECT 1575.985 1700.410 1576.265 1704.000 ;
        RECT 1574.740 1700.270 1576.265 1700.410 ;
        RECT 1574.740 44.530 1574.880 1700.270 ;
        RECT 1575.985 1700.000 1576.265 1700.270 ;
        RECT 1037.400 44.210 1037.660 44.530 ;
        RECT 1574.680 44.210 1574.940 44.530 ;
        RECT 1037.460 2.400 1037.600 44.210 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1580.630 1687.320 1580.950 1687.380 ;
        RECT 1581.550 1687.320 1581.870 1687.380 ;
        RECT 1580.630 1687.180 1581.870 1687.320 ;
        RECT 1580.630 1687.120 1580.950 1687.180 ;
        RECT 1581.550 1687.120 1581.870 1687.180 ;
        RECT 1054.850 44.100 1055.170 44.160 ;
        RECT 1580.630 44.100 1580.950 44.160 ;
        RECT 1054.850 43.960 1580.950 44.100 ;
        RECT 1054.850 43.900 1055.170 43.960 ;
        RECT 1580.630 43.900 1580.950 43.960 ;
      LAYER via ;
        RECT 1580.660 1687.120 1580.920 1687.380 ;
        RECT 1581.580 1687.120 1581.840 1687.380 ;
        RECT 1054.880 43.900 1055.140 44.160 ;
        RECT 1580.660 43.900 1580.920 44.160 ;
      LAYER met2 ;
        RECT 1583.345 1700.410 1583.625 1704.000 ;
        RECT 1581.640 1700.270 1583.625 1700.410 ;
        RECT 1581.640 1687.410 1581.780 1700.270 ;
        RECT 1583.345 1700.000 1583.625 1700.270 ;
        RECT 1580.660 1687.090 1580.920 1687.410 ;
        RECT 1581.580 1687.090 1581.840 1687.410 ;
        RECT 1580.720 44.190 1580.860 1687.090 ;
        RECT 1054.880 43.870 1055.140 44.190 ;
        RECT 1580.660 43.870 1580.920 44.190 ;
        RECT 1054.940 17.410 1055.080 43.870 ;
        RECT 1054.940 17.270 1055.540 17.410 ;
        RECT 1055.400 2.400 1055.540 17.270 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1588.525 476.085 1588.695 517.055 ;
      LAYER mcon ;
        RECT 1588.525 516.885 1588.695 517.055 ;
      LAYER met1 ;
        RECT 1587.530 1531.940 1587.850 1532.000 ;
        RECT 1588.450 1531.940 1588.770 1532.000 ;
        RECT 1587.530 1531.800 1588.770 1531.940 ;
        RECT 1587.530 1531.740 1587.850 1531.800 ;
        RECT 1588.450 1531.740 1588.770 1531.800 ;
        RECT 1587.530 1097.080 1587.850 1097.140 ;
        RECT 1588.450 1097.080 1588.770 1097.140 ;
        RECT 1587.530 1096.940 1588.770 1097.080 ;
        RECT 1587.530 1096.880 1587.850 1096.940 ;
        RECT 1588.450 1096.880 1588.770 1096.940 ;
        RECT 1587.530 1049.140 1587.850 1049.200 ;
        RECT 1588.450 1049.140 1588.770 1049.200 ;
        RECT 1587.530 1049.000 1588.770 1049.140 ;
        RECT 1587.530 1048.940 1587.850 1049.000 ;
        RECT 1588.450 1048.940 1588.770 1049.000 ;
        RECT 1587.530 1000.520 1587.850 1000.580 ;
        RECT 1588.450 1000.520 1588.770 1000.580 ;
        RECT 1587.530 1000.380 1588.770 1000.520 ;
        RECT 1587.530 1000.320 1587.850 1000.380 ;
        RECT 1588.450 1000.320 1588.770 1000.380 ;
        RECT 1587.530 952.580 1587.850 952.640 ;
        RECT 1588.450 952.580 1588.770 952.640 ;
        RECT 1587.530 952.440 1588.770 952.580 ;
        RECT 1587.530 952.380 1587.850 952.440 ;
        RECT 1588.450 952.380 1588.770 952.440 ;
        RECT 1587.530 903.960 1587.850 904.020 ;
        RECT 1588.450 903.960 1588.770 904.020 ;
        RECT 1587.530 903.820 1588.770 903.960 ;
        RECT 1587.530 903.760 1587.850 903.820 ;
        RECT 1588.450 903.760 1588.770 903.820 ;
        RECT 1588.450 517.040 1588.770 517.100 ;
        RECT 1588.255 516.900 1588.770 517.040 ;
        RECT 1588.450 516.840 1588.770 516.900 ;
        RECT 1588.465 476.240 1588.755 476.285 ;
        RECT 1588.910 476.240 1589.230 476.300 ;
        RECT 1588.465 476.100 1589.230 476.240 ;
        RECT 1588.465 476.055 1588.755 476.100 ;
        RECT 1588.910 476.040 1589.230 476.100 ;
        RECT 1588.910 448.500 1589.230 448.760 ;
        RECT 1589.000 448.020 1589.140 448.500 ;
        RECT 1589.370 448.020 1589.690 448.080 ;
        RECT 1589.000 447.880 1589.690 448.020 ;
        RECT 1589.370 447.820 1589.690 447.880 ;
        RECT 1588.450 379.680 1588.770 379.740 ;
        RECT 1589.830 379.680 1590.150 379.740 ;
        RECT 1588.450 379.540 1590.150 379.680 ;
        RECT 1588.450 379.480 1588.770 379.540 ;
        RECT 1589.830 379.480 1590.150 379.540 ;
        RECT 1587.530 276.320 1587.850 276.380 ;
        RECT 1588.450 276.320 1588.770 276.380 ;
        RECT 1587.530 276.180 1588.770 276.320 ;
        RECT 1587.530 276.120 1587.850 276.180 ;
        RECT 1588.450 276.120 1588.770 276.180 ;
        RECT 1587.530 227.700 1587.850 227.760 ;
        RECT 1588.450 227.700 1588.770 227.760 ;
        RECT 1587.530 227.560 1588.770 227.700 ;
        RECT 1587.530 227.500 1587.850 227.560 ;
        RECT 1588.450 227.500 1588.770 227.560 ;
        RECT 1587.530 159.020 1587.850 159.080 ;
        RECT 1588.450 159.020 1588.770 159.080 ;
        RECT 1587.530 158.880 1588.770 159.020 ;
        RECT 1587.530 158.820 1587.850 158.880 ;
        RECT 1588.450 158.820 1588.770 158.880 ;
        RECT 1073.250 43.760 1073.570 43.820 ;
        RECT 1587.530 43.760 1587.850 43.820 ;
        RECT 1073.250 43.620 1587.850 43.760 ;
        RECT 1073.250 43.560 1073.570 43.620 ;
        RECT 1587.530 43.560 1587.850 43.620 ;
      LAYER via ;
        RECT 1587.560 1531.740 1587.820 1532.000 ;
        RECT 1588.480 1531.740 1588.740 1532.000 ;
        RECT 1587.560 1096.880 1587.820 1097.140 ;
        RECT 1588.480 1096.880 1588.740 1097.140 ;
        RECT 1587.560 1048.940 1587.820 1049.200 ;
        RECT 1588.480 1048.940 1588.740 1049.200 ;
        RECT 1587.560 1000.320 1587.820 1000.580 ;
        RECT 1588.480 1000.320 1588.740 1000.580 ;
        RECT 1587.560 952.380 1587.820 952.640 ;
        RECT 1588.480 952.380 1588.740 952.640 ;
        RECT 1587.560 903.760 1587.820 904.020 ;
        RECT 1588.480 903.760 1588.740 904.020 ;
        RECT 1588.480 516.840 1588.740 517.100 ;
        RECT 1588.940 476.040 1589.200 476.300 ;
        RECT 1588.940 448.500 1589.200 448.760 ;
        RECT 1589.400 447.820 1589.660 448.080 ;
        RECT 1588.480 379.480 1588.740 379.740 ;
        RECT 1589.860 379.480 1590.120 379.740 ;
        RECT 1587.560 276.120 1587.820 276.380 ;
        RECT 1588.480 276.120 1588.740 276.380 ;
        RECT 1587.560 227.500 1587.820 227.760 ;
        RECT 1588.480 227.500 1588.740 227.760 ;
        RECT 1587.560 158.820 1587.820 159.080 ;
        RECT 1588.480 158.820 1588.740 159.080 ;
        RECT 1073.280 43.560 1073.540 43.820 ;
        RECT 1587.560 43.560 1587.820 43.820 ;
      LAYER met2 ;
        RECT 1590.705 1700.410 1590.985 1704.000 ;
        RECT 1589.460 1700.270 1590.985 1700.410 ;
        RECT 1589.460 1688.850 1589.600 1700.270 ;
        RECT 1590.705 1700.000 1590.985 1700.270 ;
        RECT 1588.540 1688.710 1589.600 1688.850 ;
        RECT 1588.540 1532.030 1588.680 1688.710 ;
        RECT 1587.560 1531.710 1587.820 1532.030 ;
        RECT 1588.480 1531.710 1588.740 1532.030 ;
        RECT 1587.620 1097.170 1587.760 1531.710 ;
        RECT 1587.560 1096.850 1587.820 1097.170 ;
        RECT 1588.480 1096.850 1588.740 1097.170 ;
        RECT 1588.540 1049.230 1588.680 1096.850 ;
        RECT 1587.560 1048.910 1587.820 1049.230 ;
        RECT 1588.480 1048.910 1588.740 1049.230 ;
        RECT 1587.620 1000.610 1587.760 1048.910 ;
        RECT 1587.560 1000.290 1587.820 1000.610 ;
        RECT 1588.480 1000.290 1588.740 1000.610 ;
        RECT 1588.540 952.670 1588.680 1000.290 ;
        RECT 1587.560 952.350 1587.820 952.670 ;
        RECT 1588.480 952.350 1588.740 952.670 ;
        RECT 1587.620 904.050 1587.760 952.350 ;
        RECT 1587.560 903.730 1587.820 904.050 ;
        RECT 1588.480 903.730 1588.740 904.050 ;
        RECT 1588.540 517.130 1588.680 903.730 ;
        RECT 1588.480 516.810 1588.740 517.130 ;
        RECT 1588.940 476.010 1589.200 476.330 ;
        RECT 1589.000 448.790 1589.140 476.010 ;
        RECT 1588.940 448.470 1589.200 448.790 ;
        RECT 1589.400 447.790 1589.660 448.110 ;
        RECT 1589.460 427.450 1589.600 447.790 ;
        RECT 1589.460 427.310 1590.060 427.450 ;
        RECT 1589.920 379.770 1590.060 427.310 ;
        RECT 1588.480 379.450 1588.740 379.770 ;
        RECT 1589.860 379.450 1590.120 379.770 ;
        RECT 1588.540 276.410 1588.680 379.450 ;
        RECT 1587.560 276.090 1587.820 276.410 ;
        RECT 1588.480 276.090 1588.740 276.410 ;
        RECT 1587.620 227.790 1587.760 276.090 ;
        RECT 1587.560 227.470 1587.820 227.790 ;
        RECT 1588.480 227.470 1588.740 227.790 ;
        RECT 1588.540 159.110 1588.680 227.470 ;
        RECT 1587.560 158.790 1587.820 159.110 ;
        RECT 1588.480 158.790 1588.740 159.110 ;
        RECT 1587.620 43.850 1587.760 158.790 ;
        RECT 1073.280 43.530 1073.540 43.850 ;
        RECT 1587.560 43.530 1587.820 43.850 ;
        RECT 1073.340 2.400 1073.480 43.530 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1594.430 1687.320 1594.750 1687.380 ;
        RECT 1596.270 1687.320 1596.590 1687.380 ;
        RECT 1594.430 1687.180 1596.590 1687.320 ;
        RECT 1594.430 1687.120 1594.750 1687.180 ;
        RECT 1596.270 1687.120 1596.590 1687.180 ;
        RECT 1090.730 43.420 1091.050 43.480 ;
        RECT 1594.430 43.420 1594.750 43.480 ;
        RECT 1090.730 43.280 1594.750 43.420 ;
        RECT 1090.730 43.220 1091.050 43.280 ;
        RECT 1594.430 43.220 1594.750 43.280 ;
      LAYER via ;
        RECT 1594.460 1687.120 1594.720 1687.380 ;
        RECT 1596.300 1687.120 1596.560 1687.380 ;
        RECT 1090.760 43.220 1091.020 43.480 ;
        RECT 1594.460 43.220 1594.720 43.480 ;
      LAYER met2 ;
        RECT 1598.065 1700.410 1598.345 1704.000 ;
        RECT 1596.360 1700.270 1598.345 1700.410 ;
        RECT 1596.360 1687.410 1596.500 1700.270 ;
        RECT 1598.065 1700.000 1598.345 1700.270 ;
        RECT 1594.460 1687.090 1594.720 1687.410 ;
        RECT 1596.300 1687.090 1596.560 1687.410 ;
        RECT 1594.520 43.510 1594.660 1687.090 ;
        RECT 1090.760 43.190 1091.020 43.510 ;
        RECT 1594.460 43.190 1594.720 43.510 ;
        RECT 1090.820 2.400 1090.960 43.190 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1600.870 1687.320 1601.190 1687.380 ;
        RECT 1603.630 1687.320 1603.950 1687.380 ;
        RECT 1600.870 1687.180 1603.950 1687.320 ;
        RECT 1600.870 1687.120 1601.190 1687.180 ;
        RECT 1603.630 1687.120 1603.950 1687.180 ;
        RECT 1108.670 43.080 1108.990 43.140 ;
        RECT 1600.870 43.080 1601.190 43.140 ;
        RECT 1108.670 42.940 1601.190 43.080 ;
        RECT 1108.670 42.880 1108.990 42.940 ;
        RECT 1600.870 42.880 1601.190 42.940 ;
      LAYER via ;
        RECT 1600.900 1687.120 1601.160 1687.380 ;
        RECT 1603.660 1687.120 1603.920 1687.380 ;
        RECT 1108.700 42.880 1108.960 43.140 ;
        RECT 1600.900 42.880 1601.160 43.140 ;
      LAYER met2 ;
        RECT 1605.425 1700.410 1605.705 1704.000 ;
        RECT 1603.720 1700.270 1605.705 1700.410 ;
        RECT 1603.720 1687.410 1603.860 1700.270 ;
        RECT 1605.425 1700.000 1605.705 1700.270 ;
        RECT 1600.900 1687.090 1601.160 1687.410 ;
        RECT 1603.660 1687.090 1603.920 1687.410 ;
        RECT 1600.960 43.170 1601.100 1687.090 ;
        RECT 1108.700 42.850 1108.960 43.170 ;
        RECT 1600.900 42.850 1601.160 43.170 ;
        RECT 1108.760 2.400 1108.900 42.850 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1608.230 1678.140 1608.550 1678.200 ;
        RECT 1610.990 1678.140 1611.310 1678.200 ;
        RECT 1608.230 1678.000 1611.310 1678.140 ;
        RECT 1608.230 1677.940 1608.550 1678.000 ;
        RECT 1610.990 1677.940 1611.310 1678.000 ;
        RECT 1126.610 42.740 1126.930 42.800 ;
        RECT 1608.230 42.740 1608.550 42.800 ;
        RECT 1126.610 42.600 1608.550 42.740 ;
        RECT 1126.610 42.540 1126.930 42.600 ;
        RECT 1608.230 42.540 1608.550 42.600 ;
      LAYER via ;
        RECT 1608.260 1677.940 1608.520 1678.200 ;
        RECT 1611.020 1677.940 1611.280 1678.200 ;
        RECT 1126.640 42.540 1126.900 42.800 ;
        RECT 1608.260 42.540 1608.520 42.800 ;
      LAYER met2 ;
        RECT 1612.785 1700.410 1613.065 1704.000 ;
        RECT 1611.080 1700.270 1613.065 1700.410 ;
        RECT 1611.080 1678.230 1611.220 1700.270 ;
        RECT 1612.785 1700.000 1613.065 1700.270 ;
        RECT 1608.260 1677.910 1608.520 1678.230 ;
        RECT 1611.020 1677.910 1611.280 1678.230 ;
        RECT 1608.320 42.830 1608.460 1677.910 ;
        RECT 1126.640 42.510 1126.900 42.830 ;
        RECT 1608.260 42.510 1608.520 42.830 ;
        RECT 1126.700 2.400 1126.840 42.510 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1616.585 1635.485 1616.755 1683.595 ;
        RECT 1616.125 1497.445 1616.295 1521.415 ;
        RECT 1616.585 1338.665 1616.755 1366.715 ;
        RECT 1617.045 1248.905 1617.215 1269.815 ;
        RECT 1617.045 476.085 1617.215 540.175 ;
        RECT 1617.045 282.965 1617.215 331.075 ;
        RECT 1616.585 186.405 1616.755 234.515 ;
      LAYER mcon ;
        RECT 1616.585 1683.425 1616.755 1683.595 ;
        RECT 1616.125 1521.245 1616.295 1521.415 ;
        RECT 1616.585 1366.545 1616.755 1366.715 ;
        RECT 1617.045 1269.645 1617.215 1269.815 ;
        RECT 1617.045 540.005 1617.215 540.175 ;
        RECT 1617.045 330.905 1617.215 331.075 ;
        RECT 1616.585 234.345 1616.755 234.515 ;
      LAYER met1 ;
        RECT 1616.525 1683.580 1616.815 1683.625 ;
        RECT 1618.350 1683.580 1618.670 1683.640 ;
        RECT 1616.525 1683.440 1618.670 1683.580 ;
        RECT 1616.525 1683.395 1616.815 1683.440 ;
        RECT 1618.350 1683.380 1618.670 1683.440 ;
        RECT 1616.510 1635.640 1616.830 1635.700 ;
        RECT 1616.315 1635.500 1616.830 1635.640 ;
        RECT 1616.510 1635.440 1616.830 1635.500 ;
        RECT 1616.510 1559.820 1616.830 1559.880 ;
        RECT 1616.140 1559.680 1616.830 1559.820 ;
        RECT 1616.140 1559.540 1616.280 1559.680 ;
        RECT 1616.510 1559.620 1616.830 1559.680 ;
        RECT 1616.050 1559.280 1616.370 1559.540 ;
        RECT 1616.050 1521.400 1616.370 1521.460 ;
        RECT 1615.855 1521.260 1616.370 1521.400 ;
        RECT 1616.050 1521.200 1616.370 1521.260 ;
        RECT 1616.065 1497.600 1616.355 1497.645 ;
        RECT 1616.510 1497.600 1616.830 1497.660 ;
        RECT 1616.065 1497.460 1616.830 1497.600 ;
        RECT 1616.065 1497.415 1616.355 1497.460 ;
        RECT 1616.510 1497.400 1616.830 1497.460 ;
        RECT 1616.510 1435.380 1616.830 1435.440 ;
        RECT 1617.430 1435.380 1617.750 1435.440 ;
        RECT 1616.510 1435.240 1617.750 1435.380 ;
        RECT 1616.510 1435.180 1616.830 1435.240 ;
        RECT 1617.430 1435.180 1617.750 1435.240 ;
        RECT 1616.510 1366.700 1616.830 1366.760 ;
        RECT 1616.315 1366.560 1616.830 1366.700 ;
        RECT 1616.510 1366.500 1616.830 1366.560 ;
        RECT 1616.510 1338.820 1616.830 1338.880 ;
        RECT 1616.315 1338.680 1616.830 1338.820 ;
        RECT 1616.510 1338.620 1616.830 1338.680 ;
        RECT 1616.510 1269.800 1616.830 1269.860 ;
        RECT 1616.985 1269.800 1617.275 1269.845 ;
        RECT 1616.510 1269.660 1617.275 1269.800 ;
        RECT 1616.510 1269.600 1616.830 1269.660 ;
        RECT 1616.985 1269.615 1617.275 1269.660 ;
        RECT 1616.970 1249.060 1617.290 1249.120 ;
        RECT 1616.775 1248.920 1617.290 1249.060 ;
        RECT 1616.970 1248.860 1617.290 1248.920 ;
        RECT 1616.970 1169.500 1617.290 1169.560 ;
        RECT 1617.890 1169.500 1618.210 1169.560 ;
        RECT 1616.970 1169.360 1618.210 1169.500 ;
        RECT 1616.970 1169.300 1617.290 1169.360 ;
        RECT 1617.890 1169.300 1618.210 1169.360 ;
        RECT 1616.510 869.620 1616.830 869.680 ;
        RECT 1617.430 869.620 1617.750 869.680 ;
        RECT 1616.510 869.480 1617.750 869.620 ;
        RECT 1616.510 869.420 1616.830 869.480 ;
        RECT 1617.430 869.420 1617.750 869.480 ;
        RECT 1616.970 724.440 1617.290 724.500 ;
        RECT 1617.430 724.440 1617.750 724.500 ;
        RECT 1616.970 724.300 1617.750 724.440 ;
        RECT 1616.970 724.240 1617.290 724.300 ;
        RECT 1617.430 724.240 1617.750 724.300 ;
        RECT 1616.970 540.160 1617.290 540.220 ;
        RECT 1616.775 540.020 1617.290 540.160 ;
        RECT 1616.970 539.960 1617.290 540.020 ;
        RECT 1616.970 476.240 1617.290 476.300 ;
        RECT 1616.775 476.100 1617.290 476.240 ;
        RECT 1616.970 476.040 1617.290 476.100 ;
        RECT 1616.510 434.760 1616.830 434.820 ;
        RECT 1616.970 434.760 1617.290 434.820 ;
        RECT 1616.510 434.620 1617.290 434.760 ;
        RECT 1616.510 434.560 1616.830 434.620 ;
        RECT 1616.970 434.560 1617.290 434.620 ;
        RECT 1616.970 331.060 1617.290 331.120 ;
        RECT 1616.775 330.920 1617.290 331.060 ;
        RECT 1616.970 330.860 1617.290 330.920 ;
        RECT 1616.970 283.120 1617.290 283.180 ;
        RECT 1616.775 282.980 1617.290 283.120 ;
        RECT 1616.970 282.920 1617.290 282.980 ;
        RECT 1616.510 241.300 1616.830 241.360 ;
        RECT 1616.970 241.300 1617.290 241.360 ;
        RECT 1616.510 241.160 1617.290 241.300 ;
        RECT 1616.510 241.100 1616.830 241.160 ;
        RECT 1616.970 241.100 1617.290 241.160 ;
        RECT 1616.510 234.500 1616.830 234.560 ;
        RECT 1616.315 234.360 1616.830 234.500 ;
        RECT 1616.510 234.300 1616.830 234.360 ;
        RECT 1616.510 186.560 1616.830 186.620 ;
        RECT 1616.315 186.420 1616.830 186.560 ;
        RECT 1616.510 186.360 1616.830 186.420 ;
        RECT 1616.510 144.740 1616.830 144.800 ;
        RECT 1616.970 144.740 1617.290 144.800 ;
        RECT 1616.510 144.600 1617.290 144.740 ;
        RECT 1616.510 144.540 1616.830 144.600 ;
        RECT 1616.970 144.540 1617.290 144.600 ;
        RECT 1144.550 42.400 1144.870 42.460 ;
        RECT 1616.510 42.400 1616.830 42.460 ;
        RECT 1144.550 42.260 1616.830 42.400 ;
        RECT 1144.550 42.200 1144.870 42.260 ;
        RECT 1616.510 42.200 1616.830 42.260 ;
      LAYER via ;
        RECT 1618.380 1683.380 1618.640 1683.640 ;
        RECT 1616.540 1635.440 1616.800 1635.700 ;
        RECT 1616.540 1559.620 1616.800 1559.880 ;
        RECT 1616.080 1559.280 1616.340 1559.540 ;
        RECT 1616.080 1521.200 1616.340 1521.460 ;
        RECT 1616.540 1497.400 1616.800 1497.660 ;
        RECT 1616.540 1435.180 1616.800 1435.440 ;
        RECT 1617.460 1435.180 1617.720 1435.440 ;
        RECT 1616.540 1366.500 1616.800 1366.760 ;
        RECT 1616.540 1338.620 1616.800 1338.880 ;
        RECT 1616.540 1269.600 1616.800 1269.860 ;
        RECT 1617.000 1248.860 1617.260 1249.120 ;
        RECT 1617.000 1169.300 1617.260 1169.560 ;
        RECT 1617.920 1169.300 1618.180 1169.560 ;
        RECT 1616.540 869.420 1616.800 869.680 ;
        RECT 1617.460 869.420 1617.720 869.680 ;
        RECT 1617.000 724.240 1617.260 724.500 ;
        RECT 1617.460 724.240 1617.720 724.500 ;
        RECT 1617.000 539.960 1617.260 540.220 ;
        RECT 1617.000 476.040 1617.260 476.300 ;
        RECT 1616.540 434.560 1616.800 434.820 ;
        RECT 1617.000 434.560 1617.260 434.820 ;
        RECT 1617.000 330.860 1617.260 331.120 ;
        RECT 1617.000 282.920 1617.260 283.180 ;
        RECT 1616.540 241.100 1616.800 241.360 ;
        RECT 1617.000 241.100 1617.260 241.360 ;
        RECT 1616.540 234.300 1616.800 234.560 ;
        RECT 1616.540 186.360 1616.800 186.620 ;
        RECT 1616.540 144.540 1616.800 144.800 ;
        RECT 1617.000 144.540 1617.260 144.800 ;
        RECT 1144.580 42.200 1144.840 42.460 ;
        RECT 1616.540 42.200 1616.800 42.460 ;
      LAYER met2 ;
        RECT 1620.145 1700.410 1620.425 1704.000 ;
        RECT 1618.440 1700.270 1620.425 1700.410 ;
        RECT 1618.440 1683.670 1618.580 1700.270 ;
        RECT 1620.145 1700.000 1620.425 1700.270 ;
        RECT 1618.380 1683.350 1618.640 1683.670 ;
        RECT 1616.540 1635.410 1616.800 1635.730 ;
        RECT 1616.600 1559.910 1616.740 1635.410 ;
        RECT 1616.540 1559.590 1616.800 1559.910 ;
        RECT 1616.080 1559.250 1616.340 1559.570 ;
        RECT 1616.140 1521.490 1616.280 1559.250 ;
        RECT 1616.080 1521.170 1616.340 1521.490 ;
        RECT 1616.540 1497.370 1616.800 1497.690 ;
        RECT 1616.600 1483.605 1616.740 1497.370 ;
        RECT 1616.530 1483.235 1616.810 1483.605 ;
        RECT 1617.450 1483.235 1617.730 1483.605 ;
        RECT 1617.520 1435.470 1617.660 1483.235 ;
        RECT 1616.540 1435.210 1616.800 1435.470 ;
        RECT 1616.540 1435.150 1617.200 1435.210 ;
        RECT 1617.460 1435.150 1617.720 1435.470 ;
        RECT 1616.600 1435.070 1617.200 1435.150 ;
        RECT 1617.060 1401.210 1617.200 1435.070 ;
        RECT 1617.060 1401.070 1617.660 1401.210 ;
        RECT 1617.520 1399.850 1617.660 1401.070 ;
        RECT 1616.600 1399.710 1617.660 1399.850 ;
        RECT 1616.600 1366.790 1616.740 1399.710 ;
        RECT 1616.540 1366.470 1616.800 1366.790 ;
        RECT 1616.540 1338.590 1616.800 1338.910 ;
        RECT 1616.600 1304.650 1616.740 1338.590 ;
        RECT 1616.600 1304.510 1617.200 1304.650 ;
        RECT 1617.060 1297.170 1617.200 1304.510 ;
        RECT 1616.600 1297.030 1617.200 1297.170 ;
        RECT 1616.600 1269.890 1616.740 1297.030 ;
        RECT 1616.540 1269.570 1616.800 1269.890 ;
        RECT 1617.000 1248.830 1617.260 1249.150 ;
        RECT 1617.060 1169.590 1617.200 1248.830 ;
        RECT 1617.000 1169.270 1617.260 1169.590 ;
        RECT 1617.920 1169.270 1618.180 1169.590 ;
        RECT 1617.980 1145.645 1618.120 1169.270 ;
        RECT 1616.990 1145.275 1617.270 1145.645 ;
        RECT 1617.910 1145.275 1618.190 1145.645 ;
        RECT 1617.060 1000.635 1617.200 1145.275 ;
        RECT 1616.990 1000.265 1617.270 1000.635 ;
        RECT 1616.990 999.075 1617.270 999.445 ;
        RECT 1617.060 952.410 1617.200 999.075 ;
        RECT 1617.060 952.270 1617.660 952.410 ;
        RECT 1617.520 869.710 1617.660 952.270 ;
        RECT 1616.540 869.390 1616.800 869.710 ;
        RECT 1617.460 869.390 1617.720 869.710 ;
        RECT 1616.600 821.170 1616.740 869.390 ;
        RECT 1616.600 821.030 1617.200 821.170 ;
        RECT 1617.060 787.170 1617.200 821.030 ;
        RECT 1617.060 787.030 1617.660 787.170 ;
        RECT 1617.520 776.290 1617.660 787.030 ;
        RECT 1617.060 776.150 1617.660 776.290 ;
        RECT 1617.060 724.530 1617.200 776.150 ;
        RECT 1617.000 724.210 1617.260 724.530 ;
        RECT 1617.460 724.210 1617.720 724.530 ;
        RECT 1617.520 676.445 1617.660 724.210 ;
        RECT 1616.530 676.075 1616.810 676.445 ;
        RECT 1617.450 676.075 1617.730 676.445 ;
        RECT 1616.600 628.050 1616.740 676.075 ;
        RECT 1616.600 627.910 1617.200 628.050 ;
        RECT 1617.060 594.050 1617.200 627.910 ;
        RECT 1617.060 593.910 1617.660 594.050 ;
        RECT 1617.520 590.650 1617.660 593.910 ;
        RECT 1617.060 590.510 1617.660 590.650 ;
        RECT 1617.060 540.250 1617.200 590.510 ;
        RECT 1617.000 539.930 1617.260 540.250 ;
        RECT 1617.000 476.010 1617.260 476.330 ;
        RECT 1617.060 434.850 1617.200 476.010 ;
        RECT 1616.540 434.530 1616.800 434.850 ;
        RECT 1617.000 434.530 1617.260 434.850 ;
        RECT 1616.600 362.170 1616.740 434.530 ;
        RECT 1616.600 362.030 1617.200 362.170 ;
        RECT 1617.060 331.150 1617.200 362.030 ;
        RECT 1617.000 330.830 1617.260 331.150 ;
        RECT 1617.000 282.890 1617.260 283.210 ;
        RECT 1617.060 241.390 1617.200 282.890 ;
        RECT 1616.540 241.070 1616.800 241.390 ;
        RECT 1617.000 241.070 1617.260 241.390 ;
        RECT 1616.600 234.590 1616.740 241.070 ;
        RECT 1616.540 234.270 1616.800 234.590 ;
        RECT 1616.540 186.330 1616.800 186.650 ;
        RECT 1616.600 169.050 1616.740 186.330 ;
        RECT 1616.600 168.910 1617.660 169.050 ;
        RECT 1617.520 158.170 1617.660 168.910 ;
        RECT 1617.060 158.030 1617.660 158.170 ;
        RECT 1617.060 144.830 1617.200 158.030 ;
        RECT 1616.540 144.510 1616.800 144.830 ;
        RECT 1617.000 144.510 1617.260 144.830 ;
        RECT 1616.600 42.490 1616.740 144.510 ;
        RECT 1144.580 42.170 1144.840 42.490 ;
        RECT 1616.540 42.170 1616.800 42.490 ;
        RECT 1144.640 2.400 1144.780 42.170 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
      LAYER via2 ;
        RECT 1616.530 1483.280 1616.810 1483.560 ;
        RECT 1617.450 1483.280 1617.730 1483.560 ;
        RECT 1616.990 1145.320 1617.270 1145.600 ;
        RECT 1617.910 1145.320 1618.190 1145.600 ;
        RECT 1616.990 1000.310 1617.270 1000.590 ;
        RECT 1616.990 999.120 1617.270 999.400 ;
        RECT 1616.530 676.120 1616.810 676.400 ;
        RECT 1617.450 676.120 1617.730 676.400 ;
      LAYER met3 ;
        RECT 1616.505 1483.570 1616.835 1483.585 ;
        RECT 1617.425 1483.570 1617.755 1483.585 ;
        RECT 1616.505 1483.270 1617.755 1483.570 ;
        RECT 1616.505 1483.255 1616.835 1483.270 ;
        RECT 1617.425 1483.255 1617.755 1483.270 ;
        RECT 1616.965 1145.610 1617.295 1145.625 ;
        RECT 1617.885 1145.610 1618.215 1145.625 ;
        RECT 1616.965 1145.310 1618.215 1145.610 ;
        RECT 1616.965 1145.295 1617.295 1145.310 ;
        RECT 1617.885 1145.295 1618.215 1145.310 ;
        RECT 1616.965 1000.600 1617.295 1000.615 ;
        RECT 1616.965 1000.300 1617.970 1000.600 ;
        RECT 1616.965 1000.285 1617.295 1000.300 ;
        RECT 1616.965 999.410 1617.295 999.425 ;
        RECT 1617.670 999.410 1617.970 1000.300 ;
        RECT 1616.965 999.110 1617.970 999.410 ;
        RECT 1616.965 999.095 1617.295 999.110 ;
        RECT 1616.505 676.410 1616.835 676.425 ;
        RECT 1617.425 676.410 1617.755 676.425 ;
        RECT 1616.505 676.110 1617.755 676.410 ;
        RECT 1616.505 676.095 1616.835 676.110 ;
        RECT 1617.425 676.095 1617.755 676.110 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1623.485 1449.165 1623.655 1497.275 ;
        RECT 1623.025 1290.385 1623.195 1304.495 ;
        RECT 1623.025 965.685 1623.195 1007.335 ;
        RECT 1623.945 669.545 1624.115 699.635 ;
        RECT 1623.025 565.845 1623.195 613.955 ;
        RECT 1623.025 476.085 1623.195 524.195 ;
      LAYER mcon ;
        RECT 1623.485 1497.105 1623.655 1497.275 ;
        RECT 1623.025 1304.325 1623.195 1304.495 ;
        RECT 1623.025 1007.165 1623.195 1007.335 ;
        RECT 1623.945 699.465 1624.115 699.635 ;
        RECT 1623.025 613.785 1623.195 613.955 ;
        RECT 1623.025 524.025 1623.195 524.195 ;
      LAYER met1 ;
        RECT 1623.410 1635.640 1623.730 1635.700 ;
        RECT 1625.250 1635.640 1625.570 1635.700 ;
        RECT 1623.410 1635.500 1625.570 1635.640 ;
        RECT 1623.410 1635.440 1623.730 1635.500 ;
        RECT 1625.250 1635.440 1625.570 1635.500 ;
        RECT 1623.410 1497.260 1623.730 1497.320 ;
        RECT 1623.215 1497.120 1623.730 1497.260 ;
        RECT 1623.410 1497.060 1623.730 1497.120 ;
        RECT 1623.410 1449.320 1623.730 1449.380 ;
        RECT 1623.215 1449.180 1623.730 1449.320 ;
        RECT 1623.410 1449.120 1623.730 1449.180 ;
        RECT 1622.490 1339.160 1622.810 1339.220 ;
        RECT 1623.410 1339.160 1623.730 1339.220 ;
        RECT 1622.490 1339.020 1623.730 1339.160 ;
        RECT 1622.490 1338.960 1622.810 1339.020 ;
        RECT 1623.410 1338.960 1623.730 1339.020 ;
        RECT 1622.950 1304.480 1623.270 1304.540 ;
        RECT 1622.755 1304.340 1623.270 1304.480 ;
        RECT 1622.950 1304.280 1623.270 1304.340 ;
        RECT 1622.950 1290.540 1623.270 1290.600 ;
        RECT 1622.755 1290.400 1623.270 1290.540 ;
        RECT 1622.950 1290.340 1623.270 1290.400 ;
        RECT 1623.410 1159.300 1623.730 1159.360 ;
        RECT 1623.870 1159.300 1624.190 1159.360 ;
        RECT 1623.410 1159.160 1624.190 1159.300 ;
        RECT 1623.410 1159.100 1623.730 1159.160 ;
        RECT 1623.870 1159.100 1624.190 1159.160 ;
        RECT 1623.410 1062.740 1623.730 1062.800 ;
        RECT 1623.870 1062.740 1624.190 1062.800 ;
        RECT 1623.410 1062.600 1624.190 1062.740 ;
        RECT 1623.410 1062.540 1623.730 1062.600 ;
        RECT 1623.870 1062.540 1624.190 1062.600 ;
        RECT 1622.950 1007.320 1623.270 1007.380 ;
        RECT 1622.755 1007.180 1623.270 1007.320 ;
        RECT 1622.950 1007.120 1623.270 1007.180 ;
        RECT 1622.965 965.840 1623.255 965.885 ;
        RECT 1623.410 965.840 1623.730 965.900 ;
        RECT 1622.965 965.700 1623.730 965.840 ;
        RECT 1622.965 965.655 1623.255 965.700 ;
        RECT 1623.410 965.640 1623.730 965.700 ;
        RECT 1622.950 917.900 1623.270 917.960 ;
        RECT 1623.870 917.900 1624.190 917.960 ;
        RECT 1622.950 917.760 1624.190 917.900 ;
        RECT 1622.950 917.700 1623.270 917.760 ;
        RECT 1623.870 917.700 1624.190 917.760 ;
        RECT 1622.950 869.620 1623.270 869.680 ;
        RECT 1623.410 869.620 1623.730 869.680 ;
        RECT 1622.950 869.480 1623.730 869.620 ;
        RECT 1622.950 869.420 1623.270 869.480 ;
        RECT 1623.410 869.420 1623.730 869.480 ;
        RECT 1622.950 724.440 1623.270 724.500 ;
        RECT 1623.870 724.440 1624.190 724.500 ;
        RECT 1622.950 724.300 1624.190 724.440 ;
        RECT 1622.950 724.240 1623.270 724.300 ;
        RECT 1623.870 724.240 1624.190 724.300 ;
        RECT 1623.870 699.620 1624.190 699.680 ;
        RECT 1623.675 699.480 1624.190 699.620 ;
        RECT 1623.870 699.420 1624.190 699.480 ;
        RECT 1623.870 669.700 1624.190 669.760 ;
        RECT 1623.675 669.560 1624.190 669.700 ;
        RECT 1623.870 669.500 1624.190 669.560 ;
        RECT 1622.950 613.940 1623.270 614.000 ;
        RECT 1622.755 613.800 1623.270 613.940 ;
        RECT 1622.950 613.740 1623.270 613.800 ;
        RECT 1622.950 566.000 1623.270 566.060 ;
        RECT 1622.755 565.860 1623.270 566.000 ;
        RECT 1622.950 565.800 1623.270 565.860 ;
        RECT 1622.950 524.180 1623.270 524.240 ;
        RECT 1622.755 524.040 1623.270 524.180 ;
        RECT 1622.950 523.980 1623.270 524.040 ;
        RECT 1622.950 476.240 1623.270 476.300 ;
        RECT 1622.755 476.100 1623.270 476.240 ;
        RECT 1622.950 476.040 1623.270 476.100 ;
        RECT 1622.950 434.560 1623.270 434.820 ;
        RECT 1623.040 434.420 1623.180 434.560 ;
        RECT 1623.410 434.420 1623.730 434.480 ;
        RECT 1623.040 434.280 1623.730 434.420 ;
        RECT 1623.410 434.220 1623.730 434.280 ;
        RECT 1622.950 304.000 1623.270 304.260 ;
        RECT 1623.040 303.580 1623.180 304.000 ;
        RECT 1622.950 303.320 1623.270 303.580 ;
        RECT 1622.950 193.360 1623.270 193.420 ;
        RECT 1623.410 193.360 1623.730 193.420 ;
        RECT 1622.950 193.220 1623.730 193.360 ;
        RECT 1622.950 193.160 1623.270 193.220 ;
        RECT 1623.410 193.160 1623.730 193.220 ;
        RECT 1622.950 144.740 1623.270 144.800 ;
        RECT 1623.410 144.740 1623.730 144.800 ;
        RECT 1622.950 144.600 1623.730 144.740 ;
        RECT 1622.950 144.540 1623.270 144.600 ;
        RECT 1623.410 144.540 1623.730 144.600 ;
        RECT 1162.490 42.060 1162.810 42.120 ;
        RECT 1622.950 42.060 1623.270 42.120 ;
        RECT 1162.490 41.920 1623.270 42.060 ;
        RECT 1162.490 41.860 1162.810 41.920 ;
        RECT 1622.950 41.860 1623.270 41.920 ;
      LAYER via ;
        RECT 1623.440 1635.440 1623.700 1635.700 ;
        RECT 1625.280 1635.440 1625.540 1635.700 ;
        RECT 1623.440 1497.060 1623.700 1497.320 ;
        RECT 1623.440 1449.120 1623.700 1449.380 ;
        RECT 1622.520 1338.960 1622.780 1339.220 ;
        RECT 1623.440 1338.960 1623.700 1339.220 ;
        RECT 1622.980 1304.280 1623.240 1304.540 ;
        RECT 1622.980 1290.340 1623.240 1290.600 ;
        RECT 1623.440 1159.100 1623.700 1159.360 ;
        RECT 1623.900 1159.100 1624.160 1159.360 ;
        RECT 1623.440 1062.540 1623.700 1062.800 ;
        RECT 1623.900 1062.540 1624.160 1062.800 ;
        RECT 1622.980 1007.120 1623.240 1007.380 ;
        RECT 1623.440 965.640 1623.700 965.900 ;
        RECT 1622.980 917.700 1623.240 917.960 ;
        RECT 1623.900 917.700 1624.160 917.960 ;
        RECT 1622.980 869.420 1623.240 869.680 ;
        RECT 1623.440 869.420 1623.700 869.680 ;
        RECT 1622.980 724.240 1623.240 724.500 ;
        RECT 1623.900 724.240 1624.160 724.500 ;
        RECT 1623.900 699.420 1624.160 699.680 ;
        RECT 1623.900 669.500 1624.160 669.760 ;
        RECT 1622.980 613.740 1623.240 614.000 ;
        RECT 1622.980 565.800 1623.240 566.060 ;
        RECT 1622.980 523.980 1623.240 524.240 ;
        RECT 1622.980 476.040 1623.240 476.300 ;
        RECT 1622.980 434.560 1623.240 434.820 ;
        RECT 1623.440 434.220 1623.700 434.480 ;
        RECT 1622.980 304.000 1623.240 304.260 ;
        RECT 1622.980 303.320 1623.240 303.580 ;
        RECT 1622.980 193.160 1623.240 193.420 ;
        RECT 1623.440 193.160 1623.700 193.420 ;
        RECT 1622.980 144.540 1623.240 144.800 ;
        RECT 1623.440 144.540 1623.700 144.800 ;
        RECT 1162.520 41.860 1162.780 42.120 ;
        RECT 1622.980 41.860 1623.240 42.120 ;
      LAYER met2 ;
        RECT 1627.505 1701.090 1627.785 1704.000 ;
        RECT 1625.340 1700.950 1627.785 1701.090 ;
        RECT 1625.340 1635.730 1625.480 1700.950 ;
        RECT 1627.505 1700.000 1627.785 1700.950 ;
        RECT 1623.440 1635.410 1623.700 1635.730 ;
        RECT 1625.280 1635.410 1625.540 1635.730 ;
        RECT 1623.500 1559.650 1623.640 1635.410 ;
        RECT 1623.040 1559.510 1623.640 1559.650 ;
        RECT 1623.040 1510.690 1623.180 1559.510 ;
        RECT 1623.040 1510.550 1623.640 1510.690 ;
        RECT 1623.500 1497.350 1623.640 1510.550 ;
        RECT 1623.440 1497.030 1623.700 1497.350 ;
        RECT 1623.440 1449.090 1623.700 1449.410 ;
        RECT 1623.500 1426.370 1623.640 1449.090 ;
        RECT 1623.500 1426.230 1624.100 1426.370 ;
        RECT 1623.960 1387.045 1624.100 1426.230 ;
        RECT 1622.510 1386.675 1622.790 1387.045 ;
        RECT 1623.890 1386.675 1624.170 1387.045 ;
        RECT 1622.580 1339.250 1622.720 1386.675 ;
        RECT 1622.520 1338.930 1622.780 1339.250 ;
        RECT 1623.440 1338.930 1623.700 1339.250 ;
        RECT 1623.500 1338.650 1623.640 1338.930 ;
        RECT 1623.040 1338.510 1623.640 1338.650 ;
        RECT 1623.040 1304.570 1623.180 1338.510 ;
        RECT 1622.980 1304.250 1623.240 1304.570 ;
        RECT 1622.980 1290.310 1623.240 1290.630 ;
        RECT 1623.040 1193.925 1623.180 1290.310 ;
        RECT 1622.970 1193.555 1623.250 1193.925 ;
        RECT 1623.890 1193.555 1624.170 1193.925 ;
        RECT 1623.960 1159.390 1624.100 1193.555 ;
        RECT 1623.440 1159.245 1623.700 1159.390 ;
        RECT 1623.430 1158.875 1623.710 1159.245 ;
        RECT 1623.900 1159.070 1624.160 1159.390 ;
        RECT 1623.890 1158.195 1624.170 1158.565 ;
        RECT 1623.960 1062.830 1624.100 1158.195 ;
        RECT 1623.440 1062.570 1623.700 1062.830 ;
        RECT 1623.040 1062.510 1623.700 1062.570 ;
        RECT 1623.900 1062.510 1624.160 1062.830 ;
        RECT 1623.040 1062.430 1623.640 1062.510 ;
        RECT 1623.040 1007.410 1623.180 1062.430 ;
        RECT 1622.980 1007.090 1623.240 1007.410 ;
        RECT 1623.440 965.610 1623.700 965.930 ;
        RECT 1623.500 959.210 1623.640 965.610 ;
        RECT 1623.500 959.070 1624.100 959.210 ;
        RECT 1623.960 917.990 1624.100 959.070 ;
        RECT 1622.980 917.670 1623.240 917.990 ;
        RECT 1623.900 917.670 1624.160 917.990 ;
        RECT 1623.040 869.710 1623.180 917.670 ;
        RECT 1622.980 869.390 1623.240 869.710 ;
        RECT 1623.440 869.390 1623.700 869.710 ;
        RECT 1623.500 821.170 1623.640 869.390 ;
        RECT 1623.040 821.030 1623.640 821.170 ;
        RECT 1623.040 787.170 1623.180 821.030 ;
        RECT 1622.580 787.030 1623.180 787.170 ;
        RECT 1622.580 786.490 1622.720 787.030 ;
        RECT 1622.580 786.350 1623.180 786.490 ;
        RECT 1623.040 724.530 1623.180 786.350 ;
        RECT 1622.980 724.210 1623.240 724.530 ;
        RECT 1623.900 724.210 1624.160 724.530 ;
        RECT 1623.960 699.710 1624.100 724.210 ;
        RECT 1623.900 699.390 1624.160 699.710 ;
        RECT 1623.900 669.470 1624.160 669.790 ;
        RECT 1623.960 628.165 1624.100 669.470 ;
        RECT 1622.970 627.795 1623.250 628.165 ;
        RECT 1623.890 627.795 1624.170 628.165 ;
        RECT 1623.040 614.030 1623.180 627.795 ;
        RECT 1622.980 613.710 1623.240 614.030 ;
        RECT 1622.980 565.770 1623.240 566.090 ;
        RECT 1623.040 524.270 1623.180 565.770 ;
        RECT 1622.980 523.950 1623.240 524.270 ;
        RECT 1622.980 476.010 1623.240 476.330 ;
        RECT 1623.040 434.850 1623.180 476.010 ;
        RECT 1622.980 434.530 1623.240 434.850 ;
        RECT 1623.440 434.190 1623.700 434.510 ;
        RECT 1623.500 338.370 1623.640 434.190 ;
        RECT 1623.040 338.230 1623.640 338.370 ;
        RECT 1623.040 304.290 1623.180 338.230 ;
        RECT 1622.980 303.970 1623.240 304.290 ;
        RECT 1622.980 303.290 1623.240 303.610 ;
        RECT 1623.040 193.450 1623.180 303.290 ;
        RECT 1622.980 193.130 1623.240 193.450 ;
        RECT 1623.440 193.130 1623.700 193.450 ;
        RECT 1623.500 144.830 1623.640 193.130 ;
        RECT 1622.980 144.510 1623.240 144.830 ;
        RECT 1623.440 144.510 1623.700 144.830 ;
        RECT 1623.040 42.150 1623.180 144.510 ;
        RECT 1162.520 41.830 1162.780 42.150 ;
        RECT 1622.980 41.830 1623.240 42.150 ;
        RECT 1162.580 2.400 1162.720 41.830 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
      LAYER via2 ;
        RECT 1622.510 1386.720 1622.790 1387.000 ;
        RECT 1623.890 1386.720 1624.170 1387.000 ;
        RECT 1622.970 1193.600 1623.250 1193.880 ;
        RECT 1623.890 1193.600 1624.170 1193.880 ;
        RECT 1623.430 1158.920 1623.710 1159.200 ;
        RECT 1623.890 1158.240 1624.170 1158.520 ;
        RECT 1622.970 627.840 1623.250 628.120 ;
        RECT 1623.890 627.840 1624.170 628.120 ;
      LAYER met3 ;
        RECT 1622.485 1387.010 1622.815 1387.025 ;
        RECT 1623.865 1387.010 1624.195 1387.025 ;
        RECT 1622.485 1386.710 1624.195 1387.010 ;
        RECT 1622.485 1386.695 1622.815 1386.710 ;
        RECT 1623.865 1386.695 1624.195 1386.710 ;
        RECT 1622.945 1193.890 1623.275 1193.905 ;
        RECT 1623.865 1193.890 1624.195 1193.905 ;
        RECT 1622.945 1193.590 1624.195 1193.890 ;
        RECT 1622.945 1193.575 1623.275 1193.590 ;
        RECT 1623.865 1193.575 1624.195 1193.590 ;
        RECT 1623.405 1159.210 1623.735 1159.225 ;
        RECT 1623.190 1158.895 1623.735 1159.210 ;
        RECT 1623.190 1158.530 1623.490 1158.895 ;
        RECT 1623.865 1158.530 1624.195 1158.545 ;
        RECT 1623.190 1158.230 1624.195 1158.530 ;
        RECT 1623.865 1158.215 1624.195 1158.230 ;
        RECT 1622.945 628.130 1623.275 628.145 ;
        RECT 1623.865 628.130 1624.195 628.145 ;
        RECT 1622.945 627.830 1624.195 628.130 ;
        RECT 1622.945 627.815 1623.275 627.830 ;
        RECT 1623.865 627.815 1624.195 627.830 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 680.410 46.480 680.730 46.540 ;
        RECT 1429.290 46.480 1429.610 46.540 ;
        RECT 680.410 46.340 1429.610 46.480 ;
        RECT 680.410 46.280 680.730 46.340 ;
        RECT 1429.290 46.280 1429.610 46.340 ;
      LAYER via ;
        RECT 680.440 46.280 680.700 46.540 ;
        RECT 1429.320 46.280 1429.580 46.540 ;
      LAYER met2 ;
        RECT 1428.785 1700.410 1429.065 1704.000 ;
        RECT 1428.785 1700.270 1429.520 1700.410 ;
        RECT 1428.785 1700.000 1429.065 1700.270 ;
        RECT 1429.380 46.570 1429.520 1700.270 ;
        RECT 680.440 46.250 680.700 46.570 ;
        RECT 1429.320 46.250 1429.580 46.570 ;
        RECT 680.500 2.400 680.640 46.250 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1630.385 669.545 1630.555 688.755 ;
        RECT 1629.465 571.965 1629.635 613.955 ;
      LAYER mcon ;
        RECT 1630.385 688.585 1630.555 688.755 ;
        RECT 1629.465 613.785 1629.635 613.955 ;
      LAYER met1 ;
        RECT 1629.850 1635.640 1630.170 1635.700 ;
        RECT 1633.070 1635.640 1633.390 1635.700 ;
        RECT 1629.850 1635.500 1633.390 1635.640 ;
        RECT 1629.850 1635.440 1630.170 1635.500 ;
        RECT 1633.070 1635.440 1633.390 1635.500 ;
        RECT 1629.390 1497.060 1629.710 1497.320 ;
        RECT 1629.480 1496.920 1629.620 1497.060 ;
        RECT 1629.850 1496.920 1630.170 1496.980 ;
        RECT 1629.480 1496.780 1630.170 1496.920 ;
        RECT 1629.850 1496.720 1630.170 1496.780 ;
        RECT 1629.850 1435.040 1630.170 1435.100 ;
        RECT 1630.310 1435.040 1630.630 1435.100 ;
        RECT 1629.850 1434.900 1630.630 1435.040 ;
        RECT 1629.850 1434.840 1630.170 1434.900 ;
        RECT 1630.310 1434.840 1630.630 1434.900 ;
        RECT 1629.850 1338.820 1630.170 1338.880 ;
        RECT 1630.310 1338.820 1630.630 1338.880 ;
        RECT 1629.850 1338.680 1630.630 1338.820 ;
        RECT 1629.850 1338.620 1630.170 1338.680 ;
        RECT 1630.310 1338.620 1630.630 1338.680 ;
        RECT 1629.850 1159.300 1630.170 1159.360 ;
        RECT 1630.310 1159.300 1630.630 1159.360 ;
        RECT 1629.850 1159.160 1630.630 1159.300 ;
        RECT 1629.850 1159.100 1630.170 1159.160 ;
        RECT 1630.310 1159.100 1630.630 1159.160 ;
        RECT 1629.850 1111.360 1630.170 1111.420 ;
        RECT 1629.480 1111.220 1630.170 1111.360 ;
        RECT 1629.480 1111.080 1629.620 1111.220 ;
        RECT 1629.850 1111.160 1630.170 1111.220 ;
        RECT 1629.390 1110.820 1629.710 1111.080 ;
        RECT 1629.390 1062.740 1629.710 1062.800 ;
        RECT 1629.850 1062.740 1630.170 1062.800 ;
        RECT 1629.390 1062.600 1630.170 1062.740 ;
        RECT 1629.390 1062.540 1629.710 1062.600 ;
        RECT 1629.850 1062.540 1630.170 1062.600 ;
        RECT 1629.850 1014.800 1630.170 1014.860 ;
        RECT 1629.480 1014.660 1630.170 1014.800 ;
        RECT 1629.480 1014.520 1629.620 1014.660 ;
        RECT 1629.850 1014.600 1630.170 1014.660 ;
        RECT 1629.390 1014.260 1629.710 1014.520 ;
        RECT 1629.390 869.620 1629.710 869.680 ;
        RECT 1629.850 869.620 1630.170 869.680 ;
        RECT 1629.390 869.480 1630.170 869.620 ;
        RECT 1629.390 869.420 1629.710 869.480 ;
        RECT 1629.850 869.420 1630.170 869.480 ;
        RECT 1629.850 786.120 1630.170 786.380 ;
        RECT 1629.940 785.700 1630.080 786.120 ;
        RECT 1629.850 785.440 1630.170 785.700 ;
        RECT 1629.390 724.440 1629.710 724.500 ;
        RECT 1630.310 724.440 1630.630 724.500 ;
        RECT 1629.390 724.300 1630.630 724.440 ;
        RECT 1629.390 724.240 1629.710 724.300 ;
        RECT 1630.310 724.240 1630.630 724.300 ;
        RECT 1630.310 688.740 1630.630 688.800 ;
        RECT 1630.115 688.600 1630.630 688.740 ;
        RECT 1630.310 688.540 1630.630 688.600 ;
        RECT 1630.310 669.700 1630.630 669.760 ;
        RECT 1630.115 669.560 1630.630 669.700 ;
        RECT 1630.310 669.500 1630.630 669.560 ;
        RECT 1629.390 613.940 1629.710 614.000 ;
        RECT 1629.195 613.800 1629.710 613.940 ;
        RECT 1629.390 613.740 1629.710 613.800 ;
        RECT 1629.405 572.120 1629.695 572.165 ;
        RECT 1630.310 572.120 1630.630 572.180 ;
        RECT 1629.405 571.980 1630.630 572.120 ;
        RECT 1629.405 571.935 1629.695 571.980 ;
        RECT 1630.310 571.920 1630.630 571.980 ;
        RECT 1629.850 524.520 1630.170 524.580 ;
        RECT 1630.310 524.520 1630.630 524.580 ;
        RECT 1629.850 524.380 1630.630 524.520 ;
        RECT 1629.850 524.320 1630.170 524.380 ;
        RECT 1630.310 524.320 1630.630 524.380 ;
        RECT 1629.390 303.660 1629.710 303.920 ;
        RECT 1629.480 303.180 1629.620 303.660 ;
        RECT 1629.850 303.180 1630.170 303.240 ;
        RECT 1629.480 303.040 1630.170 303.180 ;
        RECT 1629.850 302.980 1630.170 303.040 ;
        RECT 1629.390 241.640 1629.710 241.700 ;
        RECT 1630.310 241.640 1630.630 241.700 ;
        RECT 1629.390 241.500 1630.630 241.640 ;
        RECT 1629.390 241.440 1629.710 241.500 ;
        RECT 1630.310 241.440 1630.630 241.500 ;
        RECT 1629.390 193.500 1629.710 193.760 ;
        RECT 1629.480 193.080 1629.620 193.500 ;
        RECT 1629.390 192.820 1629.710 193.080 ;
        RECT 1629.390 144.740 1629.710 144.800 ;
        RECT 1629.850 144.740 1630.170 144.800 ;
        RECT 1629.390 144.600 1630.170 144.740 ;
        RECT 1629.390 144.540 1629.710 144.600 ;
        RECT 1629.850 144.540 1630.170 144.600 ;
        RECT 1179.970 44.780 1180.290 44.840 ;
        RECT 1629.850 44.780 1630.170 44.840 ;
        RECT 1179.970 44.640 1630.170 44.780 ;
        RECT 1179.970 44.580 1180.290 44.640 ;
        RECT 1629.850 44.580 1630.170 44.640 ;
      LAYER via ;
        RECT 1629.880 1635.440 1630.140 1635.700 ;
        RECT 1633.100 1635.440 1633.360 1635.700 ;
        RECT 1629.420 1497.060 1629.680 1497.320 ;
        RECT 1629.880 1496.720 1630.140 1496.980 ;
        RECT 1629.880 1434.840 1630.140 1435.100 ;
        RECT 1630.340 1434.840 1630.600 1435.100 ;
        RECT 1629.880 1338.620 1630.140 1338.880 ;
        RECT 1630.340 1338.620 1630.600 1338.880 ;
        RECT 1629.880 1159.100 1630.140 1159.360 ;
        RECT 1630.340 1159.100 1630.600 1159.360 ;
        RECT 1629.880 1111.160 1630.140 1111.420 ;
        RECT 1629.420 1110.820 1629.680 1111.080 ;
        RECT 1629.420 1062.540 1629.680 1062.800 ;
        RECT 1629.880 1062.540 1630.140 1062.800 ;
        RECT 1629.880 1014.600 1630.140 1014.860 ;
        RECT 1629.420 1014.260 1629.680 1014.520 ;
        RECT 1629.420 869.420 1629.680 869.680 ;
        RECT 1629.880 869.420 1630.140 869.680 ;
        RECT 1629.880 786.120 1630.140 786.380 ;
        RECT 1629.880 785.440 1630.140 785.700 ;
        RECT 1629.420 724.240 1629.680 724.500 ;
        RECT 1630.340 724.240 1630.600 724.500 ;
        RECT 1630.340 688.540 1630.600 688.800 ;
        RECT 1630.340 669.500 1630.600 669.760 ;
        RECT 1629.420 613.740 1629.680 614.000 ;
        RECT 1630.340 571.920 1630.600 572.180 ;
        RECT 1629.880 524.320 1630.140 524.580 ;
        RECT 1630.340 524.320 1630.600 524.580 ;
        RECT 1629.420 303.660 1629.680 303.920 ;
        RECT 1629.880 302.980 1630.140 303.240 ;
        RECT 1629.420 241.440 1629.680 241.700 ;
        RECT 1630.340 241.440 1630.600 241.700 ;
        RECT 1629.420 193.500 1629.680 193.760 ;
        RECT 1629.420 192.820 1629.680 193.080 ;
        RECT 1629.420 144.540 1629.680 144.800 ;
        RECT 1629.880 144.540 1630.140 144.800 ;
        RECT 1180.000 44.580 1180.260 44.840 ;
        RECT 1629.880 44.580 1630.140 44.840 ;
      LAYER met2 ;
        RECT 1634.865 1700.410 1635.145 1704.000 ;
        RECT 1633.160 1700.270 1635.145 1700.410 ;
        RECT 1633.160 1635.730 1633.300 1700.270 ;
        RECT 1634.865 1700.000 1635.145 1700.270 ;
        RECT 1629.880 1635.410 1630.140 1635.730 ;
        RECT 1633.100 1635.410 1633.360 1635.730 ;
        RECT 1629.940 1511.370 1630.080 1635.410 ;
        RECT 1629.480 1511.230 1630.080 1511.370 ;
        RECT 1629.480 1497.350 1629.620 1511.230 ;
        RECT 1629.420 1497.030 1629.680 1497.350 ;
        RECT 1629.880 1496.690 1630.140 1497.010 ;
        RECT 1629.940 1435.130 1630.080 1496.690 ;
        RECT 1629.880 1434.810 1630.140 1435.130 ;
        RECT 1630.340 1434.810 1630.600 1435.130 ;
        RECT 1630.400 1338.910 1630.540 1434.810 ;
        RECT 1629.880 1338.590 1630.140 1338.910 ;
        RECT 1630.340 1338.590 1630.600 1338.910 ;
        RECT 1629.940 1314.850 1630.080 1338.590 ;
        RECT 1629.940 1314.710 1630.540 1314.850 ;
        RECT 1630.400 1159.390 1630.540 1314.710 ;
        RECT 1629.880 1159.070 1630.140 1159.390 ;
        RECT 1630.340 1159.070 1630.600 1159.390 ;
        RECT 1629.940 1111.450 1630.080 1159.070 ;
        RECT 1629.880 1111.130 1630.140 1111.450 ;
        RECT 1629.420 1110.790 1629.680 1111.110 ;
        RECT 1629.480 1062.830 1629.620 1110.790 ;
        RECT 1629.420 1062.510 1629.680 1062.830 ;
        RECT 1629.880 1062.510 1630.140 1062.830 ;
        RECT 1629.940 1014.890 1630.080 1062.510 ;
        RECT 1629.880 1014.570 1630.140 1014.890 ;
        RECT 1629.420 1014.405 1629.680 1014.550 ;
        RECT 1629.410 1014.035 1629.690 1014.405 ;
        RECT 1629.870 1013.355 1630.150 1013.725 ;
        RECT 1629.940 942.210 1630.080 1013.355 ;
        RECT 1629.480 942.070 1630.080 942.210 ;
        RECT 1629.480 869.710 1629.620 942.070 ;
        RECT 1629.420 869.390 1629.680 869.710 ;
        RECT 1629.880 869.390 1630.140 869.710 ;
        RECT 1629.940 821.170 1630.080 869.390 ;
        RECT 1629.480 821.030 1630.080 821.170 ;
        RECT 1629.480 789.890 1629.620 821.030 ;
        RECT 1629.480 789.750 1630.080 789.890 ;
        RECT 1629.940 786.410 1630.080 789.750 ;
        RECT 1629.880 786.090 1630.140 786.410 ;
        RECT 1629.880 785.410 1630.140 785.730 ;
        RECT 1629.940 749.090 1630.080 785.410 ;
        RECT 1629.940 748.950 1630.540 749.090 ;
        RECT 1630.400 724.725 1630.540 748.950 ;
        RECT 1629.410 724.355 1629.690 724.725 ;
        RECT 1630.330 724.355 1630.610 724.725 ;
        RECT 1629.420 724.210 1629.680 724.355 ;
        RECT 1630.340 724.210 1630.600 724.355 ;
        RECT 1630.400 688.830 1630.540 724.210 ;
        RECT 1630.340 688.510 1630.600 688.830 ;
        RECT 1630.340 669.470 1630.600 669.790 ;
        RECT 1630.400 628.165 1630.540 669.470 ;
        RECT 1629.410 627.795 1629.690 628.165 ;
        RECT 1630.330 627.795 1630.610 628.165 ;
        RECT 1629.480 614.030 1629.620 627.795 ;
        RECT 1629.420 613.710 1629.680 614.030 ;
        RECT 1630.340 571.890 1630.600 572.210 ;
        RECT 1630.400 524.610 1630.540 571.890 ;
        RECT 1629.880 524.290 1630.140 524.610 ;
        RECT 1630.340 524.290 1630.600 524.610 ;
        RECT 1629.940 338.370 1630.080 524.290 ;
        RECT 1629.480 338.230 1630.080 338.370 ;
        RECT 1629.480 303.950 1629.620 338.230 ;
        RECT 1629.420 303.630 1629.680 303.950 ;
        RECT 1629.880 302.950 1630.140 303.270 ;
        RECT 1629.940 266.290 1630.080 302.950 ;
        RECT 1629.940 266.150 1630.540 266.290 ;
        RECT 1630.400 241.730 1630.540 266.150 ;
        RECT 1629.420 241.410 1629.680 241.730 ;
        RECT 1630.340 241.410 1630.600 241.730 ;
        RECT 1629.480 193.790 1629.620 241.410 ;
        RECT 1629.420 193.470 1629.680 193.790 ;
        RECT 1629.420 192.790 1629.680 193.110 ;
        RECT 1629.480 144.830 1629.620 192.790 ;
        RECT 1629.420 144.510 1629.680 144.830 ;
        RECT 1629.880 144.510 1630.140 144.830 ;
        RECT 1629.940 44.870 1630.080 144.510 ;
        RECT 1180.000 44.550 1180.260 44.870 ;
        RECT 1629.880 44.550 1630.140 44.870 ;
        RECT 1180.060 2.400 1180.200 44.550 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
      LAYER via2 ;
        RECT 1629.410 1014.080 1629.690 1014.360 ;
        RECT 1629.870 1013.400 1630.150 1013.680 ;
        RECT 1629.410 724.400 1629.690 724.680 ;
        RECT 1630.330 724.400 1630.610 724.680 ;
        RECT 1629.410 627.840 1629.690 628.120 ;
        RECT 1630.330 627.840 1630.610 628.120 ;
      LAYER met3 ;
        RECT 1629.385 1014.370 1629.715 1014.385 ;
        RECT 1629.385 1014.055 1629.930 1014.370 ;
        RECT 1629.630 1013.705 1629.930 1014.055 ;
        RECT 1629.630 1013.390 1630.175 1013.705 ;
        RECT 1629.845 1013.375 1630.175 1013.390 ;
        RECT 1629.385 724.690 1629.715 724.705 ;
        RECT 1630.305 724.690 1630.635 724.705 ;
        RECT 1629.385 724.390 1630.635 724.690 ;
        RECT 1629.385 724.375 1629.715 724.390 ;
        RECT 1630.305 724.375 1630.635 724.390 ;
        RECT 1629.385 628.130 1629.715 628.145 ;
        RECT 1630.305 628.130 1630.635 628.145 ;
        RECT 1629.385 627.830 1630.635 628.130 ;
        RECT 1629.385 627.815 1629.715 627.830 ;
        RECT 1630.305 627.815 1630.635 627.830 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1197.910 45.120 1198.230 45.180 ;
        RECT 1643.190 45.120 1643.510 45.180 ;
        RECT 1197.910 44.980 1643.510 45.120 ;
        RECT 1197.910 44.920 1198.230 44.980 ;
        RECT 1643.190 44.920 1643.510 44.980 ;
      LAYER via ;
        RECT 1197.940 44.920 1198.200 45.180 ;
        RECT 1643.220 44.920 1643.480 45.180 ;
      LAYER met2 ;
        RECT 1642.225 1700.410 1642.505 1704.000 ;
        RECT 1642.225 1700.270 1643.420 1700.410 ;
        RECT 1642.225 1700.000 1642.505 1700.270 ;
        RECT 1643.280 45.210 1643.420 1700.270 ;
        RECT 1197.940 44.890 1198.200 45.210 ;
        RECT 1643.220 44.890 1643.480 45.210 ;
        RECT 1198.000 2.400 1198.140 44.890 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1650.090 1249.200 1650.410 1249.460 ;
        RECT 1650.180 1248.780 1650.320 1249.200 ;
        RECT 1650.090 1248.520 1650.410 1248.780 ;
        RECT 1650.090 386.620 1650.410 386.880 ;
        RECT 1650.180 386.200 1650.320 386.620 ;
        RECT 1650.090 385.940 1650.410 386.200 ;
        RECT 1215.850 45.460 1216.170 45.520 ;
        RECT 1650.090 45.460 1650.410 45.520 ;
        RECT 1215.850 45.320 1650.410 45.460 ;
        RECT 1215.850 45.260 1216.170 45.320 ;
        RECT 1650.090 45.260 1650.410 45.320 ;
      LAYER via ;
        RECT 1650.120 1249.200 1650.380 1249.460 ;
        RECT 1650.120 1248.520 1650.380 1248.780 ;
        RECT 1650.120 386.620 1650.380 386.880 ;
        RECT 1650.120 385.940 1650.380 386.200 ;
        RECT 1215.880 45.260 1216.140 45.520 ;
        RECT 1650.120 45.260 1650.380 45.520 ;
      LAYER met2 ;
        RECT 1649.585 1700.410 1649.865 1704.000 ;
        RECT 1649.585 1700.270 1650.320 1700.410 ;
        RECT 1649.585 1700.000 1649.865 1700.270 ;
        RECT 1650.180 1249.490 1650.320 1700.270 ;
        RECT 1650.120 1249.170 1650.380 1249.490 ;
        RECT 1650.120 1248.490 1650.380 1248.810 ;
        RECT 1650.180 386.910 1650.320 1248.490 ;
        RECT 1650.120 386.590 1650.380 386.910 ;
        RECT 1650.120 385.910 1650.380 386.230 ;
        RECT 1650.180 45.550 1650.320 385.910 ;
        RECT 1215.880 45.230 1216.140 45.550 ;
        RECT 1650.120 45.230 1650.380 45.550 ;
        RECT 1215.940 2.400 1216.080 45.230 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1657.065 1594.345 1657.235 1659.455 ;
        RECT 1657.065 1497.785 1657.235 1587.035 ;
        RECT 1657.065 1338.665 1657.235 1386.775 ;
        RECT 1657.065 1183.285 1657.235 1297.015 ;
        RECT 1657.065 1104.065 1657.235 1111.035 ;
        RECT 1657.065 958.885 1657.235 1000.535 ;
        RECT 1657.985 807.245 1658.155 855.355 ;
        RECT 1657.065 669.545 1657.235 730.235 ;
        RECT 1657.065 469.285 1657.235 517.395 ;
        RECT 1657.065 48.365 1657.235 131.155 ;
      LAYER mcon ;
        RECT 1657.065 1659.285 1657.235 1659.455 ;
        RECT 1657.065 1586.865 1657.235 1587.035 ;
        RECT 1657.065 1386.605 1657.235 1386.775 ;
        RECT 1657.065 1296.845 1657.235 1297.015 ;
        RECT 1657.065 1110.865 1657.235 1111.035 ;
        RECT 1657.065 1000.365 1657.235 1000.535 ;
        RECT 1657.985 855.185 1658.155 855.355 ;
        RECT 1657.065 730.065 1657.235 730.235 ;
        RECT 1657.065 517.225 1657.235 517.395 ;
        RECT 1657.065 130.985 1657.235 131.155 ;
      LAYER met1 ;
        RECT 1656.990 1659.440 1657.310 1659.500 ;
        RECT 1656.795 1659.300 1657.310 1659.440 ;
        RECT 1656.990 1659.240 1657.310 1659.300 ;
        RECT 1656.990 1594.500 1657.310 1594.560 ;
        RECT 1656.795 1594.360 1657.310 1594.500 ;
        RECT 1656.990 1594.300 1657.310 1594.360 ;
        RECT 1656.990 1587.020 1657.310 1587.080 ;
        RECT 1656.795 1586.880 1657.310 1587.020 ;
        RECT 1656.990 1586.820 1657.310 1586.880 ;
        RECT 1656.990 1497.940 1657.310 1498.000 ;
        RECT 1656.795 1497.800 1657.310 1497.940 ;
        RECT 1656.990 1497.740 1657.310 1497.800 ;
        RECT 1656.990 1442.180 1657.310 1442.240 ;
        RECT 1657.450 1442.180 1657.770 1442.240 ;
        RECT 1656.990 1442.040 1657.770 1442.180 ;
        RECT 1656.990 1441.980 1657.310 1442.040 ;
        RECT 1657.450 1441.980 1657.770 1442.040 ;
        RECT 1657.450 1394.240 1657.770 1394.300 ;
        RECT 1657.080 1394.100 1657.770 1394.240 ;
        RECT 1657.080 1393.620 1657.220 1394.100 ;
        RECT 1657.450 1394.040 1657.770 1394.100 ;
        RECT 1656.990 1393.360 1657.310 1393.620 ;
        RECT 1656.990 1386.760 1657.310 1386.820 ;
        RECT 1656.795 1386.620 1657.310 1386.760 ;
        RECT 1656.990 1386.560 1657.310 1386.620 ;
        RECT 1656.990 1338.820 1657.310 1338.880 ;
        RECT 1656.795 1338.680 1657.310 1338.820 ;
        RECT 1656.990 1338.620 1657.310 1338.680 ;
        RECT 1656.990 1297.000 1657.310 1297.060 ;
        RECT 1656.795 1296.860 1657.310 1297.000 ;
        RECT 1656.990 1296.800 1657.310 1296.860 ;
        RECT 1656.990 1183.440 1657.310 1183.500 ;
        RECT 1656.795 1183.300 1657.310 1183.440 ;
        RECT 1656.990 1183.240 1657.310 1183.300 ;
        RECT 1656.990 1111.020 1657.310 1111.080 ;
        RECT 1656.795 1110.880 1657.310 1111.020 ;
        RECT 1656.990 1110.820 1657.310 1110.880 ;
        RECT 1656.990 1104.220 1657.310 1104.280 ;
        RECT 1656.795 1104.080 1657.310 1104.220 ;
        RECT 1656.990 1104.020 1657.310 1104.080 ;
        RECT 1656.990 1014.940 1657.310 1015.200 ;
        RECT 1657.080 1014.520 1657.220 1014.940 ;
        RECT 1656.990 1014.260 1657.310 1014.520 ;
        RECT 1656.990 1000.520 1657.310 1000.580 ;
        RECT 1656.795 1000.380 1657.310 1000.520 ;
        RECT 1656.990 1000.320 1657.310 1000.380 ;
        RECT 1657.005 959.040 1657.295 959.085 ;
        RECT 1657.910 959.040 1658.230 959.100 ;
        RECT 1657.005 958.900 1658.230 959.040 ;
        RECT 1657.005 958.855 1657.295 958.900 ;
        RECT 1657.910 958.840 1658.230 958.900 ;
        RECT 1656.990 952.240 1657.310 952.300 ;
        RECT 1658.370 952.240 1658.690 952.300 ;
        RECT 1656.990 952.100 1658.690 952.240 ;
        RECT 1656.990 952.040 1657.310 952.100 ;
        RECT 1658.370 952.040 1658.690 952.100 ;
        RECT 1657.910 862.620 1658.230 862.880 ;
        RECT 1658.000 862.200 1658.140 862.620 ;
        RECT 1657.910 861.940 1658.230 862.200 ;
        RECT 1657.910 855.340 1658.230 855.400 ;
        RECT 1657.715 855.200 1658.230 855.340 ;
        RECT 1657.910 855.140 1658.230 855.200 ;
        RECT 1657.925 807.400 1658.215 807.445 ;
        RECT 1658.370 807.400 1658.690 807.460 ;
        RECT 1657.925 807.260 1658.690 807.400 ;
        RECT 1657.925 807.215 1658.215 807.260 ;
        RECT 1658.370 807.200 1658.690 807.260 ;
        RECT 1656.990 730.220 1657.310 730.280 ;
        RECT 1656.795 730.080 1657.310 730.220 ;
        RECT 1656.990 730.020 1657.310 730.080 ;
        RECT 1656.990 669.700 1657.310 669.760 ;
        RECT 1656.795 669.560 1657.310 669.700 ;
        RECT 1656.990 669.500 1657.310 669.560 ;
        RECT 1656.990 627.880 1657.310 627.940 ;
        RECT 1657.910 627.880 1658.230 627.940 ;
        RECT 1656.990 627.740 1658.230 627.880 ;
        RECT 1656.990 627.680 1657.310 627.740 ;
        RECT 1657.910 627.680 1658.230 627.740 ;
        RECT 1656.990 517.380 1657.310 517.440 ;
        RECT 1656.795 517.240 1657.310 517.380 ;
        RECT 1656.990 517.180 1657.310 517.240 ;
        RECT 1656.990 469.440 1657.310 469.500 ;
        RECT 1656.795 469.300 1657.310 469.440 ;
        RECT 1656.990 469.240 1657.310 469.300 ;
        RECT 1656.990 427.960 1657.310 428.020 ;
        RECT 1658.370 427.960 1658.690 428.020 ;
        RECT 1656.990 427.820 1658.690 427.960 ;
        RECT 1656.990 427.760 1657.310 427.820 ;
        RECT 1658.370 427.760 1658.690 427.820 ;
        RECT 1656.990 379.680 1657.310 379.740 ;
        RECT 1658.370 379.680 1658.690 379.740 ;
        RECT 1656.990 379.540 1658.690 379.680 ;
        RECT 1656.990 379.480 1657.310 379.540 ;
        RECT 1658.370 379.480 1658.690 379.540 ;
        RECT 1655.610 193.360 1655.930 193.420 ;
        RECT 1657.450 193.360 1657.770 193.420 ;
        RECT 1655.610 193.220 1657.770 193.360 ;
        RECT 1655.610 193.160 1655.930 193.220 ;
        RECT 1657.450 193.160 1657.770 193.220 ;
        RECT 1656.990 131.140 1657.310 131.200 ;
        RECT 1656.795 131.000 1657.310 131.140 ;
        RECT 1656.990 130.940 1657.310 131.000 ;
        RECT 1656.990 48.520 1657.310 48.580 ;
        RECT 1656.795 48.380 1657.310 48.520 ;
        RECT 1656.990 48.320 1657.310 48.380 ;
        RECT 1233.790 41.720 1234.110 41.780 ;
        RECT 1656.990 41.720 1657.310 41.780 ;
        RECT 1233.790 41.580 1657.310 41.720 ;
        RECT 1233.790 41.520 1234.110 41.580 ;
        RECT 1656.990 41.520 1657.310 41.580 ;
      LAYER via ;
        RECT 1657.020 1659.240 1657.280 1659.500 ;
        RECT 1657.020 1594.300 1657.280 1594.560 ;
        RECT 1657.020 1586.820 1657.280 1587.080 ;
        RECT 1657.020 1497.740 1657.280 1498.000 ;
        RECT 1657.020 1441.980 1657.280 1442.240 ;
        RECT 1657.480 1441.980 1657.740 1442.240 ;
        RECT 1657.480 1394.040 1657.740 1394.300 ;
        RECT 1657.020 1393.360 1657.280 1393.620 ;
        RECT 1657.020 1386.560 1657.280 1386.820 ;
        RECT 1657.020 1338.620 1657.280 1338.880 ;
        RECT 1657.020 1296.800 1657.280 1297.060 ;
        RECT 1657.020 1183.240 1657.280 1183.500 ;
        RECT 1657.020 1110.820 1657.280 1111.080 ;
        RECT 1657.020 1104.020 1657.280 1104.280 ;
        RECT 1657.020 1014.940 1657.280 1015.200 ;
        RECT 1657.020 1014.260 1657.280 1014.520 ;
        RECT 1657.020 1000.320 1657.280 1000.580 ;
        RECT 1657.940 958.840 1658.200 959.100 ;
        RECT 1657.020 952.040 1657.280 952.300 ;
        RECT 1658.400 952.040 1658.660 952.300 ;
        RECT 1657.940 862.620 1658.200 862.880 ;
        RECT 1657.940 861.940 1658.200 862.200 ;
        RECT 1657.940 855.140 1658.200 855.400 ;
        RECT 1658.400 807.200 1658.660 807.460 ;
        RECT 1657.020 730.020 1657.280 730.280 ;
        RECT 1657.020 669.500 1657.280 669.760 ;
        RECT 1657.020 627.680 1657.280 627.940 ;
        RECT 1657.940 627.680 1658.200 627.940 ;
        RECT 1657.020 517.180 1657.280 517.440 ;
        RECT 1657.020 469.240 1657.280 469.500 ;
        RECT 1657.020 427.760 1657.280 428.020 ;
        RECT 1658.400 427.760 1658.660 428.020 ;
        RECT 1657.020 379.480 1657.280 379.740 ;
        RECT 1658.400 379.480 1658.660 379.740 ;
        RECT 1655.640 193.160 1655.900 193.420 ;
        RECT 1657.480 193.160 1657.740 193.420 ;
        RECT 1657.020 130.940 1657.280 131.200 ;
        RECT 1657.020 48.320 1657.280 48.580 ;
        RECT 1233.820 41.520 1234.080 41.780 ;
        RECT 1657.020 41.520 1657.280 41.780 ;
      LAYER met2 ;
        RECT 1656.945 1700.000 1657.225 1704.000 ;
        RECT 1657.080 1659.530 1657.220 1700.000 ;
        RECT 1657.020 1659.210 1657.280 1659.530 ;
        RECT 1657.020 1594.270 1657.280 1594.590 ;
        RECT 1657.080 1587.110 1657.220 1594.270 ;
        RECT 1657.020 1586.790 1657.280 1587.110 ;
        RECT 1657.020 1497.710 1657.280 1498.030 ;
        RECT 1657.080 1442.270 1657.220 1497.710 ;
        RECT 1657.020 1441.950 1657.280 1442.270 ;
        RECT 1657.480 1441.950 1657.740 1442.270 ;
        RECT 1657.540 1394.330 1657.680 1441.950 ;
        RECT 1657.480 1394.010 1657.740 1394.330 ;
        RECT 1657.020 1393.330 1657.280 1393.650 ;
        RECT 1657.080 1386.850 1657.220 1393.330 ;
        RECT 1657.020 1386.530 1657.280 1386.850 ;
        RECT 1657.020 1338.590 1657.280 1338.910 ;
        RECT 1657.080 1297.090 1657.220 1338.590 ;
        RECT 1657.020 1296.770 1657.280 1297.090 ;
        RECT 1657.020 1183.210 1657.280 1183.530 ;
        RECT 1657.080 1111.110 1657.220 1183.210 ;
        RECT 1657.020 1110.790 1657.280 1111.110 ;
        RECT 1657.080 1104.310 1657.220 1104.465 ;
        RECT 1657.020 1104.050 1657.280 1104.310 ;
        RECT 1657.020 1103.990 1657.680 1104.050 ;
        RECT 1657.080 1103.910 1657.680 1103.990 ;
        RECT 1657.540 1055.770 1657.680 1103.910 ;
        RECT 1657.080 1055.630 1657.680 1055.770 ;
        RECT 1657.080 1015.230 1657.220 1055.630 ;
        RECT 1657.020 1014.910 1657.280 1015.230 ;
        RECT 1657.020 1014.230 1657.280 1014.550 ;
        RECT 1657.080 1000.610 1657.220 1014.230 ;
        RECT 1657.020 1000.290 1657.280 1000.610 ;
        RECT 1657.940 958.810 1658.200 959.130 ;
        RECT 1658.000 952.410 1658.140 958.810 ;
        RECT 1658.000 952.330 1658.600 952.410 ;
        RECT 1657.020 952.010 1657.280 952.330 ;
        RECT 1658.000 952.270 1658.660 952.330 ;
        RECT 1658.400 952.010 1658.660 952.270 ;
        RECT 1657.080 904.245 1657.220 952.010 ;
        RECT 1658.460 951.855 1658.600 952.010 ;
        RECT 1657.010 903.875 1657.290 904.245 ;
        RECT 1657.930 903.875 1658.210 904.245 ;
        RECT 1658.000 862.910 1658.140 903.875 ;
        RECT 1657.940 862.590 1658.200 862.910 ;
        RECT 1657.940 861.910 1658.200 862.230 ;
        RECT 1658.000 855.430 1658.140 861.910 ;
        RECT 1657.940 855.110 1658.200 855.430 ;
        RECT 1658.400 807.170 1658.660 807.490 ;
        RECT 1658.460 759.405 1658.600 807.170 ;
        RECT 1657.470 759.290 1657.750 759.405 ;
        RECT 1657.080 759.150 1657.750 759.290 ;
        RECT 1657.080 730.310 1657.220 759.150 ;
        RECT 1657.470 759.035 1657.750 759.150 ;
        RECT 1658.390 759.035 1658.670 759.405 ;
        RECT 1657.020 729.990 1657.280 730.310 ;
        RECT 1657.020 669.470 1657.280 669.790 ;
        RECT 1657.080 627.970 1657.220 669.470 ;
        RECT 1657.020 627.650 1657.280 627.970 ;
        RECT 1657.940 627.650 1658.200 627.970 ;
        RECT 1658.000 592.010 1658.140 627.650 ;
        RECT 1657.540 591.870 1658.140 592.010 ;
        RECT 1657.540 524.690 1657.680 591.870 ;
        RECT 1657.080 524.550 1657.680 524.690 ;
        RECT 1657.080 517.470 1657.220 524.550 ;
        RECT 1657.020 517.150 1657.280 517.470 ;
        RECT 1657.020 469.210 1657.280 469.530 ;
        RECT 1657.080 428.050 1657.220 469.210 ;
        RECT 1657.020 427.730 1657.280 428.050 ;
        RECT 1658.400 427.730 1658.660 428.050 ;
        RECT 1658.460 379.770 1658.600 427.730 ;
        RECT 1657.020 379.450 1657.280 379.770 ;
        RECT 1658.400 379.450 1658.660 379.770 ;
        RECT 1657.080 331.005 1657.220 379.450 ;
        RECT 1657.010 330.635 1657.290 331.005 ;
        RECT 1657.930 329.955 1658.210 330.325 ;
        RECT 1658.000 241.925 1658.140 329.955 ;
        RECT 1657.930 241.555 1658.210 241.925 ;
        RECT 1655.630 240.875 1655.910 241.245 ;
        RECT 1655.700 193.450 1655.840 240.875 ;
        RECT 1655.640 193.130 1655.900 193.450 ;
        RECT 1657.480 193.130 1657.740 193.450 ;
        RECT 1657.540 139.245 1657.680 193.130 ;
        RECT 1657.470 138.875 1657.750 139.245 ;
        RECT 1657.010 138.195 1657.290 138.565 ;
        RECT 1657.080 131.230 1657.220 138.195 ;
        RECT 1657.020 130.910 1657.280 131.230 ;
        RECT 1657.020 48.290 1657.280 48.610 ;
        RECT 1657.080 41.810 1657.220 48.290 ;
        RECT 1233.820 41.490 1234.080 41.810 ;
        RECT 1657.020 41.490 1657.280 41.810 ;
        RECT 1233.880 2.400 1234.020 41.490 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
      LAYER via2 ;
        RECT 1657.010 903.920 1657.290 904.200 ;
        RECT 1657.930 903.920 1658.210 904.200 ;
        RECT 1657.470 759.080 1657.750 759.360 ;
        RECT 1658.390 759.080 1658.670 759.360 ;
        RECT 1657.010 330.680 1657.290 330.960 ;
        RECT 1657.930 330.000 1658.210 330.280 ;
        RECT 1657.930 241.600 1658.210 241.880 ;
        RECT 1655.630 240.920 1655.910 241.200 ;
        RECT 1657.470 138.920 1657.750 139.200 ;
        RECT 1657.010 138.240 1657.290 138.520 ;
      LAYER met3 ;
        RECT 1656.985 904.210 1657.315 904.225 ;
        RECT 1657.905 904.210 1658.235 904.225 ;
        RECT 1656.985 903.910 1658.235 904.210 ;
        RECT 1656.985 903.895 1657.315 903.910 ;
        RECT 1657.905 903.895 1658.235 903.910 ;
        RECT 1657.445 759.370 1657.775 759.385 ;
        RECT 1658.365 759.370 1658.695 759.385 ;
        RECT 1657.445 759.070 1658.695 759.370 ;
        RECT 1657.445 759.055 1657.775 759.070 ;
        RECT 1658.365 759.055 1658.695 759.070 ;
        RECT 1656.985 330.970 1657.315 330.985 ;
        RECT 1656.310 330.670 1657.315 330.970 ;
        RECT 1656.310 330.290 1656.610 330.670 ;
        RECT 1656.985 330.655 1657.315 330.670 ;
        RECT 1657.905 330.290 1658.235 330.305 ;
        RECT 1656.310 329.990 1658.235 330.290 ;
        RECT 1657.905 329.975 1658.235 329.990 ;
        RECT 1657.905 241.890 1658.235 241.905 ;
        RECT 1656.310 241.590 1658.235 241.890 ;
        RECT 1655.605 241.210 1655.935 241.225 ;
        RECT 1656.310 241.210 1656.610 241.590 ;
        RECT 1657.905 241.575 1658.235 241.590 ;
        RECT 1655.605 240.910 1656.610 241.210 ;
        RECT 1655.605 240.895 1655.935 240.910 ;
        RECT 1657.445 139.210 1657.775 139.225 ;
        RECT 1656.310 138.910 1657.775 139.210 ;
        RECT 1656.310 138.530 1656.610 138.910 ;
        RECT 1657.445 138.895 1657.775 138.910 ;
        RECT 1656.985 138.530 1657.315 138.545 ;
        RECT 1656.310 138.230 1657.315 138.530 ;
        RECT 1656.985 138.215 1657.315 138.230 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1251.730 45.800 1252.050 45.860 ;
        RECT 1663.890 45.800 1664.210 45.860 ;
        RECT 1251.730 45.660 1664.210 45.800 ;
        RECT 1251.730 45.600 1252.050 45.660 ;
        RECT 1663.890 45.600 1664.210 45.660 ;
      LAYER via ;
        RECT 1251.760 45.600 1252.020 45.860 ;
        RECT 1663.920 45.600 1664.180 45.860 ;
      LAYER met2 ;
        RECT 1664.305 1700.410 1664.585 1704.000 ;
        RECT 1663.980 1700.270 1664.585 1700.410 ;
        RECT 1663.980 45.890 1664.120 1700.270 ;
        RECT 1664.305 1700.000 1664.585 1700.270 ;
        RECT 1251.760 45.570 1252.020 45.890 ;
        RECT 1663.920 45.570 1664.180 45.890 ;
        RECT 1251.820 2.400 1251.960 45.570 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1269.210 46.140 1269.530 46.200 ;
        RECT 1670.790 46.140 1671.110 46.200 ;
        RECT 1269.210 46.000 1671.110 46.140 ;
        RECT 1269.210 45.940 1269.530 46.000 ;
        RECT 1670.790 45.940 1671.110 46.000 ;
      LAYER via ;
        RECT 1269.240 45.940 1269.500 46.200 ;
        RECT 1670.820 45.940 1671.080 46.200 ;
      LAYER met2 ;
        RECT 1671.665 1700.410 1671.945 1704.000 ;
        RECT 1670.880 1700.270 1671.945 1700.410 ;
        RECT 1670.880 46.230 1671.020 1700.270 ;
        RECT 1671.665 1700.000 1671.945 1700.270 ;
        RECT 1269.240 45.910 1269.500 46.230 ;
        RECT 1670.820 45.910 1671.080 46.230 ;
        RECT 1269.300 2.400 1269.440 45.910 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1438.105 19.805 1438.275 20.995 ;
      LAYER mcon ;
        RECT 1438.105 20.825 1438.275 20.995 ;
      LAYER met1 ;
        RECT 1479.430 33.220 1479.750 33.280 ;
        RECT 1677.230 33.220 1677.550 33.280 ;
        RECT 1479.430 33.080 1677.550 33.220 ;
        RECT 1479.430 33.020 1479.750 33.080 ;
        RECT 1677.230 33.020 1677.550 33.080 ;
        RECT 1438.045 20.980 1438.335 21.025 ;
        RECT 1438.045 20.840 1439.640 20.980 ;
        RECT 1438.045 20.795 1438.335 20.840 ;
        RECT 1439.500 20.640 1439.640 20.840 ;
        RECT 1479.430 20.640 1479.750 20.700 ;
        RECT 1439.500 20.500 1479.750 20.640 ;
        RECT 1479.430 20.440 1479.750 20.500 ;
        RECT 1287.150 19.960 1287.470 20.020 ;
        RECT 1438.045 19.960 1438.335 20.005 ;
        RECT 1287.150 19.820 1438.335 19.960 ;
        RECT 1287.150 19.760 1287.470 19.820 ;
        RECT 1438.045 19.775 1438.335 19.820 ;
      LAYER via ;
        RECT 1479.460 33.020 1479.720 33.280 ;
        RECT 1677.260 33.020 1677.520 33.280 ;
        RECT 1479.460 20.440 1479.720 20.700 ;
        RECT 1287.180 19.760 1287.440 20.020 ;
      LAYER met2 ;
        RECT 1679.025 1700.410 1679.305 1704.000 ;
        RECT 1677.320 1700.270 1679.305 1700.410 ;
        RECT 1677.320 33.310 1677.460 1700.270 ;
        RECT 1679.025 1700.000 1679.305 1700.270 ;
        RECT 1479.460 32.990 1479.720 33.310 ;
        RECT 1677.260 32.990 1677.520 33.310 ;
        RECT 1479.520 20.730 1479.660 32.990 ;
        RECT 1479.460 20.410 1479.720 20.730 ;
        RECT 1287.180 19.730 1287.440 20.050 ;
        RECT 1287.240 2.400 1287.380 19.730 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1323.105 5.525 1323.275 20.315 ;
        RECT 1345.645 20.145 1345.815 21.335 ;
        RECT 1393.485 20.145 1393.655 21.335 ;
        RECT 1414.645 18.445 1414.815 20.315 ;
        RECT 1438.565 18.445 1438.735 19.975 ;
      LAYER mcon ;
        RECT 1345.645 21.165 1345.815 21.335 ;
        RECT 1323.105 20.145 1323.275 20.315 ;
        RECT 1393.485 21.165 1393.655 21.335 ;
        RECT 1414.645 20.145 1414.815 20.315 ;
        RECT 1438.565 19.805 1438.735 19.975 ;
      LAYER met1 ;
        RECT 1685.050 1635.980 1685.370 1636.040 ;
        RECT 1684.220 1635.840 1685.370 1635.980 ;
        RECT 1684.220 1635.700 1684.360 1635.840 ;
        RECT 1685.050 1635.780 1685.370 1635.840 ;
        RECT 1684.130 1635.440 1684.450 1635.700 ;
        RECT 1486.790 33.560 1487.110 33.620 ;
        RECT 1684.130 33.560 1684.450 33.620 ;
        RECT 1486.790 33.420 1684.450 33.560 ;
        RECT 1486.790 33.360 1487.110 33.420 ;
        RECT 1684.130 33.360 1684.450 33.420 ;
        RECT 1345.585 21.320 1345.875 21.365 ;
        RECT 1393.425 21.320 1393.715 21.365 ;
        RECT 1345.585 21.180 1393.715 21.320 ;
        RECT 1345.585 21.135 1345.875 21.180 ;
        RECT 1393.425 21.135 1393.715 21.180 ;
        RECT 1323.045 20.300 1323.335 20.345 ;
        RECT 1345.585 20.300 1345.875 20.345 ;
        RECT 1323.045 20.160 1345.875 20.300 ;
        RECT 1323.045 20.115 1323.335 20.160 ;
        RECT 1345.585 20.115 1345.875 20.160 ;
        RECT 1393.425 20.300 1393.715 20.345 ;
        RECT 1414.585 20.300 1414.875 20.345 ;
        RECT 1393.425 20.160 1414.875 20.300 ;
        RECT 1393.425 20.115 1393.715 20.160 ;
        RECT 1414.585 20.115 1414.875 20.160 ;
        RECT 1438.505 19.960 1438.795 20.005 ;
        RECT 1486.790 19.960 1487.110 20.020 ;
        RECT 1438.505 19.820 1487.110 19.960 ;
        RECT 1438.505 19.775 1438.795 19.820 ;
        RECT 1486.790 19.760 1487.110 19.820 ;
        RECT 1414.585 18.600 1414.875 18.645 ;
        RECT 1438.505 18.600 1438.795 18.645 ;
        RECT 1414.585 18.460 1438.795 18.600 ;
        RECT 1414.585 18.415 1414.875 18.460 ;
        RECT 1438.505 18.415 1438.795 18.460 ;
        RECT 1305.090 5.680 1305.410 5.740 ;
        RECT 1323.045 5.680 1323.335 5.725 ;
        RECT 1305.090 5.540 1323.335 5.680 ;
        RECT 1305.090 5.480 1305.410 5.540 ;
        RECT 1323.045 5.495 1323.335 5.540 ;
      LAYER via ;
        RECT 1685.080 1635.780 1685.340 1636.040 ;
        RECT 1684.160 1635.440 1684.420 1635.700 ;
        RECT 1486.820 33.360 1487.080 33.620 ;
        RECT 1684.160 33.360 1684.420 33.620 ;
        RECT 1486.820 19.760 1487.080 20.020 ;
        RECT 1305.120 5.480 1305.380 5.740 ;
      LAYER met2 ;
        RECT 1686.385 1700.410 1686.665 1704.000 ;
        RECT 1685.140 1700.270 1686.665 1700.410 ;
        RECT 1685.140 1636.070 1685.280 1700.270 ;
        RECT 1686.385 1700.000 1686.665 1700.270 ;
        RECT 1685.080 1635.750 1685.340 1636.070 ;
        RECT 1684.160 1635.410 1684.420 1635.730 ;
        RECT 1684.220 33.650 1684.360 1635.410 ;
        RECT 1486.820 33.330 1487.080 33.650 ;
        RECT 1684.160 33.330 1684.420 33.650 ;
        RECT 1486.880 20.050 1487.020 33.330 ;
        RECT 1486.820 19.730 1487.080 20.050 ;
        RECT 1305.120 5.450 1305.380 5.770 ;
        RECT 1305.180 2.400 1305.320 5.450 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1367.265 19.125 1367.435 20.655 ;
      LAYER mcon ;
        RECT 1367.265 20.485 1367.435 20.655 ;
      LAYER met1 ;
        RECT 1490.470 32.880 1490.790 32.940 ;
        RECT 1691.950 32.880 1692.270 32.940 ;
        RECT 1490.470 32.740 1692.270 32.880 ;
        RECT 1490.470 32.680 1490.790 32.740 ;
        RECT 1691.950 32.680 1692.270 32.740 ;
        RECT 1423.400 20.840 1428.600 20.980 ;
        RECT 1367.205 20.640 1367.495 20.685 ;
        RECT 1423.400 20.640 1423.540 20.840 ;
        RECT 1367.205 20.500 1423.540 20.640 ;
        RECT 1428.460 20.640 1428.600 20.840 ;
        RECT 1428.460 20.500 1439.180 20.640 ;
        RECT 1367.205 20.455 1367.495 20.500 ;
        RECT 1439.040 20.300 1439.180 20.500 ;
        RECT 1490.470 20.300 1490.790 20.360 ;
        RECT 1439.040 20.160 1490.790 20.300 ;
        RECT 1490.470 20.100 1490.790 20.160 ;
        RECT 1323.030 19.280 1323.350 19.340 ;
        RECT 1367.205 19.280 1367.495 19.325 ;
        RECT 1323.030 19.140 1367.495 19.280 ;
        RECT 1323.030 19.080 1323.350 19.140 ;
        RECT 1367.205 19.095 1367.495 19.140 ;
      LAYER via ;
        RECT 1490.500 32.680 1490.760 32.940 ;
        RECT 1691.980 32.680 1692.240 32.940 ;
        RECT 1490.500 20.100 1490.760 20.360 ;
        RECT 1323.060 19.080 1323.320 19.340 ;
      LAYER met2 ;
        RECT 1693.745 1700.410 1694.025 1704.000 ;
        RECT 1692.040 1700.270 1694.025 1700.410 ;
        RECT 1692.040 32.970 1692.180 1700.270 ;
        RECT 1693.745 1700.000 1694.025 1700.270 ;
        RECT 1490.500 32.650 1490.760 32.970 ;
        RECT 1691.980 32.650 1692.240 32.970 ;
        RECT 1490.560 20.390 1490.700 32.650 ;
        RECT 1490.500 20.070 1490.760 20.390 ;
        RECT 1323.060 19.050 1323.320 19.370 ;
        RECT 1323.120 2.400 1323.260 19.050 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1345.110 1686.980 1345.430 1687.040 ;
        RECT 1701.150 1686.980 1701.470 1687.040 ;
        RECT 1345.110 1686.840 1701.470 1686.980 ;
        RECT 1345.110 1686.780 1345.430 1686.840 ;
        RECT 1701.150 1686.780 1701.470 1686.840 ;
        RECT 1340.510 20.640 1340.830 20.700 ;
        RECT 1345.110 20.640 1345.430 20.700 ;
        RECT 1340.510 20.500 1345.430 20.640 ;
        RECT 1340.510 20.440 1340.830 20.500 ;
        RECT 1345.110 20.440 1345.430 20.500 ;
      LAYER via ;
        RECT 1345.140 1686.780 1345.400 1687.040 ;
        RECT 1701.180 1686.780 1701.440 1687.040 ;
        RECT 1340.540 20.440 1340.800 20.700 ;
        RECT 1345.140 20.440 1345.400 20.700 ;
      LAYER met2 ;
        RECT 1701.105 1700.000 1701.385 1704.000 ;
        RECT 1701.240 1687.070 1701.380 1700.000 ;
        RECT 1345.140 1686.750 1345.400 1687.070 ;
        RECT 1701.180 1686.750 1701.440 1687.070 ;
        RECT 1345.200 20.730 1345.340 1686.750 ;
        RECT 1340.540 20.410 1340.800 20.730 ;
        RECT 1345.140 20.410 1345.400 20.730 ;
        RECT 1340.600 2.400 1340.740 20.410 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 698.350 46.820 698.670 46.880 ;
        RECT 1435.730 46.820 1436.050 46.880 ;
        RECT 698.350 46.680 1436.050 46.820 ;
        RECT 698.350 46.620 698.670 46.680 ;
        RECT 1435.730 46.620 1436.050 46.680 ;
      LAYER via ;
        RECT 698.380 46.620 698.640 46.880 ;
        RECT 1435.760 46.620 1436.020 46.880 ;
      LAYER met2 ;
        RECT 1436.145 1700.410 1436.425 1704.000 ;
        RECT 1435.820 1700.270 1436.425 1700.410 ;
        RECT 1435.820 46.910 1435.960 1700.270 ;
        RECT 1436.145 1700.000 1436.425 1700.270 ;
        RECT 698.380 46.590 698.640 46.910 ;
        RECT 1435.760 46.590 1436.020 46.910 ;
        RECT 698.440 2.400 698.580 46.590 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1376.465 1685.805 1376.635 1689.035 ;
        RECT 1393.945 1688.865 1394.115 1690.055 ;
        RECT 1435.345 1689.885 1435.515 1690.735 ;
        RECT 1483.185 1689.205 1483.355 1690.735 ;
        RECT 1531.945 1689.205 1532.115 1690.735 ;
        RECT 1579.785 1689.205 1579.955 1690.735 ;
        RECT 1635.445 1687.165 1635.615 1689.375 ;
        RECT 1683.745 1687.165 1683.915 1694.135 ;
      LAYER mcon ;
        RECT 1683.745 1693.965 1683.915 1694.135 ;
        RECT 1435.345 1690.565 1435.515 1690.735 ;
        RECT 1393.945 1689.885 1394.115 1690.055 ;
        RECT 1483.185 1690.565 1483.355 1690.735 ;
        RECT 1531.945 1690.565 1532.115 1690.735 ;
        RECT 1579.785 1690.565 1579.955 1690.735 ;
        RECT 1635.445 1689.205 1635.615 1689.375 ;
        RECT 1376.465 1688.865 1376.635 1689.035 ;
      LAYER met1 ;
        RECT 1683.685 1694.120 1683.975 1694.165 ;
        RECT 1708.050 1694.120 1708.370 1694.180 ;
        RECT 1683.685 1693.980 1708.370 1694.120 ;
        RECT 1683.685 1693.935 1683.975 1693.980 ;
        RECT 1708.050 1693.920 1708.370 1693.980 ;
        RECT 1435.285 1690.720 1435.575 1690.765 ;
        RECT 1483.125 1690.720 1483.415 1690.765 ;
        RECT 1435.285 1690.580 1483.415 1690.720 ;
        RECT 1435.285 1690.535 1435.575 1690.580 ;
        RECT 1483.125 1690.535 1483.415 1690.580 ;
        RECT 1531.885 1690.720 1532.175 1690.765 ;
        RECT 1579.725 1690.720 1580.015 1690.765 ;
        RECT 1531.885 1690.580 1580.015 1690.720 ;
        RECT 1531.885 1690.535 1532.175 1690.580 ;
        RECT 1579.725 1690.535 1580.015 1690.580 ;
        RECT 1393.885 1690.040 1394.175 1690.085 ;
        RECT 1435.285 1690.040 1435.575 1690.085 ;
        RECT 1393.885 1689.900 1435.575 1690.040 ;
        RECT 1393.885 1689.855 1394.175 1689.900 ;
        RECT 1435.285 1689.855 1435.575 1689.900 ;
        RECT 1483.125 1689.360 1483.415 1689.405 ;
        RECT 1531.885 1689.360 1532.175 1689.405 ;
        RECT 1483.125 1689.220 1532.175 1689.360 ;
        RECT 1483.125 1689.175 1483.415 1689.220 ;
        RECT 1531.885 1689.175 1532.175 1689.220 ;
        RECT 1579.725 1689.360 1580.015 1689.405 ;
        RECT 1587.070 1689.360 1587.390 1689.420 ;
        RECT 1579.725 1689.220 1587.390 1689.360 ;
        RECT 1579.725 1689.175 1580.015 1689.220 ;
        RECT 1587.070 1689.160 1587.390 1689.220 ;
        RECT 1634.910 1689.360 1635.230 1689.420 ;
        RECT 1635.385 1689.360 1635.675 1689.405 ;
        RECT 1634.910 1689.220 1635.675 1689.360 ;
        RECT 1634.910 1689.160 1635.230 1689.220 ;
        RECT 1635.385 1689.175 1635.675 1689.220 ;
        RECT 1376.405 1689.020 1376.695 1689.065 ;
        RECT 1393.885 1689.020 1394.175 1689.065 ;
        RECT 1376.405 1688.880 1394.175 1689.020 ;
        RECT 1376.405 1688.835 1376.695 1688.880 ;
        RECT 1393.885 1688.835 1394.175 1688.880 ;
        RECT 1635.385 1687.320 1635.675 1687.365 ;
        RECT 1683.685 1687.320 1683.975 1687.365 ;
        RECT 1635.385 1687.180 1683.975 1687.320 ;
        RECT 1635.385 1687.135 1635.675 1687.180 ;
        RECT 1683.685 1687.135 1683.975 1687.180 ;
        RECT 1358.910 1685.960 1359.230 1686.020 ;
        RECT 1376.405 1685.960 1376.695 1686.005 ;
        RECT 1358.910 1685.820 1376.695 1685.960 ;
        RECT 1358.910 1685.760 1359.230 1685.820 ;
        RECT 1376.405 1685.775 1376.695 1685.820 ;
      LAYER via ;
        RECT 1708.080 1693.920 1708.340 1694.180 ;
        RECT 1587.100 1689.160 1587.360 1689.420 ;
        RECT 1634.940 1689.160 1635.200 1689.420 ;
        RECT 1358.940 1685.760 1359.200 1686.020 ;
      LAYER met2 ;
        RECT 1708.005 1700.000 1708.285 1704.000 ;
        RECT 1708.140 1694.210 1708.280 1700.000 ;
        RECT 1708.080 1693.890 1708.340 1694.210 ;
        RECT 1587.100 1689.130 1587.360 1689.450 ;
        RECT 1634.940 1689.130 1635.200 1689.450 ;
        RECT 1587.160 1688.965 1587.300 1689.130 ;
        RECT 1635.000 1688.965 1635.140 1689.130 ;
        RECT 1587.090 1688.595 1587.370 1688.965 ;
        RECT 1634.930 1688.595 1635.210 1688.965 ;
        RECT 1358.940 1685.730 1359.200 1686.050 ;
        RECT 1359.000 3.130 1359.140 1685.730 ;
        RECT 1358.540 2.990 1359.140 3.130 ;
        RECT 1358.540 2.400 1358.680 2.990 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
      LAYER via2 ;
        RECT 1587.090 1688.640 1587.370 1688.920 ;
        RECT 1634.930 1688.640 1635.210 1688.920 ;
      LAYER met3 ;
        RECT 1587.065 1688.930 1587.395 1688.945 ;
        RECT 1634.905 1688.930 1635.235 1688.945 ;
        RECT 1587.065 1688.630 1635.235 1688.930 ;
        RECT 1587.065 1688.615 1587.395 1688.630 ;
        RECT 1634.905 1688.615 1635.235 1688.630 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1635.905 1684.105 1636.075 1687.675 ;
      LAYER mcon ;
        RECT 1635.905 1687.505 1636.075 1687.675 ;
      LAYER met1 ;
        RECT 1379.610 1687.660 1379.930 1687.720 ;
        RECT 1635.845 1687.660 1636.135 1687.705 ;
        RECT 1379.610 1687.520 1636.135 1687.660 ;
        RECT 1379.610 1687.460 1379.930 1687.520 ;
        RECT 1635.845 1687.475 1636.135 1687.520 ;
        RECT 1635.845 1684.260 1636.135 1684.305 ;
        RECT 1715.410 1684.260 1715.730 1684.320 ;
        RECT 1635.845 1684.120 1715.730 1684.260 ;
        RECT 1635.845 1684.075 1636.135 1684.120 ;
        RECT 1715.410 1684.060 1715.730 1684.120 ;
        RECT 1376.390 14.520 1376.710 14.580 ;
        RECT 1379.610 14.520 1379.930 14.580 ;
        RECT 1376.390 14.380 1379.930 14.520 ;
        RECT 1376.390 14.320 1376.710 14.380 ;
        RECT 1379.610 14.320 1379.930 14.380 ;
      LAYER via ;
        RECT 1379.640 1687.460 1379.900 1687.720 ;
        RECT 1715.440 1684.060 1715.700 1684.320 ;
        RECT 1376.420 14.320 1376.680 14.580 ;
        RECT 1379.640 14.320 1379.900 14.580 ;
      LAYER met2 ;
        RECT 1715.365 1700.000 1715.645 1704.000 ;
        RECT 1379.640 1687.430 1379.900 1687.750 ;
        RECT 1379.700 14.610 1379.840 1687.430 ;
        RECT 1715.500 1684.350 1715.640 1700.000 ;
        RECT 1715.440 1684.030 1715.700 1684.350 ;
        RECT 1376.420 14.290 1376.680 14.610 ;
        RECT 1379.640 14.290 1379.900 14.610 ;
        RECT 1376.480 2.400 1376.620 14.290 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1443.165 16.405 1443.335 19.295 ;
        RECT 1462.485 16.405 1462.655 18.615 ;
        RECT 1631.765 18.445 1631.935 19.635 ;
        RECT 1661.205 18.785 1661.375 19.635 ;
      LAYER mcon ;
        RECT 1631.765 19.465 1631.935 19.635 ;
        RECT 1443.165 19.125 1443.335 19.295 ;
        RECT 1661.205 19.465 1661.375 19.635 ;
        RECT 1462.485 18.445 1462.655 18.615 ;
      LAYER met1 ;
        RECT 1680.450 1689.360 1680.770 1689.420 ;
        RECT 1722.770 1689.360 1723.090 1689.420 ;
        RECT 1680.450 1689.220 1723.090 1689.360 ;
        RECT 1680.450 1689.160 1680.770 1689.220 ;
        RECT 1722.770 1689.160 1723.090 1689.220 ;
        RECT 1631.705 19.620 1631.995 19.665 ;
        RECT 1661.145 19.620 1661.435 19.665 ;
        RECT 1631.705 19.480 1661.435 19.620 ;
        RECT 1631.705 19.435 1631.995 19.480 ;
        RECT 1661.145 19.435 1661.435 19.480 ;
        RECT 1443.105 19.280 1443.395 19.325 ;
        RECT 1429.380 19.140 1443.395 19.280 ;
        RECT 1394.330 18.940 1394.650 19.000 ;
        RECT 1429.380 18.940 1429.520 19.140 ;
        RECT 1443.105 19.095 1443.395 19.140 ;
        RECT 1394.330 18.800 1429.520 18.940 ;
        RECT 1661.145 18.940 1661.435 18.985 ;
        RECT 1677.690 18.940 1678.010 19.000 ;
        RECT 1661.145 18.800 1678.010 18.940 ;
        RECT 1394.330 18.740 1394.650 18.800 ;
        RECT 1661.145 18.755 1661.435 18.800 ;
        RECT 1677.690 18.740 1678.010 18.800 ;
        RECT 1462.425 18.600 1462.715 18.645 ;
        RECT 1631.705 18.600 1631.995 18.645 ;
        RECT 1462.425 18.460 1631.995 18.600 ;
        RECT 1462.425 18.415 1462.715 18.460 ;
        RECT 1631.705 18.415 1631.995 18.460 ;
        RECT 1443.105 16.560 1443.395 16.605 ;
        RECT 1462.425 16.560 1462.715 16.605 ;
        RECT 1443.105 16.420 1462.715 16.560 ;
        RECT 1443.105 16.375 1443.395 16.420 ;
        RECT 1462.425 16.375 1462.715 16.420 ;
      LAYER via ;
        RECT 1680.480 1689.160 1680.740 1689.420 ;
        RECT 1722.800 1689.160 1723.060 1689.420 ;
        RECT 1394.360 18.740 1394.620 19.000 ;
        RECT 1677.720 18.740 1677.980 19.000 ;
      LAYER met2 ;
        RECT 1722.725 1700.000 1723.005 1704.000 ;
        RECT 1722.860 1689.450 1723.000 1700.000 ;
        RECT 1680.480 1689.130 1680.740 1689.450 ;
        RECT 1722.800 1689.130 1723.060 1689.450 ;
        RECT 1680.540 1665.050 1680.680 1689.130 ;
        RECT 1680.080 1664.910 1680.680 1665.050 ;
        RECT 1394.360 18.710 1394.620 19.030 ;
        RECT 1677.720 18.770 1677.980 19.030 ;
        RECT 1680.080 18.770 1680.220 1664.910 ;
        RECT 1677.720 18.710 1680.220 18.770 ;
        RECT 1394.420 2.400 1394.560 18.710 ;
        RECT 1677.780 18.630 1680.220 18.710 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1604.165 17.765 1604.335 19.635 ;
        RECT 1613.825 15.385 1613.995 17.935 ;
      LAYER mcon ;
        RECT 1604.165 19.465 1604.335 19.635 ;
        RECT 1613.825 17.765 1613.995 17.935 ;
      LAYER met1 ;
        RECT 1638.590 1684.600 1638.910 1684.660 ;
        RECT 1727.370 1684.600 1727.690 1684.660 ;
        RECT 1638.590 1684.460 1727.690 1684.600 ;
        RECT 1638.590 1684.400 1638.910 1684.460 ;
        RECT 1727.370 1684.400 1727.690 1684.460 ;
        RECT 1412.270 19.620 1412.590 19.680 ;
        RECT 1604.105 19.620 1604.395 19.665 ;
        RECT 1412.270 19.480 1604.395 19.620 ;
        RECT 1412.270 19.420 1412.590 19.480 ;
        RECT 1604.105 19.435 1604.395 19.480 ;
        RECT 1604.105 17.920 1604.395 17.965 ;
        RECT 1613.765 17.920 1614.055 17.965 ;
        RECT 1604.105 17.780 1614.055 17.920 ;
        RECT 1604.105 17.735 1604.395 17.780 ;
        RECT 1613.765 17.735 1614.055 17.780 ;
        RECT 1613.765 15.540 1614.055 15.585 ;
        RECT 1638.590 15.540 1638.910 15.600 ;
        RECT 1613.765 15.400 1638.910 15.540 ;
        RECT 1613.765 15.355 1614.055 15.400 ;
        RECT 1638.590 15.340 1638.910 15.400 ;
      LAYER via ;
        RECT 1638.620 1684.400 1638.880 1684.660 ;
        RECT 1727.400 1684.400 1727.660 1684.660 ;
        RECT 1412.300 19.420 1412.560 19.680 ;
        RECT 1638.620 15.340 1638.880 15.600 ;
      LAYER met2 ;
        RECT 1730.085 1700.410 1730.365 1704.000 ;
        RECT 1728.380 1700.270 1730.365 1700.410 ;
        RECT 1728.380 1685.450 1728.520 1700.270 ;
        RECT 1730.085 1700.000 1730.365 1700.270 ;
        RECT 1727.460 1685.310 1728.520 1685.450 ;
        RECT 1727.460 1684.690 1727.600 1685.310 ;
        RECT 1638.620 1684.370 1638.880 1684.690 ;
        RECT 1727.400 1684.370 1727.660 1684.690 ;
        RECT 1412.300 19.390 1412.560 19.710 ;
        RECT 1412.360 2.400 1412.500 19.390 ;
        RECT 1638.680 15.630 1638.820 1684.370 ;
        RECT 1638.620 15.310 1638.880 15.630 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1660.745 17.765 1660.915 18.955 ;
        RECT 1676.845 17.765 1677.015 20.655 ;
      LAYER mcon ;
        RECT 1676.845 20.485 1677.015 20.655 ;
        RECT 1660.745 18.785 1660.915 18.955 ;
      LAYER met1 ;
        RECT 1693.790 1687.320 1694.110 1687.380 ;
        RECT 1737.490 1687.320 1737.810 1687.380 ;
        RECT 1693.790 1687.180 1737.810 1687.320 ;
        RECT 1693.790 1687.120 1694.110 1687.180 ;
        RECT 1737.490 1687.120 1737.810 1687.180 ;
        RECT 1676.785 20.640 1677.075 20.685 ;
        RECT 1693.790 20.640 1694.110 20.700 ;
        RECT 1676.785 20.500 1694.110 20.640 ;
        RECT 1676.785 20.455 1677.075 20.500 ;
        RECT 1693.790 20.440 1694.110 20.500 ;
        RECT 1429.750 18.940 1430.070 19.000 ;
        RECT 1660.685 18.940 1660.975 18.985 ;
        RECT 1429.750 18.800 1660.975 18.940 ;
        RECT 1429.750 18.740 1430.070 18.800 ;
        RECT 1660.685 18.755 1660.975 18.800 ;
        RECT 1660.685 17.920 1660.975 17.965 ;
        RECT 1676.785 17.920 1677.075 17.965 ;
        RECT 1660.685 17.780 1677.075 17.920 ;
        RECT 1660.685 17.735 1660.975 17.780 ;
        RECT 1676.785 17.735 1677.075 17.780 ;
      LAYER via ;
        RECT 1693.820 1687.120 1694.080 1687.380 ;
        RECT 1737.520 1687.120 1737.780 1687.380 ;
        RECT 1693.820 20.440 1694.080 20.700 ;
        RECT 1429.780 18.740 1430.040 19.000 ;
      LAYER met2 ;
        RECT 1737.445 1700.000 1737.725 1704.000 ;
        RECT 1737.580 1687.410 1737.720 1700.000 ;
        RECT 1693.820 1687.090 1694.080 1687.410 ;
        RECT 1737.520 1687.090 1737.780 1687.410 ;
        RECT 1693.880 20.730 1694.020 1687.090 ;
        RECT 1693.820 20.410 1694.080 20.730 ;
        RECT 1429.780 18.710 1430.040 19.030 ;
        RECT 1429.840 2.400 1429.980 18.710 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1709.430 1685.620 1709.750 1685.680 ;
        RECT 1744.850 1685.620 1745.170 1685.680 ;
        RECT 1709.430 1685.480 1745.170 1685.620 ;
        RECT 1709.430 1685.420 1709.750 1685.480 ;
        RECT 1744.850 1685.420 1745.170 1685.480 ;
        RECT 1447.690 19.280 1448.010 19.340 ;
        RECT 1447.690 19.140 1678.840 19.280 ;
        RECT 1447.690 19.080 1448.010 19.140 ;
        RECT 1678.700 18.940 1678.840 19.140 ;
        RECT 1707.590 18.940 1707.910 19.000 ;
        RECT 1678.700 18.800 1707.910 18.940 ;
        RECT 1707.590 18.740 1707.910 18.800 ;
      LAYER via ;
        RECT 1709.460 1685.420 1709.720 1685.680 ;
        RECT 1744.880 1685.420 1745.140 1685.680 ;
        RECT 1447.720 19.080 1447.980 19.340 ;
        RECT 1707.620 18.740 1707.880 19.000 ;
      LAYER met2 ;
        RECT 1744.805 1700.000 1745.085 1704.000 ;
        RECT 1744.940 1685.710 1745.080 1700.000 ;
        RECT 1709.460 1685.390 1709.720 1685.710 ;
        RECT 1744.880 1685.390 1745.140 1685.710 ;
        RECT 1709.520 1656.210 1709.660 1685.390 ;
        RECT 1707.680 1656.070 1709.660 1656.210 ;
        RECT 1447.720 19.050 1447.980 19.370 ;
        RECT 1447.780 2.400 1447.920 19.050 ;
        RECT 1707.680 19.030 1707.820 1656.070 ;
        RECT 1707.620 18.710 1707.880 19.030 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1562.690 1686.300 1563.010 1686.360 ;
        RECT 1752.210 1686.300 1752.530 1686.360 ;
        RECT 1562.690 1686.160 1752.530 1686.300 ;
        RECT 1562.690 1686.100 1563.010 1686.160 ;
        RECT 1752.210 1686.100 1752.530 1686.160 ;
        RECT 1465.630 15.200 1465.950 15.260 ;
        RECT 1562.690 15.200 1563.010 15.260 ;
        RECT 1465.630 15.060 1563.010 15.200 ;
        RECT 1465.630 15.000 1465.950 15.060 ;
        RECT 1562.690 15.000 1563.010 15.060 ;
      LAYER via ;
        RECT 1562.720 1686.100 1562.980 1686.360 ;
        RECT 1752.240 1686.100 1752.500 1686.360 ;
        RECT 1465.660 15.000 1465.920 15.260 ;
        RECT 1562.720 15.000 1562.980 15.260 ;
      LAYER met2 ;
        RECT 1752.165 1700.000 1752.445 1704.000 ;
        RECT 1752.300 1686.390 1752.440 1700.000 ;
        RECT 1562.720 1686.070 1562.980 1686.390 ;
        RECT 1752.240 1686.070 1752.500 1686.390 ;
        RECT 1562.780 15.290 1562.920 1686.070 ;
        RECT 1465.660 14.970 1465.920 15.290 ;
        RECT 1562.720 14.970 1562.980 15.290 ;
        RECT 1465.720 2.400 1465.860 14.970 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1535.165 1687.165 1535.335 1689.035 ;
      LAYER mcon ;
        RECT 1535.165 1688.865 1535.335 1689.035 ;
      LAYER met1 ;
        RECT 1535.105 1689.020 1535.395 1689.065 ;
        RECT 1759.570 1689.020 1759.890 1689.080 ;
        RECT 1535.105 1688.880 1759.890 1689.020 ;
        RECT 1535.105 1688.835 1535.395 1688.880 ;
        RECT 1759.570 1688.820 1759.890 1688.880 ;
        RECT 1489.550 1687.320 1489.870 1687.380 ;
        RECT 1535.105 1687.320 1535.395 1687.365 ;
        RECT 1489.550 1687.180 1535.395 1687.320 ;
        RECT 1489.550 1687.120 1489.870 1687.180 ;
        RECT 1535.105 1687.135 1535.395 1687.180 ;
        RECT 1483.570 20.640 1483.890 20.700 ;
        RECT 1489.550 20.640 1489.870 20.700 ;
        RECT 1483.570 20.500 1489.870 20.640 ;
        RECT 1483.570 20.440 1483.890 20.500 ;
        RECT 1489.550 20.440 1489.870 20.500 ;
      LAYER via ;
        RECT 1759.600 1688.820 1759.860 1689.080 ;
        RECT 1489.580 1687.120 1489.840 1687.380 ;
        RECT 1483.600 20.440 1483.860 20.700 ;
        RECT 1489.580 20.440 1489.840 20.700 ;
      LAYER met2 ;
        RECT 1759.525 1700.000 1759.805 1704.000 ;
        RECT 1759.660 1689.110 1759.800 1700.000 ;
        RECT 1759.600 1688.790 1759.860 1689.110 ;
        RECT 1489.580 1687.090 1489.840 1687.410 ;
        RECT 1489.640 20.730 1489.780 1687.090 ;
        RECT 1483.600 20.410 1483.860 20.730 ;
        RECT 1489.580 20.410 1489.840 20.730 ;
        RECT 1483.660 2.400 1483.800 20.410 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1661.665 19.465 1661.835 20.655 ;
      LAYER mcon ;
        RECT 1661.665 20.485 1661.835 20.655 ;
      LAYER met1 ;
        RECT 1714.490 1687.660 1714.810 1687.720 ;
        RECT 1766.930 1687.660 1767.250 1687.720 ;
        RECT 1714.490 1687.520 1767.250 1687.660 ;
        RECT 1714.490 1687.460 1714.810 1687.520 ;
        RECT 1766.930 1687.460 1767.250 1687.520 ;
        RECT 1501.510 20.640 1501.830 20.700 ;
        RECT 1661.605 20.640 1661.895 20.685 ;
        RECT 1501.510 20.500 1661.895 20.640 ;
        RECT 1501.510 20.440 1501.830 20.500 ;
        RECT 1661.605 20.455 1661.895 20.500 ;
        RECT 1661.605 19.620 1661.895 19.665 ;
        RECT 1661.605 19.480 1679.300 19.620 ;
        RECT 1661.605 19.435 1661.895 19.480 ;
        RECT 1679.160 19.280 1679.300 19.480 ;
        RECT 1714.490 19.280 1714.810 19.340 ;
        RECT 1679.160 19.140 1714.810 19.280 ;
        RECT 1714.490 19.080 1714.810 19.140 ;
      LAYER via ;
        RECT 1714.520 1687.460 1714.780 1687.720 ;
        RECT 1766.960 1687.460 1767.220 1687.720 ;
        RECT 1501.540 20.440 1501.800 20.700 ;
        RECT 1714.520 19.080 1714.780 19.340 ;
      LAYER met2 ;
        RECT 1766.885 1700.000 1767.165 1704.000 ;
        RECT 1767.020 1687.750 1767.160 1700.000 ;
        RECT 1714.520 1687.430 1714.780 1687.750 ;
        RECT 1766.960 1687.430 1767.220 1687.750 ;
        RECT 1501.540 20.410 1501.800 20.730 ;
        RECT 1501.600 2.400 1501.740 20.410 ;
        RECT 1714.580 19.370 1714.720 1687.430 ;
        RECT 1714.520 19.050 1714.780 19.370 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1774.290 1684.260 1774.610 1684.320 ;
        RECT 1762.420 1684.120 1774.610 1684.260 ;
        RECT 1721.850 1683.920 1722.170 1683.980 ;
        RECT 1762.420 1683.920 1762.560 1684.120 ;
        RECT 1774.290 1684.060 1774.610 1684.120 ;
        RECT 1721.850 1683.780 1762.560 1683.920 ;
        RECT 1721.850 1683.720 1722.170 1683.780 ;
        RECT 1518.990 16.560 1519.310 16.620 ;
        RECT 1721.850 16.560 1722.170 16.620 ;
        RECT 1518.990 16.420 1722.170 16.560 ;
        RECT 1518.990 16.360 1519.310 16.420 ;
        RECT 1721.850 16.360 1722.170 16.420 ;
      LAYER via ;
        RECT 1721.880 1683.720 1722.140 1683.980 ;
        RECT 1774.320 1684.060 1774.580 1684.320 ;
        RECT 1519.020 16.360 1519.280 16.620 ;
        RECT 1721.880 16.360 1722.140 16.620 ;
      LAYER met2 ;
        RECT 1774.245 1700.000 1774.525 1704.000 ;
        RECT 1774.380 1684.350 1774.520 1700.000 ;
        RECT 1774.320 1684.030 1774.580 1684.350 ;
        RECT 1721.880 1683.690 1722.140 1684.010 ;
        RECT 1721.940 16.650 1722.080 1683.690 ;
        RECT 1519.020 16.330 1519.280 16.650 ;
        RECT 1721.880 16.330 1722.140 16.650 ;
        RECT 1519.080 2.400 1519.220 16.330 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 717.210 50.220 717.530 50.280 ;
        RECT 1442.630 50.220 1442.950 50.280 ;
        RECT 717.210 50.080 1442.950 50.220 ;
        RECT 717.210 50.020 717.530 50.080 ;
        RECT 1442.630 50.020 1442.950 50.080 ;
      LAYER via ;
        RECT 717.240 50.020 717.500 50.280 ;
        RECT 1442.660 50.020 1442.920 50.280 ;
      LAYER met2 ;
        RECT 1443.505 1700.410 1443.785 1704.000 ;
        RECT 1442.720 1700.270 1443.785 1700.410 ;
        RECT 1442.720 50.310 1442.860 1700.270 ;
        RECT 1443.505 1700.000 1443.785 1700.270 ;
        RECT 717.240 49.990 717.500 50.310 ;
        RECT 1442.660 49.990 1442.920 50.310 ;
        RECT 717.300 17.410 717.440 49.990 ;
        RECT 716.380 17.270 717.440 17.410 ;
        RECT 716.380 2.400 716.520 17.270 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1781.605 1700.410 1781.885 1704.000 ;
        RECT 1781.280 1700.270 1781.885 1700.410 ;
        RECT 1781.280 16.845 1781.420 1700.270 ;
        RECT 1781.605 1700.000 1781.885 1700.270 ;
        RECT 1536.950 16.475 1537.230 16.845 ;
        RECT 1781.210 16.475 1781.490 16.845 ;
        RECT 1537.020 2.400 1537.160 16.475 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
      LAYER via2 ;
        RECT 1536.950 16.520 1537.230 16.800 ;
        RECT 1781.210 16.520 1781.490 16.800 ;
      LAYER met3 ;
        RECT 1536.925 16.810 1537.255 16.825 ;
        RECT 1781.185 16.810 1781.515 16.825 ;
        RECT 1536.925 16.510 1781.515 16.810 ;
        RECT 1536.925 16.495 1537.255 16.510 ;
        RECT 1781.185 16.495 1781.515 16.510 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1727.445 16.575 1727.615 16.915 ;
        RECT 1727.445 16.405 1728.535 16.575 ;
        RECT 1728.365 16.065 1728.535 16.405 ;
        RECT 1750.905 16.065 1751.075 22.355 ;
      LAYER mcon ;
        RECT 1750.905 22.185 1751.075 22.355 ;
        RECT 1727.445 16.745 1727.615 16.915 ;
      LAYER met1 ;
        RECT 1762.790 1683.920 1763.110 1683.980 ;
        RECT 1789.010 1683.920 1789.330 1683.980 ;
        RECT 1762.790 1683.780 1789.330 1683.920 ;
        RECT 1762.790 1683.720 1763.110 1683.780 ;
        RECT 1789.010 1683.720 1789.330 1683.780 ;
        RECT 1750.845 22.340 1751.135 22.385 ;
        RECT 1762.790 22.340 1763.110 22.400 ;
        RECT 1750.845 22.200 1763.110 22.340 ;
        RECT 1750.845 22.155 1751.135 22.200 ;
        RECT 1762.790 22.140 1763.110 22.200 ;
        RECT 1554.870 16.900 1555.190 16.960 ;
        RECT 1727.385 16.900 1727.675 16.945 ;
        RECT 1554.870 16.760 1727.675 16.900 ;
        RECT 1554.870 16.700 1555.190 16.760 ;
        RECT 1727.385 16.715 1727.675 16.760 ;
        RECT 1728.305 16.220 1728.595 16.265 ;
        RECT 1750.845 16.220 1751.135 16.265 ;
        RECT 1728.305 16.080 1751.135 16.220 ;
        RECT 1728.305 16.035 1728.595 16.080 ;
        RECT 1750.845 16.035 1751.135 16.080 ;
      LAYER via ;
        RECT 1762.820 1683.720 1763.080 1683.980 ;
        RECT 1789.040 1683.720 1789.300 1683.980 ;
        RECT 1762.820 22.140 1763.080 22.400 ;
        RECT 1554.900 16.700 1555.160 16.960 ;
      LAYER met2 ;
        RECT 1788.965 1700.000 1789.245 1704.000 ;
        RECT 1789.100 1684.010 1789.240 1700.000 ;
        RECT 1762.820 1683.690 1763.080 1684.010 ;
        RECT 1789.040 1683.690 1789.300 1684.010 ;
        RECT 1762.880 22.430 1763.020 1683.690 ;
        RECT 1762.820 22.110 1763.080 22.430 ;
        RECT 1554.900 16.670 1555.160 16.990 ;
        RECT 1554.960 2.400 1555.100 16.670 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1752.745 20.145 1753.375 20.315 ;
        RECT 1753.205 18.105 1753.375 20.145 ;
        RECT 1775.285 19.805 1777.295 19.975 ;
        RECT 1775.285 18.105 1775.455 19.805 ;
      LAYER mcon ;
        RECT 1777.125 19.805 1777.295 19.975 ;
      LAYER met1 ;
        RECT 1572.810 20.300 1573.130 20.360 ;
        RECT 1752.685 20.300 1752.975 20.345 ;
        RECT 1572.810 20.160 1752.975 20.300 ;
        RECT 1572.810 20.100 1573.130 20.160 ;
        RECT 1752.685 20.115 1752.975 20.160 ;
        RECT 1777.065 19.960 1777.355 20.005 ;
        RECT 1795.450 19.960 1795.770 20.020 ;
        RECT 1777.065 19.820 1795.770 19.960 ;
        RECT 1777.065 19.775 1777.355 19.820 ;
        RECT 1795.450 19.760 1795.770 19.820 ;
        RECT 1753.145 18.260 1753.435 18.305 ;
        RECT 1775.225 18.260 1775.515 18.305 ;
        RECT 1753.145 18.120 1775.515 18.260 ;
        RECT 1753.145 18.075 1753.435 18.120 ;
        RECT 1775.225 18.075 1775.515 18.120 ;
      LAYER via ;
        RECT 1572.840 20.100 1573.100 20.360 ;
        RECT 1795.480 19.760 1795.740 20.020 ;
      LAYER met2 ;
        RECT 1796.325 1700.410 1796.605 1704.000 ;
        RECT 1795.540 1700.270 1796.605 1700.410 ;
        RECT 1572.840 20.070 1573.100 20.390 ;
        RECT 1572.900 2.400 1573.040 20.070 ;
        RECT 1795.540 20.050 1795.680 1700.270 ;
        RECT 1796.325 1700.000 1796.605 1700.270 ;
        RECT 1795.480 19.730 1795.740 20.050 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1727.905 14.025 1728.075 16.235 ;
        RECT 1778.505 14.025 1780.055 14.195 ;
      LAYER mcon ;
        RECT 1727.905 16.065 1728.075 16.235 ;
        RECT 1779.885 14.025 1780.055 14.195 ;
      LAYER met1 ;
        RECT 1783.490 1688.340 1783.810 1688.400 ;
        RECT 1803.730 1688.340 1804.050 1688.400 ;
        RECT 1783.490 1688.200 1804.050 1688.340 ;
        RECT 1783.490 1688.140 1783.810 1688.200 ;
        RECT 1803.730 1688.140 1804.050 1688.200 ;
        RECT 1590.290 16.220 1590.610 16.280 ;
        RECT 1727.845 16.220 1728.135 16.265 ;
        RECT 1590.290 16.080 1728.135 16.220 ;
        RECT 1590.290 16.020 1590.610 16.080 ;
        RECT 1727.845 16.035 1728.135 16.080 ;
        RECT 1727.845 14.180 1728.135 14.225 ;
        RECT 1778.445 14.180 1778.735 14.225 ;
        RECT 1727.845 14.040 1778.735 14.180 ;
        RECT 1727.845 13.995 1728.135 14.040 ;
        RECT 1778.445 13.995 1778.735 14.040 ;
        RECT 1779.825 14.180 1780.115 14.225 ;
        RECT 1783.490 14.180 1783.810 14.240 ;
        RECT 1779.825 14.040 1783.810 14.180 ;
        RECT 1779.825 13.995 1780.115 14.040 ;
        RECT 1783.490 13.980 1783.810 14.040 ;
      LAYER via ;
        RECT 1783.520 1688.140 1783.780 1688.400 ;
        RECT 1803.760 1688.140 1804.020 1688.400 ;
        RECT 1590.320 16.020 1590.580 16.280 ;
        RECT 1783.520 13.980 1783.780 14.240 ;
      LAYER met2 ;
        RECT 1803.685 1700.000 1803.965 1704.000 ;
        RECT 1803.820 1688.430 1803.960 1700.000 ;
        RECT 1783.520 1688.110 1783.780 1688.430 ;
        RECT 1803.760 1688.110 1804.020 1688.430 ;
        RECT 1590.320 15.990 1590.580 16.310 ;
        RECT 1590.380 2.400 1590.520 15.990 ;
        RECT 1783.580 14.270 1783.720 1688.110 ;
        RECT 1783.520 13.950 1783.780 14.270 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1809.250 17.920 1809.570 17.980 ;
        RECT 1776.220 17.780 1809.570 17.920 ;
        RECT 1608.230 17.580 1608.550 17.640 ;
        RECT 1776.220 17.580 1776.360 17.780 ;
        RECT 1809.250 17.720 1809.570 17.780 ;
        RECT 1608.230 17.440 1776.360 17.580 ;
        RECT 1608.230 17.380 1608.550 17.440 ;
      LAYER via ;
        RECT 1608.260 17.380 1608.520 17.640 ;
        RECT 1809.280 17.720 1809.540 17.980 ;
      LAYER met2 ;
        RECT 1811.045 1700.410 1811.325 1704.000 ;
        RECT 1809.340 1700.270 1811.325 1700.410 ;
        RECT 1809.340 18.010 1809.480 1700.270 ;
        RECT 1811.045 1700.000 1811.325 1700.270 ;
        RECT 1809.280 17.690 1809.540 18.010 ;
        RECT 1608.260 17.350 1608.520 17.670 ;
        RECT 1608.320 2.400 1608.460 17.350 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1752.745 14.535 1752.915 18.275 ;
        RECT 1752.745 14.365 1754.295 14.535 ;
        RECT 1778.045 14.365 1778.215 15.555 ;
      LAYER mcon ;
        RECT 1752.745 18.105 1752.915 18.275 ;
        RECT 1778.045 15.385 1778.215 15.555 ;
        RECT 1754.125 14.365 1754.295 14.535 ;
      LAYER met1 ;
        RECT 1797.290 1687.660 1797.610 1687.720 ;
        RECT 1818.450 1687.660 1818.770 1687.720 ;
        RECT 1797.290 1687.520 1818.770 1687.660 ;
        RECT 1797.290 1687.460 1797.610 1687.520 ;
        RECT 1818.450 1687.460 1818.770 1687.520 ;
        RECT 1626.170 18.260 1626.490 18.320 ;
        RECT 1752.685 18.260 1752.975 18.305 ;
        RECT 1626.170 18.120 1752.975 18.260 ;
        RECT 1626.170 18.060 1626.490 18.120 ;
        RECT 1752.685 18.075 1752.975 18.120 ;
        RECT 1777.985 15.540 1778.275 15.585 ;
        RECT 1797.290 15.540 1797.610 15.600 ;
        RECT 1777.985 15.400 1797.610 15.540 ;
        RECT 1777.985 15.355 1778.275 15.400 ;
        RECT 1797.290 15.340 1797.610 15.400 ;
        RECT 1754.065 14.520 1754.355 14.565 ;
        RECT 1777.985 14.520 1778.275 14.565 ;
        RECT 1754.065 14.380 1778.275 14.520 ;
        RECT 1754.065 14.335 1754.355 14.380 ;
        RECT 1777.985 14.335 1778.275 14.380 ;
      LAYER via ;
        RECT 1797.320 1687.460 1797.580 1687.720 ;
        RECT 1818.480 1687.460 1818.740 1687.720 ;
        RECT 1626.200 18.060 1626.460 18.320 ;
        RECT 1797.320 15.340 1797.580 15.600 ;
      LAYER met2 ;
        RECT 1818.405 1700.000 1818.685 1704.000 ;
        RECT 1818.540 1687.750 1818.680 1700.000 ;
        RECT 1797.320 1687.430 1797.580 1687.750 ;
        RECT 1818.480 1687.430 1818.740 1687.750 ;
        RECT 1626.200 18.030 1626.460 18.350 ;
        RECT 1626.260 2.400 1626.400 18.030 ;
        RECT 1797.380 15.630 1797.520 1687.430 ;
        RECT 1797.320 15.310 1797.580 15.630 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1777.585 13.685 1777.755 15.555 ;
      LAYER mcon ;
        RECT 1777.585 15.385 1777.755 15.555 ;
      LAYER met1 ;
        RECT 1811.090 1684.260 1811.410 1684.320 ;
        RECT 1825.810 1684.260 1826.130 1684.320 ;
        RECT 1811.090 1684.120 1826.130 1684.260 ;
        RECT 1811.090 1684.060 1811.410 1684.120 ;
        RECT 1825.810 1684.060 1826.130 1684.120 ;
        RECT 1644.110 15.540 1644.430 15.600 ;
        RECT 1777.525 15.540 1777.815 15.585 ;
        RECT 1644.110 15.400 1777.815 15.540 ;
        RECT 1644.110 15.340 1644.430 15.400 ;
        RECT 1777.525 15.355 1777.815 15.400 ;
        RECT 1811.090 14.520 1811.410 14.580 ;
        RECT 1778.980 14.380 1811.410 14.520 ;
        RECT 1777.525 13.840 1777.815 13.885 ;
        RECT 1778.980 13.840 1779.120 14.380 ;
        RECT 1811.090 14.320 1811.410 14.380 ;
        RECT 1777.525 13.700 1779.120 13.840 ;
        RECT 1777.525 13.655 1777.815 13.700 ;
      LAYER via ;
        RECT 1811.120 1684.060 1811.380 1684.320 ;
        RECT 1825.840 1684.060 1826.100 1684.320 ;
        RECT 1644.140 15.340 1644.400 15.600 ;
        RECT 1811.120 14.320 1811.380 14.580 ;
      LAYER met2 ;
        RECT 1825.765 1700.000 1826.045 1704.000 ;
        RECT 1825.900 1684.350 1826.040 1700.000 ;
        RECT 1811.120 1684.030 1811.380 1684.350 ;
        RECT 1825.840 1684.030 1826.100 1684.350 ;
        RECT 1644.140 15.310 1644.400 15.630 ;
        RECT 1644.200 2.400 1644.340 15.310 ;
        RECT 1811.180 14.610 1811.320 1684.030 ;
        RECT 1811.120 14.290 1811.380 14.610 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1666.190 1685.960 1666.510 1686.020 ;
        RECT 1833.170 1685.960 1833.490 1686.020 ;
        RECT 1666.190 1685.820 1833.490 1685.960 ;
        RECT 1666.190 1685.760 1666.510 1685.820 ;
        RECT 1833.170 1685.760 1833.490 1685.820 ;
        RECT 1662.050 20.640 1662.370 20.700 ;
        RECT 1666.190 20.640 1666.510 20.700 ;
        RECT 1662.050 20.500 1666.510 20.640 ;
        RECT 1662.050 20.440 1662.370 20.500 ;
        RECT 1666.190 20.440 1666.510 20.500 ;
      LAYER via ;
        RECT 1666.220 1685.760 1666.480 1686.020 ;
        RECT 1833.200 1685.760 1833.460 1686.020 ;
        RECT 1662.080 20.440 1662.340 20.700 ;
        RECT 1666.220 20.440 1666.480 20.700 ;
      LAYER met2 ;
        RECT 1833.125 1700.000 1833.405 1704.000 ;
        RECT 1833.260 1686.050 1833.400 1700.000 ;
        RECT 1666.220 1685.730 1666.480 1686.050 ;
        RECT 1833.200 1685.730 1833.460 1686.050 ;
        RECT 1666.280 20.730 1666.420 1685.730 ;
        RECT 1662.080 20.410 1662.340 20.730 ;
        RECT 1666.220 20.410 1666.480 20.730 ;
        RECT 1662.140 2.400 1662.280 20.410 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1801.505 14.875 1801.675 15.215 ;
        RECT 1801.505 14.705 1802.595 14.875 ;
      LAYER mcon ;
        RECT 1801.505 15.045 1801.675 15.215 ;
        RECT 1802.425 14.705 1802.595 14.875 ;
      LAYER met1 ;
        RECT 1836.390 1676.780 1836.710 1676.840 ;
        RECT 1839.610 1676.780 1839.930 1676.840 ;
        RECT 1836.390 1676.640 1839.930 1676.780 ;
        RECT 1836.390 1676.580 1836.710 1676.640 ;
        RECT 1839.610 1676.580 1839.930 1676.640 ;
        RECT 1679.530 15.200 1679.850 15.260 ;
        RECT 1801.445 15.200 1801.735 15.245 ;
        RECT 1679.530 15.060 1801.735 15.200 ;
        RECT 1679.530 15.000 1679.850 15.060 ;
        RECT 1801.445 15.015 1801.735 15.060 ;
        RECT 1802.365 14.860 1802.655 14.905 ;
        RECT 1802.365 14.720 1811.780 14.860 ;
        RECT 1802.365 14.675 1802.655 14.720 ;
        RECT 1811.640 14.520 1811.780 14.720 ;
        RECT 1836.390 14.520 1836.710 14.580 ;
        RECT 1811.640 14.380 1836.710 14.520 ;
        RECT 1836.390 14.320 1836.710 14.380 ;
      LAYER via ;
        RECT 1836.420 1676.580 1836.680 1676.840 ;
        RECT 1839.640 1676.580 1839.900 1676.840 ;
        RECT 1679.560 15.000 1679.820 15.260 ;
        RECT 1836.420 14.320 1836.680 14.580 ;
      LAYER met2 ;
        RECT 1840.485 1700.410 1840.765 1704.000 ;
        RECT 1839.700 1700.270 1840.765 1700.410 ;
        RECT 1839.700 1676.870 1839.840 1700.270 ;
        RECT 1840.485 1700.000 1840.765 1700.270 ;
        RECT 1836.420 1676.550 1836.680 1676.870 ;
        RECT 1839.640 1676.550 1839.900 1676.870 ;
        RECT 1679.560 14.970 1679.820 15.290 ;
        RECT 1679.620 2.400 1679.760 14.970 ;
        RECT 1836.480 14.610 1836.620 1676.550 ;
        RECT 1836.420 14.290 1836.680 14.610 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1703.910 1686.980 1704.230 1687.040 ;
        RECT 1847.890 1686.980 1848.210 1687.040 ;
        RECT 1703.910 1686.840 1848.210 1686.980 ;
        RECT 1703.910 1686.780 1704.230 1686.840 ;
        RECT 1847.890 1686.780 1848.210 1686.840 ;
        RECT 1697.470 20.640 1697.790 20.700 ;
        RECT 1703.910 20.640 1704.230 20.700 ;
        RECT 1697.470 20.500 1704.230 20.640 ;
        RECT 1697.470 20.440 1697.790 20.500 ;
        RECT 1703.910 20.440 1704.230 20.500 ;
      LAYER via ;
        RECT 1703.940 1686.780 1704.200 1687.040 ;
        RECT 1847.920 1686.780 1848.180 1687.040 ;
        RECT 1697.500 20.440 1697.760 20.700 ;
        RECT 1703.940 20.440 1704.200 20.700 ;
      LAYER met2 ;
        RECT 1847.845 1700.000 1848.125 1704.000 ;
        RECT 1847.980 1687.070 1848.120 1700.000 ;
        RECT 1703.940 1686.750 1704.200 1687.070 ;
        RECT 1847.920 1686.750 1848.180 1687.070 ;
        RECT 1704.000 20.730 1704.140 1686.750 ;
        RECT 1697.500 20.410 1697.760 20.730 ;
        RECT 1703.940 20.410 1704.200 20.730 ;
        RECT 1697.560 2.400 1697.700 20.410 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 737.910 49.880 738.230 49.940 ;
        RECT 1449.070 49.880 1449.390 49.940 ;
        RECT 737.910 49.740 1449.390 49.880 ;
        RECT 737.910 49.680 738.230 49.740 ;
        RECT 1449.070 49.680 1449.390 49.740 ;
      LAYER via ;
        RECT 737.940 49.680 738.200 49.940 ;
        RECT 1449.100 49.680 1449.360 49.940 ;
      LAYER met2 ;
        RECT 1450.865 1700.410 1451.145 1704.000 ;
        RECT 1449.160 1700.270 1451.145 1700.410 ;
        RECT 1449.160 49.970 1449.300 1700.270 ;
        RECT 1450.865 1700.000 1451.145 1700.270 ;
        RECT 737.940 49.650 738.200 49.970 ;
        RECT 1449.100 49.650 1449.360 49.970 ;
        RECT 738.000 17.410 738.140 49.650 ;
        RECT 734.320 17.270 738.140 17.410 ;
        RECT 734.320 2.400 734.460 17.270 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1845.590 1688.000 1845.910 1688.060 ;
        RECT 1855.250 1688.000 1855.570 1688.060 ;
        RECT 1845.590 1687.860 1855.570 1688.000 ;
        RECT 1845.590 1687.800 1845.910 1687.860 ;
        RECT 1855.250 1687.800 1855.570 1687.860 ;
        RECT 1715.410 19.280 1715.730 19.340 ;
        RECT 1845.590 19.280 1845.910 19.340 ;
        RECT 1715.410 19.140 1845.910 19.280 ;
        RECT 1715.410 19.080 1715.730 19.140 ;
        RECT 1845.590 19.080 1845.910 19.140 ;
      LAYER via ;
        RECT 1845.620 1687.800 1845.880 1688.060 ;
        RECT 1855.280 1687.800 1855.540 1688.060 ;
        RECT 1715.440 19.080 1715.700 19.340 ;
        RECT 1845.620 19.080 1845.880 19.340 ;
      LAYER met2 ;
        RECT 1855.205 1700.000 1855.485 1704.000 ;
        RECT 1855.340 1688.090 1855.480 1700.000 ;
        RECT 1845.620 1687.770 1845.880 1688.090 ;
        RECT 1855.280 1687.770 1855.540 1688.090 ;
        RECT 1845.680 19.370 1845.820 1687.770 ;
        RECT 1715.440 19.050 1715.700 19.370 ;
        RECT 1845.620 19.050 1845.880 19.370 ;
        RECT 1715.500 2.400 1715.640 19.050 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1852.490 1683.920 1852.810 1683.980 ;
        RECT 1862.610 1683.920 1862.930 1683.980 ;
        RECT 1852.490 1683.780 1862.930 1683.920 ;
        RECT 1852.490 1683.720 1852.810 1683.780 ;
        RECT 1862.610 1683.720 1862.930 1683.780 ;
        RECT 1733.350 15.880 1733.670 15.940 ;
        RECT 1852.490 15.880 1852.810 15.940 ;
        RECT 1733.350 15.740 1852.810 15.880 ;
        RECT 1733.350 15.680 1733.670 15.740 ;
        RECT 1852.490 15.680 1852.810 15.740 ;
      LAYER via ;
        RECT 1852.520 1683.720 1852.780 1683.980 ;
        RECT 1862.640 1683.720 1862.900 1683.980 ;
        RECT 1733.380 15.680 1733.640 15.940 ;
        RECT 1852.520 15.680 1852.780 15.940 ;
      LAYER met2 ;
        RECT 1862.565 1700.000 1862.845 1704.000 ;
        RECT 1862.700 1684.010 1862.840 1700.000 ;
        RECT 1852.520 1683.690 1852.780 1684.010 ;
        RECT 1862.640 1683.690 1862.900 1684.010 ;
        RECT 1852.580 15.970 1852.720 1683.690 ;
        RECT 1733.380 15.650 1733.640 15.970 ;
        RECT 1852.520 15.650 1852.780 15.970 ;
        RECT 1733.440 2.400 1733.580 15.650 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1762.405 16.065 1762.575 19.975 ;
      LAYER mcon ;
        RECT 1762.405 19.805 1762.575 19.975 ;
      LAYER met1 ;
        RECT 1869.970 20.300 1870.290 20.360 ;
        RECT 1763.800 20.160 1870.290 20.300 ;
        RECT 1762.345 19.960 1762.635 20.005 ;
        RECT 1763.800 19.960 1763.940 20.160 ;
        RECT 1869.970 20.100 1870.290 20.160 ;
        RECT 1762.345 19.820 1763.940 19.960 ;
        RECT 1762.345 19.775 1762.635 19.820 ;
        RECT 1751.290 16.220 1751.610 16.280 ;
        RECT 1762.345 16.220 1762.635 16.265 ;
        RECT 1751.290 16.080 1762.635 16.220 ;
        RECT 1751.290 16.020 1751.610 16.080 ;
        RECT 1762.345 16.035 1762.635 16.080 ;
      LAYER via ;
        RECT 1870.000 20.100 1870.260 20.360 ;
        RECT 1751.320 16.020 1751.580 16.280 ;
      LAYER met2 ;
        RECT 1869.925 1700.000 1870.205 1704.000 ;
        RECT 1870.060 20.390 1870.200 1700.000 ;
        RECT 1870.000 20.070 1870.260 20.390 ;
        RECT 1751.320 15.990 1751.580 16.310 ;
        RECT 1751.380 2.400 1751.520 15.990 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1768.770 16.900 1769.090 16.960 ;
        RECT 1878.250 16.900 1878.570 16.960 ;
        RECT 1768.770 16.760 1878.570 16.900 ;
        RECT 1768.770 16.700 1769.090 16.760 ;
        RECT 1878.250 16.700 1878.570 16.760 ;
      LAYER via ;
        RECT 1768.800 16.700 1769.060 16.960 ;
        RECT 1878.280 16.700 1878.540 16.960 ;
      LAYER met2 ;
        RECT 1877.285 1700.410 1877.565 1704.000 ;
        RECT 1877.285 1700.270 1878.480 1700.410 ;
        RECT 1877.285 1700.000 1877.565 1700.270 ;
        RECT 1878.340 16.990 1878.480 1700.270 ;
        RECT 1768.800 16.670 1769.060 16.990 ;
        RECT 1878.280 16.670 1878.540 16.990 ;
        RECT 1768.860 2.400 1769.000 16.670 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1880.090 1683.920 1880.410 1683.980 ;
        RECT 1884.690 1683.920 1885.010 1683.980 ;
        RECT 1880.090 1683.780 1885.010 1683.920 ;
        RECT 1880.090 1683.720 1880.410 1683.780 ;
        RECT 1884.690 1683.720 1885.010 1683.780 ;
        RECT 1786.710 16.220 1787.030 16.280 ;
        RECT 1880.090 16.220 1880.410 16.280 ;
        RECT 1786.710 16.080 1880.410 16.220 ;
        RECT 1786.710 16.020 1787.030 16.080 ;
        RECT 1880.090 16.020 1880.410 16.080 ;
      LAYER via ;
        RECT 1880.120 1683.720 1880.380 1683.980 ;
        RECT 1884.720 1683.720 1884.980 1683.980 ;
        RECT 1786.740 16.020 1787.000 16.280 ;
        RECT 1880.120 16.020 1880.380 16.280 ;
      LAYER met2 ;
        RECT 1884.645 1700.000 1884.925 1704.000 ;
        RECT 1884.780 1684.010 1884.920 1700.000 ;
        RECT 1880.120 1683.690 1880.380 1684.010 ;
        RECT 1884.720 1683.690 1884.980 1684.010 ;
        RECT 1880.180 16.310 1880.320 1683.690 ;
        RECT 1786.740 15.990 1787.000 16.310 ;
        RECT 1880.120 15.990 1880.380 16.310 ;
        RECT 1786.800 2.400 1786.940 15.990 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1888.370 1683.920 1888.690 1683.980 ;
        RECT 1892.050 1683.920 1892.370 1683.980 ;
        RECT 1888.370 1683.780 1892.370 1683.920 ;
        RECT 1888.370 1683.720 1888.690 1683.780 ;
        RECT 1892.050 1683.720 1892.370 1683.780 ;
        RECT 1804.650 18.260 1804.970 18.320 ;
        RECT 1886.990 18.260 1887.310 18.320 ;
        RECT 1804.650 18.120 1887.310 18.260 ;
        RECT 1804.650 18.060 1804.970 18.120 ;
        RECT 1886.990 18.060 1887.310 18.120 ;
      LAYER via ;
        RECT 1888.400 1683.720 1888.660 1683.980 ;
        RECT 1892.080 1683.720 1892.340 1683.980 ;
        RECT 1804.680 18.060 1804.940 18.320 ;
        RECT 1887.020 18.060 1887.280 18.320 ;
      LAYER met2 ;
        RECT 1892.005 1700.000 1892.285 1704.000 ;
        RECT 1892.140 1684.010 1892.280 1700.000 ;
        RECT 1888.400 1683.690 1888.660 1684.010 ;
        RECT 1892.080 1683.690 1892.340 1684.010 ;
        RECT 1888.460 1677.290 1888.600 1683.690 ;
        RECT 1887.080 1677.150 1888.600 1677.290 ;
        RECT 1887.080 18.350 1887.220 1677.150 ;
        RECT 1804.680 18.030 1804.940 18.350 ;
        RECT 1887.020 18.030 1887.280 18.350 ;
        RECT 1804.740 2.400 1804.880 18.030 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1851.645 16.575 1851.815 17.255 ;
        RECT 1849.345 16.405 1851.815 16.575 ;
      LAYER mcon ;
        RECT 1851.645 17.085 1851.815 17.255 ;
      LAYER met1 ;
        RECT 1851.585 17.240 1851.875 17.285 ;
        RECT 1898.490 17.240 1898.810 17.300 ;
        RECT 1851.585 17.100 1898.810 17.240 ;
        RECT 1851.585 17.055 1851.875 17.100 ;
        RECT 1898.490 17.040 1898.810 17.100 ;
        RECT 1827.650 16.560 1827.970 16.620 ;
        RECT 1849.285 16.560 1849.575 16.605 ;
        RECT 1827.650 16.420 1849.575 16.560 ;
        RECT 1827.650 16.360 1827.970 16.420 ;
        RECT 1849.285 16.375 1849.575 16.420 ;
        RECT 1822.590 15.200 1822.910 15.260 ;
        RECT 1827.650 15.200 1827.970 15.260 ;
        RECT 1822.590 15.060 1827.970 15.200 ;
        RECT 1822.590 15.000 1822.910 15.060 ;
        RECT 1827.650 15.000 1827.970 15.060 ;
      LAYER via ;
        RECT 1898.520 17.040 1898.780 17.300 ;
        RECT 1827.680 16.360 1827.940 16.620 ;
        RECT 1822.620 15.000 1822.880 15.260 ;
        RECT 1827.680 15.000 1827.940 15.260 ;
      LAYER met2 ;
        RECT 1899.365 1700.410 1899.645 1704.000 ;
        RECT 1898.580 1700.270 1899.645 1700.410 ;
        RECT 1898.580 17.330 1898.720 1700.270 ;
        RECT 1899.365 1700.000 1899.645 1700.270 ;
        RECT 1898.520 17.010 1898.780 17.330 ;
        RECT 1827.680 16.330 1827.940 16.650 ;
        RECT 1827.740 15.290 1827.880 16.330 ;
        RECT 1822.620 14.970 1822.880 15.290 ;
        RECT 1827.680 14.970 1827.940 15.290 ;
        RECT 1822.680 2.400 1822.820 14.970 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1884.305 17.595 1884.475 25.075 ;
        RECT 1883.845 17.425 1884.475 17.595 ;
      LAYER mcon ;
        RECT 1884.305 24.905 1884.475 25.075 ;
      LAYER met1 ;
        RECT 1900.790 1688.680 1901.110 1688.740 ;
        RECT 1906.770 1688.680 1907.090 1688.740 ;
        RECT 1900.790 1688.540 1907.090 1688.680 ;
        RECT 1900.790 1688.480 1901.110 1688.540 ;
        RECT 1906.770 1688.480 1907.090 1688.540 ;
        RECT 1884.245 25.060 1884.535 25.105 ;
        RECT 1900.790 25.060 1901.110 25.120 ;
        RECT 1884.245 24.920 1901.110 25.060 ;
        RECT 1884.245 24.875 1884.535 24.920 ;
        RECT 1900.790 24.860 1901.110 24.920 ;
        RECT 1883.785 17.580 1884.075 17.625 ;
        RECT 1851.200 17.440 1884.075 17.580 ;
        RECT 1840.070 17.240 1840.390 17.300 ;
        RECT 1851.200 17.240 1851.340 17.440 ;
        RECT 1883.785 17.395 1884.075 17.440 ;
        RECT 1840.070 17.100 1851.340 17.240 ;
        RECT 1840.070 17.040 1840.390 17.100 ;
      LAYER via ;
        RECT 1900.820 1688.480 1901.080 1688.740 ;
        RECT 1906.800 1688.480 1907.060 1688.740 ;
        RECT 1900.820 24.860 1901.080 25.120 ;
        RECT 1840.100 17.040 1840.360 17.300 ;
      LAYER met2 ;
        RECT 1906.725 1700.000 1907.005 1704.000 ;
        RECT 1906.860 1688.770 1907.000 1700.000 ;
        RECT 1900.820 1688.450 1901.080 1688.770 ;
        RECT 1906.800 1688.450 1907.060 1688.770 ;
        RECT 1900.880 25.150 1901.020 1688.450 ;
        RECT 1900.820 24.830 1901.080 25.150 ;
        RECT 1840.100 17.010 1840.360 17.330 ;
        RECT 1840.160 2.400 1840.300 17.010 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1883.845 19.465 1884.015 24.735 ;
      LAYER mcon ;
        RECT 1883.845 24.565 1884.015 24.735 ;
      LAYER met1 ;
        RECT 1907.690 1688.680 1908.010 1688.740 ;
        RECT 1914.130 1688.680 1914.450 1688.740 ;
        RECT 1907.690 1688.540 1914.450 1688.680 ;
        RECT 1907.690 1688.480 1908.010 1688.540 ;
        RECT 1914.130 1688.480 1914.450 1688.540 ;
        RECT 1883.785 24.720 1884.075 24.765 ;
        RECT 1907.690 24.720 1908.010 24.780 ;
        RECT 1883.785 24.580 1908.010 24.720 ;
        RECT 1883.785 24.535 1884.075 24.580 ;
        RECT 1907.690 24.520 1908.010 24.580 ;
        RECT 1858.010 19.620 1858.330 19.680 ;
        RECT 1883.785 19.620 1884.075 19.665 ;
        RECT 1858.010 19.480 1884.075 19.620 ;
        RECT 1858.010 19.420 1858.330 19.480 ;
        RECT 1883.785 19.435 1884.075 19.480 ;
      LAYER via ;
        RECT 1907.720 1688.480 1907.980 1688.740 ;
        RECT 1914.160 1688.480 1914.420 1688.740 ;
        RECT 1907.720 24.520 1907.980 24.780 ;
        RECT 1858.040 19.420 1858.300 19.680 ;
      LAYER met2 ;
        RECT 1914.085 1700.000 1914.365 1704.000 ;
        RECT 1914.220 1688.770 1914.360 1700.000 ;
        RECT 1907.720 1688.450 1907.980 1688.770 ;
        RECT 1914.160 1688.450 1914.420 1688.770 ;
        RECT 1907.780 24.810 1907.920 1688.450 ;
        RECT 1907.720 24.490 1907.980 24.810 ;
        RECT 1858.040 19.390 1858.300 19.710 ;
        RECT 1858.100 2.400 1858.240 19.390 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1875.950 18.600 1876.270 18.660 ;
        RECT 1919.190 18.600 1919.510 18.660 ;
        RECT 1875.950 18.460 1919.510 18.600 ;
        RECT 1875.950 18.400 1876.270 18.460 ;
        RECT 1919.190 18.400 1919.510 18.460 ;
      LAYER via ;
        RECT 1875.980 18.400 1876.240 18.660 ;
        RECT 1919.220 18.400 1919.480 18.660 ;
      LAYER met2 ;
        RECT 1921.445 1700.410 1921.725 1704.000 ;
        RECT 1919.280 1700.270 1921.725 1700.410 ;
        RECT 1919.280 18.690 1919.420 1700.270 ;
        RECT 1921.445 1700.000 1921.725 1700.270 ;
        RECT 1875.980 18.370 1876.240 18.690 ;
        RECT 1919.220 18.370 1919.480 18.690 ;
        RECT 1876.040 2.400 1876.180 18.370 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 758.150 49.540 758.470 49.600 ;
        RECT 1456.430 49.540 1456.750 49.600 ;
        RECT 758.150 49.400 1456.750 49.540 ;
        RECT 758.150 49.340 758.470 49.400 ;
        RECT 1456.430 49.340 1456.750 49.400 ;
        RECT 752.170 20.980 752.490 21.040 ;
        RECT 758.150 20.980 758.470 21.040 ;
        RECT 752.170 20.840 758.470 20.980 ;
        RECT 752.170 20.780 752.490 20.840 ;
        RECT 758.150 20.780 758.470 20.840 ;
      LAYER via ;
        RECT 758.180 49.340 758.440 49.600 ;
        RECT 1456.460 49.340 1456.720 49.600 ;
        RECT 752.200 20.780 752.460 21.040 ;
        RECT 758.180 20.780 758.440 21.040 ;
      LAYER met2 ;
        RECT 1458.225 1700.410 1458.505 1704.000 ;
        RECT 1456.520 1700.270 1458.505 1700.410 ;
        RECT 1456.520 49.630 1456.660 1700.270 ;
        RECT 1458.225 1700.000 1458.505 1700.270 ;
        RECT 758.180 49.310 758.440 49.630 ;
        RECT 1456.460 49.310 1456.720 49.630 ;
        RECT 758.240 21.070 758.380 49.310 ;
        RECT 752.200 20.750 752.460 21.070 ;
        RECT 758.180 20.750 758.440 21.070 ;
        RECT 752.260 2.400 752.400 20.750 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1893.890 20.640 1894.210 20.700 ;
        RECT 1926.550 20.640 1926.870 20.700 ;
        RECT 1893.890 20.500 1926.870 20.640 ;
        RECT 1893.890 20.440 1894.210 20.500 ;
        RECT 1926.550 20.440 1926.870 20.500 ;
      LAYER via ;
        RECT 1893.920 20.440 1894.180 20.700 ;
        RECT 1926.580 20.440 1926.840 20.700 ;
      LAYER met2 ;
        RECT 1928.805 1700.410 1929.085 1704.000 ;
        RECT 1926.640 1700.270 1929.085 1700.410 ;
        RECT 1926.640 20.730 1926.780 1700.270 ;
        RECT 1928.805 1700.000 1929.085 1700.270 ;
        RECT 1893.920 20.410 1894.180 20.730 ;
        RECT 1926.580 20.410 1926.840 20.730 ;
        RECT 1893.980 2.400 1894.120 20.410 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1911.830 17.920 1912.150 17.980 ;
        RECT 1932.990 17.920 1933.310 17.980 ;
        RECT 1911.830 17.780 1933.310 17.920 ;
        RECT 1911.830 17.720 1912.150 17.780 ;
        RECT 1932.990 17.720 1933.310 17.780 ;
      LAYER via ;
        RECT 1911.860 17.720 1912.120 17.980 ;
        RECT 1933.020 17.720 1933.280 17.980 ;
      LAYER met2 ;
        RECT 1936.165 1701.090 1936.445 1704.000 ;
        RECT 1934.000 1700.950 1936.445 1701.090 ;
        RECT 1934.000 1686.130 1934.140 1700.950 ;
        RECT 1936.165 1700.000 1936.445 1700.950 ;
        RECT 1933.080 1685.990 1934.140 1686.130 ;
        RECT 1933.080 18.010 1933.220 1685.990 ;
        RECT 1911.860 17.690 1912.120 18.010 ;
        RECT 1933.020 17.690 1933.280 18.010 ;
        RECT 1911.920 2.400 1912.060 17.690 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1935.290 1687.320 1935.610 1687.380 ;
        RECT 1943.570 1687.320 1943.890 1687.380 ;
        RECT 1935.290 1687.180 1943.890 1687.320 ;
        RECT 1935.290 1687.120 1935.610 1687.180 ;
        RECT 1943.570 1687.120 1943.890 1687.180 ;
        RECT 1929.310 14.520 1929.630 14.580 ;
        RECT 1935.290 14.520 1935.610 14.580 ;
        RECT 1929.310 14.380 1935.610 14.520 ;
        RECT 1929.310 14.320 1929.630 14.380 ;
        RECT 1935.290 14.320 1935.610 14.380 ;
      LAYER via ;
        RECT 1935.320 1687.120 1935.580 1687.380 ;
        RECT 1943.600 1687.120 1943.860 1687.380 ;
        RECT 1929.340 14.320 1929.600 14.580 ;
        RECT 1935.320 14.320 1935.580 14.580 ;
      LAYER met2 ;
        RECT 1943.525 1700.000 1943.805 1704.000 ;
        RECT 1943.660 1687.410 1943.800 1700.000 ;
        RECT 1935.320 1687.090 1935.580 1687.410 ;
        RECT 1943.600 1687.090 1943.860 1687.410 ;
        RECT 1935.380 14.610 1935.520 1687.090 ;
        RECT 1929.340 14.290 1929.600 14.610 ;
        RECT 1935.320 14.290 1935.580 14.610 ;
        RECT 1929.400 2.400 1929.540 14.290 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1947.325 1594.005 1947.495 1642.115 ;
        RECT 1946.865 1400.885 1947.035 1448.995 ;
        RECT 1946.865 1304.325 1947.035 1352.435 ;
        RECT 1946.865 517.565 1947.035 607.155 ;
        RECT 1946.405 448.205 1946.575 493.595 ;
        RECT 1946.865 331.245 1947.035 379.355 ;
        RECT 1945.945 241.485 1946.115 287.895 ;
        RECT 1946.865 83.045 1947.035 131.155 ;
        RECT 1947.325 2.805 1947.495 17.595 ;
      LAYER mcon ;
        RECT 1947.325 1641.945 1947.495 1642.115 ;
        RECT 1946.865 1448.825 1947.035 1448.995 ;
        RECT 1946.865 1352.265 1947.035 1352.435 ;
        RECT 1946.865 606.985 1947.035 607.155 ;
        RECT 1946.405 493.425 1946.575 493.595 ;
        RECT 1946.865 379.185 1947.035 379.355 ;
        RECT 1945.945 287.725 1946.115 287.895 ;
        RECT 1946.865 130.985 1947.035 131.155 ;
        RECT 1947.325 17.425 1947.495 17.595 ;
      LAYER met1 ;
        RECT 1946.330 1656.040 1946.650 1656.100 ;
        RECT 1947.250 1656.040 1947.570 1656.100 ;
        RECT 1946.330 1655.900 1947.570 1656.040 ;
        RECT 1946.330 1655.840 1946.650 1655.900 ;
        RECT 1947.250 1655.840 1947.570 1655.900 ;
        RECT 1947.250 1642.100 1947.570 1642.160 ;
        RECT 1947.055 1641.960 1947.570 1642.100 ;
        RECT 1947.250 1641.900 1947.570 1641.960 ;
        RECT 1947.265 1594.160 1947.555 1594.205 ;
        RECT 1947.710 1594.160 1948.030 1594.220 ;
        RECT 1947.265 1594.020 1948.030 1594.160 ;
        RECT 1947.265 1593.975 1947.555 1594.020 ;
        RECT 1947.710 1593.960 1948.030 1594.020 ;
        RECT 1946.790 1559.480 1947.110 1559.540 ;
        RECT 1947.710 1559.480 1948.030 1559.540 ;
        RECT 1946.790 1559.340 1948.030 1559.480 ;
        RECT 1946.790 1559.280 1947.110 1559.340 ;
        RECT 1947.710 1559.280 1948.030 1559.340 ;
        RECT 1945.870 1511.200 1946.190 1511.260 ;
        RECT 1946.790 1511.200 1947.110 1511.260 ;
        RECT 1945.870 1511.060 1947.110 1511.200 ;
        RECT 1945.870 1511.000 1946.190 1511.060 ;
        RECT 1946.790 1511.000 1947.110 1511.060 ;
        RECT 1946.805 1448.980 1947.095 1449.025 ;
        RECT 1947.250 1448.980 1947.570 1449.040 ;
        RECT 1946.805 1448.840 1947.570 1448.980 ;
        RECT 1946.805 1448.795 1947.095 1448.840 ;
        RECT 1947.250 1448.780 1947.570 1448.840 ;
        RECT 1946.790 1401.040 1947.110 1401.100 ;
        RECT 1946.595 1400.900 1947.110 1401.040 ;
        RECT 1946.790 1400.840 1947.110 1400.900 ;
        RECT 1946.805 1352.420 1947.095 1352.465 ;
        RECT 1947.250 1352.420 1947.570 1352.480 ;
        RECT 1946.805 1352.280 1947.570 1352.420 ;
        RECT 1946.805 1352.235 1947.095 1352.280 ;
        RECT 1947.250 1352.220 1947.570 1352.280 ;
        RECT 1946.790 1304.480 1947.110 1304.540 ;
        RECT 1946.595 1304.340 1947.110 1304.480 ;
        RECT 1946.790 1304.280 1947.110 1304.340 ;
        RECT 1945.870 1256.200 1946.190 1256.260 ;
        RECT 1946.790 1256.200 1947.110 1256.260 ;
        RECT 1945.870 1256.060 1947.110 1256.200 ;
        RECT 1945.870 1256.000 1946.190 1256.060 ;
        RECT 1946.790 1256.000 1947.110 1256.060 ;
        RECT 1946.330 1111.020 1946.650 1111.080 ;
        RECT 1947.710 1111.020 1948.030 1111.080 ;
        RECT 1946.330 1110.880 1948.030 1111.020 ;
        RECT 1946.330 1110.820 1946.650 1110.880 ;
        RECT 1947.710 1110.820 1948.030 1110.880 ;
        RECT 1947.710 1077.020 1948.030 1077.080 ;
        RECT 1947.340 1076.880 1948.030 1077.020 ;
        RECT 1947.340 1076.400 1947.480 1076.880 ;
        RECT 1947.710 1076.820 1948.030 1076.880 ;
        RECT 1947.250 1076.140 1947.570 1076.400 ;
        RECT 1946.330 1014.460 1946.650 1014.520 ;
        RECT 1947.710 1014.460 1948.030 1014.520 ;
        RECT 1946.330 1014.320 1948.030 1014.460 ;
        RECT 1946.330 1014.260 1946.650 1014.320 ;
        RECT 1947.710 1014.260 1948.030 1014.320 ;
        RECT 1947.710 980.460 1948.030 980.520 ;
        RECT 1947.340 980.320 1948.030 980.460 ;
        RECT 1947.340 979.840 1947.480 980.320 ;
        RECT 1947.710 980.260 1948.030 980.320 ;
        RECT 1947.250 979.580 1947.570 979.840 ;
        RECT 1946.330 917.900 1946.650 917.960 ;
        RECT 1947.710 917.900 1948.030 917.960 ;
        RECT 1946.330 917.760 1948.030 917.900 ;
        RECT 1946.330 917.700 1946.650 917.760 ;
        RECT 1947.710 917.700 1948.030 917.760 ;
        RECT 1947.710 883.900 1948.030 883.960 ;
        RECT 1947.340 883.760 1948.030 883.900 ;
        RECT 1947.340 883.280 1947.480 883.760 ;
        RECT 1947.710 883.700 1948.030 883.760 ;
        RECT 1947.250 883.020 1947.570 883.280 ;
        RECT 1946.790 607.140 1947.110 607.200 ;
        RECT 1946.595 607.000 1947.110 607.140 ;
        RECT 1946.790 606.940 1947.110 607.000 ;
        RECT 1946.790 517.720 1947.110 517.780 ;
        RECT 1946.595 517.580 1947.110 517.720 ;
        RECT 1946.790 517.520 1947.110 517.580 ;
        RECT 1946.345 493.580 1946.635 493.625 ;
        RECT 1946.790 493.580 1947.110 493.640 ;
        RECT 1946.345 493.440 1947.110 493.580 ;
        RECT 1946.345 493.395 1946.635 493.440 ;
        RECT 1946.790 493.380 1947.110 493.440 ;
        RECT 1946.330 448.360 1946.650 448.420 ;
        RECT 1946.135 448.220 1946.650 448.360 ;
        RECT 1946.330 448.160 1946.650 448.220 ;
        RECT 1946.790 400.220 1947.110 400.480 ;
        RECT 1946.880 399.740 1947.020 400.220 ;
        RECT 1947.250 399.740 1947.570 399.800 ;
        RECT 1946.880 399.600 1947.570 399.740 ;
        RECT 1947.250 399.540 1947.570 399.600 ;
        RECT 1946.805 379.340 1947.095 379.385 ;
        RECT 1947.250 379.340 1947.570 379.400 ;
        RECT 1946.805 379.200 1947.570 379.340 ;
        RECT 1946.805 379.155 1947.095 379.200 ;
        RECT 1947.250 379.140 1947.570 379.200 ;
        RECT 1946.790 331.400 1947.110 331.460 ;
        RECT 1946.595 331.260 1947.110 331.400 ;
        RECT 1946.790 331.200 1947.110 331.260 ;
        RECT 1945.885 287.880 1946.175 287.925 ;
        RECT 1946.790 287.880 1947.110 287.940 ;
        RECT 1945.885 287.740 1947.110 287.880 ;
        RECT 1945.885 287.695 1946.175 287.740 ;
        RECT 1946.790 287.680 1947.110 287.740 ;
        RECT 1945.885 241.640 1946.175 241.685 ;
        RECT 1946.330 241.640 1946.650 241.700 ;
        RECT 1945.885 241.500 1946.650 241.640 ;
        RECT 1945.885 241.455 1946.175 241.500 ;
        RECT 1946.330 241.440 1946.650 241.500 ;
        RECT 1945.870 186.560 1946.190 186.620 ;
        RECT 1946.790 186.560 1947.110 186.620 ;
        RECT 1945.870 186.420 1947.110 186.560 ;
        RECT 1945.870 186.360 1946.190 186.420 ;
        RECT 1946.790 186.360 1947.110 186.420 ;
        RECT 1946.330 138.620 1946.650 138.680 ;
        RECT 1946.790 138.620 1947.110 138.680 ;
        RECT 1946.330 138.480 1947.110 138.620 ;
        RECT 1946.330 138.420 1946.650 138.480 ;
        RECT 1946.790 138.420 1947.110 138.480 ;
        RECT 1946.790 131.140 1947.110 131.200 ;
        RECT 1946.595 131.000 1947.110 131.140 ;
        RECT 1946.790 130.940 1947.110 131.000 ;
        RECT 1946.790 83.200 1947.110 83.260 ;
        RECT 1946.595 83.060 1947.110 83.200 ;
        RECT 1946.790 83.000 1947.110 83.060 ;
        RECT 1946.790 34.580 1947.110 34.640 ;
        RECT 1947.710 34.580 1948.030 34.640 ;
        RECT 1946.790 34.440 1948.030 34.580 ;
        RECT 1946.790 34.380 1947.110 34.440 ;
        RECT 1947.710 34.380 1948.030 34.440 ;
        RECT 1946.330 17.580 1946.650 17.640 ;
        RECT 1947.265 17.580 1947.555 17.625 ;
        RECT 1946.330 17.440 1947.555 17.580 ;
        RECT 1946.330 17.380 1946.650 17.440 ;
        RECT 1947.265 17.395 1947.555 17.440 ;
        RECT 1947.250 2.960 1947.570 3.020 ;
        RECT 1947.055 2.820 1947.570 2.960 ;
        RECT 1947.250 2.760 1947.570 2.820 ;
      LAYER via ;
        RECT 1946.360 1655.840 1946.620 1656.100 ;
        RECT 1947.280 1655.840 1947.540 1656.100 ;
        RECT 1947.280 1641.900 1947.540 1642.160 ;
        RECT 1947.740 1593.960 1948.000 1594.220 ;
        RECT 1946.820 1559.280 1947.080 1559.540 ;
        RECT 1947.740 1559.280 1948.000 1559.540 ;
        RECT 1945.900 1511.000 1946.160 1511.260 ;
        RECT 1946.820 1511.000 1947.080 1511.260 ;
        RECT 1947.280 1448.780 1947.540 1449.040 ;
        RECT 1946.820 1400.840 1947.080 1401.100 ;
        RECT 1947.280 1352.220 1947.540 1352.480 ;
        RECT 1946.820 1304.280 1947.080 1304.540 ;
        RECT 1945.900 1256.000 1946.160 1256.260 ;
        RECT 1946.820 1256.000 1947.080 1256.260 ;
        RECT 1946.360 1110.820 1946.620 1111.080 ;
        RECT 1947.740 1110.820 1948.000 1111.080 ;
        RECT 1947.740 1076.820 1948.000 1077.080 ;
        RECT 1947.280 1076.140 1947.540 1076.400 ;
        RECT 1946.360 1014.260 1946.620 1014.520 ;
        RECT 1947.740 1014.260 1948.000 1014.520 ;
        RECT 1947.740 980.260 1948.000 980.520 ;
        RECT 1947.280 979.580 1947.540 979.840 ;
        RECT 1946.360 917.700 1946.620 917.960 ;
        RECT 1947.740 917.700 1948.000 917.960 ;
        RECT 1947.740 883.700 1948.000 883.960 ;
        RECT 1947.280 883.020 1947.540 883.280 ;
        RECT 1946.820 606.940 1947.080 607.200 ;
        RECT 1946.820 517.520 1947.080 517.780 ;
        RECT 1946.820 493.380 1947.080 493.640 ;
        RECT 1946.360 448.160 1946.620 448.420 ;
        RECT 1946.820 400.220 1947.080 400.480 ;
        RECT 1947.280 399.540 1947.540 399.800 ;
        RECT 1947.280 379.140 1947.540 379.400 ;
        RECT 1946.820 331.200 1947.080 331.460 ;
        RECT 1946.820 287.680 1947.080 287.940 ;
        RECT 1946.360 241.440 1946.620 241.700 ;
        RECT 1945.900 186.360 1946.160 186.620 ;
        RECT 1946.820 186.360 1947.080 186.620 ;
        RECT 1946.360 138.420 1946.620 138.680 ;
        RECT 1946.820 138.420 1947.080 138.680 ;
        RECT 1946.820 130.940 1947.080 131.200 ;
        RECT 1946.820 83.000 1947.080 83.260 ;
        RECT 1946.820 34.380 1947.080 34.640 ;
        RECT 1947.740 34.380 1948.000 34.640 ;
        RECT 1946.360 17.380 1946.620 17.640 ;
        RECT 1947.280 2.760 1947.540 3.020 ;
      LAYER met2 ;
        RECT 1950.885 1701.090 1951.165 1704.000 ;
        RECT 1948.720 1700.950 1951.165 1701.090 ;
        RECT 1948.720 1656.210 1948.860 1700.950 ;
        RECT 1950.885 1700.000 1951.165 1700.950 ;
        RECT 1946.420 1656.130 1948.860 1656.210 ;
        RECT 1946.360 1656.070 1948.860 1656.130 ;
        RECT 1946.360 1655.810 1946.620 1656.070 ;
        RECT 1947.280 1655.810 1947.540 1656.070 ;
        RECT 1947.340 1642.190 1947.480 1655.810 ;
        RECT 1947.280 1641.870 1947.540 1642.190 ;
        RECT 1947.740 1593.930 1948.000 1594.250 ;
        RECT 1947.800 1559.570 1947.940 1593.930 ;
        RECT 1946.820 1559.250 1947.080 1559.570 ;
        RECT 1947.740 1559.250 1948.000 1559.570 ;
        RECT 1946.880 1511.290 1947.020 1559.250 ;
        RECT 1945.900 1510.970 1946.160 1511.290 ;
        RECT 1946.820 1510.970 1947.080 1511.290 ;
        RECT 1945.960 1510.690 1946.100 1510.970 ;
        RECT 1945.960 1510.550 1946.560 1510.690 ;
        RECT 1946.420 1463.090 1946.560 1510.550 ;
        RECT 1946.420 1462.950 1947.480 1463.090 ;
        RECT 1947.340 1449.070 1947.480 1462.950 ;
        RECT 1947.280 1448.750 1947.540 1449.070 ;
        RECT 1946.820 1400.810 1947.080 1401.130 ;
        RECT 1946.880 1366.530 1947.020 1400.810 ;
        RECT 1946.880 1366.390 1947.480 1366.530 ;
        RECT 1947.340 1352.510 1947.480 1366.390 ;
        RECT 1947.280 1352.190 1947.540 1352.510 ;
        RECT 1946.820 1304.250 1947.080 1304.570 ;
        RECT 1946.880 1256.290 1947.020 1304.250 ;
        RECT 1945.900 1255.970 1946.160 1256.290 ;
        RECT 1946.820 1255.970 1947.080 1256.290 ;
        RECT 1945.960 1221.010 1946.100 1255.970 ;
        RECT 1945.960 1220.870 1946.560 1221.010 ;
        RECT 1946.420 1173.410 1946.560 1220.870 ;
        RECT 1946.420 1173.270 1947.480 1173.410 ;
        RECT 1947.340 1159.245 1947.480 1173.270 ;
        RECT 1946.350 1158.875 1946.630 1159.245 ;
        RECT 1947.270 1158.875 1947.550 1159.245 ;
        RECT 1946.420 1111.110 1946.560 1158.875 ;
        RECT 1946.360 1110.790 1946.620 1111.110 ;
        RECT 1947.740 1110.790 1948.000 1111.110 ;
        RECT 1947.800 1077.110 1947.940 1110.790 ;
        RECT 1947.740 1076.790 1948.000 1077.110 ;
        RECT 1947.280 1076.110 1947.540 1076.430 ;
        RECT 1947.340 1062.685 1947.480 1076.110 ;
        RECT 1946.350 1062.315 1946.630 1062.685 ;
        RECT 1947.270 1062.315 1947.550 1062.685 ;
        RECT 1946.420 1014.550 1946.560 1062.315 ;
        RECT 1946.360 1014.230 1946.620 1014.550 ;
        RECT 1947.740 1014.230 1948.000 1014.550 ;
        RECT 1947.800 980.550 1947.940 1014.230 ;
        RECT 1947.740 980.230 1948.000 980.550 ;
        RECT 1947.280 979.550 1947.540 979.870 ;
        RECT 1947.340 966.125 1947.480 979.550 ;
        RECT 1946.350 965.755 1946.630 966.125 ;
        RECT 1947.270 965.755 1947.550 966.125 ;
        RECT 1946.420 917.990 1946.560 965.755 ;
        RECT 1946.360 917.670 1946.620 917.990 ;
        RECT 1947.740 917.670 1948.000 917.990 ;
        RECT 1947.800 883.990 1947.940 917.670 ;
        RECT 1947.740 883.670 1948.000 883.990 ;
        RECT 1947.280 882.990 1947.540 883.310 ;
        RECT 1947.340 614.450 1947.480 882.990 ;
        RECT 1946.880 614.310 1947.480 614.450 ;
        RECT 1946.880 607.230 1947.020 614.310 ;
        RECT 1946.820 606.910 1947.080 607.230 ;
        RECT 1946.820 517.490 1947.080 517.810 ;
        RECT 1946.880 493.670 1947.020 517.490 ;
        RECT 1946.820 493.350 1947.080 493.670 ;
        RECT 1946.360 448.130 1946.620 448.450 ;
        RECT 1946.420 434.930 1946.560 448.130 ;
        RECT 1946.420 434.790 1947.020 434.930 ;
        RECT 1946.880 400.510 1947.020 434.790 ;
        RECT 1946.820 400.190 1947.080 400.510 ;
        RECT 1947.280 399.510 1947.540 399.830 ;
        RECT 1947.340 379.430 1947.480 399.510 ;
        RECT 1947.280 379.110 1947.540 379.430 ;
        RECT 1946.820 331.170 1947.080 331.490 ;
        RECT 1946.880 287.970 1947.020 331.170 ;
        RECT 1946.820 287.650 1947.080 287.970 ;
        RECT 1946.360 241.410 1946.620 241.730 ;
        RECT 1946.420 210.530 1946.560 241.410 ;
        RECT 1945.960 210.390 1946.560 210.530 ;
        RECT 1945.960 186.650 1946.100 210.390 ;
        RECT 1945.900 186.330 1946.160 186.650 ;
        RECT 1946.820 186.330 1947.080 186.650 ;
        RECT 1946.880 158.170 1947.020 186.330 ;
        RECT 1946.420 158.030 1947.020 158.170 ;
        RECT 1946.420 138.710 1946.560 158.030 ;
        RECT 1946.360 138.390 1946.620 138.710 ;
        RECT 1946.820 138.390 1947.080 138.710 ;
        RECT 1946.880 131.230 1947.020 138.390 ;
        RECT 1946.820 130.910 1947.080 131.230 ;
        RECT 1946.820 82.970 1947.080 83.290 ;
        RECT 1946.880 82.805 1947.020 82.970 ;
        RECT 1946.810 82.435 1947.090 82.805 ;
        RECT 1947.730 82.435 1948.010 82.805 ;
        RECT 1946.880 34.670 1947.020 34.825 ;
        RECT 1947.800 34.670 1947.940 82.435 ;
        RECT 1946.820 34.410 1947.080 34.670 ;
        RECT 1946.420 34.350 1947.080 34.410 ;
        RECT 1947.740 34.350 1948.000 34.670 ;
        RECT 1946.420 34.270 1947.020 34.350 ;
        RECT 1946.420 17.670 1946.560 34.270 ;
        RECT 1946.360 17.350 1946.620 17.670 ;
        RECT 1947.280 2.730 1947.540 3.050 ;
        RECT 1947.340 2.400 1947.480 2.730 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
      LAYER via2 ;
        RECT 1946.350 1158.920 1946.630 1159.200 ;
        RECT 1947.270 1158.920 1947.550 1159.200 ;
        RECT 1946.350 1062.360 1946.630 1062.640 ;
        RECT 1947.270 1062.360 1947.550 1062.640 ;
        RECT 1946.350 965.800 1946.630 966.080 ;
        RECT 1947.270 965.800 1947.550 966.080 ;
        RECT 1946.810 82.480 1947.090 82.760 ;
        RECT 1947.730 82.480 1948.010 82.760 ;
      LAYER met3 ;
        RECT 1946.325 1159.210 1946.655 1159.225 ;
        RECT 1947.245 1159.210 1947.575 1159.225 ;
        RECT 1946.325 1158.910 1947.575 1159.210 ;
        RECT 1946.325 1158.895 1946.655 1158.910 ;
        RECT 1947.245 1158.895 1947.575 1158.910 ;
        RECT 1946.325 1062.650 1946.655 1062.665 ;
        RECT 1947.245 1062.650 1947.575 1062.665 ;
        RECT 1946.325 1062.350 1947.575 1062.650 ;
        RECT 1946.325 1062.335 1946.655 1062.350 ;
        RECT 1947.245 1062.335 1947.575 1062.350 ;
        RECT 1946.325 966.090 1946.655 966.105 ;
        RECT 1947.245 966.090 1947.575 966.105 ;
        RECT 1946.325 965.790 1947.575 966.090 ;
        RECT 1946.325 965.775 1946.655 965.790 ;
        RECT 1947.245 965.775 1947.575 965.790 ;
        RECT 1946.785 82.770 1947.115 82.785 ;
        RECT 1947.705 82.770 1948.035 82.785 ;
        RECT 1946.785 82.470 1948.035 82.770 ;
        RECT 1946.785 82.455 1947.115 82.470 ;
        RECT 1947.705 82.455 1948.035 82.470 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1958.245 1700.410 1958.525 1704.000 ;
        RECT 1958.245 1700.270 1959.440 1700.410 ;
        RECT 1958.245 1700.000 1958.525 1700.270 ;
        RECT 1959.300 1684.090 1959.440 1700.270 ;
        RECT 1959.300 1683.950 1960.820 1684.090 ;
        RECT 1960.680 7.210 1960.820 1683.950 ;
        RECT 1960.680 7.070 1965.420 7.210 ;
        RECT 1965.280 2.400 1965.420 7.070 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1965.650 20.300 1965.970 20.360 ;
        RECT 1983.130 20.300 1983.450 20.360 ;
        RECT 1965.650 20.160 1983.450 20.300 ;
        RECT 1965.650 20.100 1965.970 20.160 ;
        RECT 1983.130 20.100 1983.450 20.160 ;
      LAYER via ;
        RECT 1965.680 20.100 1965.940 20.360 ;
        RECT 1983.160 20.100 1983.420 20.360 ;
      LAYER met2 ;
        RECT 1965.605 1700.000 1965.885 1704.000 ;
        RECT 1965.740 20.390 1965.880 1700.000 ;
        RECT 1965.680 20.070 1965.940 20.390 ;
        RECT 1983.160 20.070 1983.420 20.390 ;
        RECT 1983.220 2.400 1983.360 20.070 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1972.550 16.560 1972.870 16.620 ;
        RECT 2001.070 16.560 2001.390 16.620 ;
        RECT 1972.550 16.420 2001.390 16.560 ;
        RECT 1972.550 16.360 1972.870 16.420 ;
        RECT 2001.070 16.360 2001.390 16.420 ;
      LAYER via ;
        RECT 1972.580 16.360 1972.840 16.620 ;
        RECT 2001.100 16.360 2001.360 16.620 ;
      LAYER met2 ;
        RECT 1972.965 1700.410 1973.245 1704.000 ;
        RECT 1972.640 1700.270 1973.245 1700.410 ;
        RECT 1972.640 16.650 1972.780 1700.270 ;
        RECT 1972.965 1700.000 1973.245 1700.270 ;
        RECT 1972.580 16.330 1972.840 16.650 ;
        RECT 2001.100 16.330 2001.360 16.650 ;
        RECT 2001.160 2.400 2001.300 16.330 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1980.370 1684.260 1980.690 1684.320 ;
        RECT 1990.490 1684.260 1990.810 1684.320 ;
        RECT 1980.370 1684.120 1990.810 1684.260 ;
        RECT 1980.370 1684.060 1980.690 1684.120 ;
        RECT 1990.490 1684.060 1990.810 1684.120 ;
        RECT 1990.490 20.640 1990.810 20.700 ;
        RECT 2018.550 20.640 2018.870 20.700 ;
        RECT 1990.490 20.500 2018.870 20.640 ;
        RECT 1990.490 20.440 1990.810 20.500 ;
        RECT 2018.550 20.440 2018.870 20.500 ;
      LAYER via ;
        RECT 1980.400 1684.060 1980.660 1684.320 ;
        RECT 1990.520 1684.060 1990.780 1684.320 ;
        RECT 1990.520 20.440 1990.780 20.700 ;
        RECT 2018.580 20.440 2018.840 20.700 ;
      LAYER met2 ;
        RECT 1980.325 1700.000 1980.605 1704.000 ;
        RECT 1980.460 1684.350 1980.600 1700.000 ;
        RECT 1980.400 1684.030 1980.660 1684.350 ;
        RECT 1990.520 1684.030 1990.780 1684.350 ;
        RECT 1990.580 20.730 1990.720 1684.030 ;
        RECT 1990.520 20.410 1990.780 20.730 ;
        RECT 2018.580 20.410 2018.840 20.730 ;
        RECT 2018.640 2.400 2018.780 20.410 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1987.270 1689.360 1987.590 1689.420 ;
        RECT 1997.390 1689.360 1997.710 1689.420 ;
        RECT 1987.270 1689.220 1997.710 1689.360 ;
        RECT 1987.270 1689.160 1987.590 1689.220 ;
        RECT 1997.390 1689.160 1997.710 1689.220 ;
        RECT 1997.390 19.280 1997.710 19.340 ;
        RECT 2036.490 19.280 2036.810 19.340 ;
        RECT 1997.390 19.140 2036.810 19.280 ;
        RECT 1997.390 19.080 1997.710 19.140 ;
        RECT 2036.490 19.080 2036.810 19.140 ;
      LAYER via ;
        RECT 1987.300 1689.160 1987.560 1689.420 ;
        RECT 1997.420 1689.160 1997.680 1689.420 ;
        RECT 1997.420 19.080 1997.680 19.340 ;
        RECT 2036.520 19.080 2036.780 19.340 ;
      LAYER met2 ;
        RECT 1987.225 1700.000 1987.505 1704.000 ;
        RECT 1987.360 1689.450 1987.500 1700.000 ;
        RECT 1987.300 1689.130 1987.560 1689.450 ;
        RECT 1997.420 1689.130 1997.680 1689.450 ;
        RECT 1997.480 19.370 1997.620 1689.130 ;
        RECT 1997.420 19.050 1997.680 19.370 ;
        RECT 2036.520 19.050 2036.780 19.370 ;
        RECT 2036.580 2.400 2036.720 19.050 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1994.630 1684.940 1994.950 1685.000 ;
        RECT 2018.090 1684.940 2018.410 1685.000 ;
        RECT 1994.630 1684.800 2018.410 1684.940 ;
        RECT 1994.630 1684.740 1994.950 1684.800 ;
        RECT 2018.090 1684.740 2018.410 1684.800 ;
        RECT 2018.090 16.560 2018.410 16.620 ;
        RECT 2054.430 16.560 2054.750 16.620 ;
        RECT 2018.090 16.420 2054.750 16.560 ;
        RECT 2018.090 16.360 2018.410 16.420 ;
        RECT 2054.430 16.360 2054.750 16.420 ;
      LAYER via ;
        RECT 1994.660 1684.740 1994.920 1685.000 ;
        RECT 2018.120 1684.740 2018.380 1685.000 ;
        RECT 2018.120 16.360 2018.380 16.620 ;
        RECT 2054.460 16.360 2054.720 16.620 ;
      LAYER met2 ;
        RECT 1994.585 1700.000 1994.865 1704.000 ;
        RECT 1994.720 1685.030 1994.860 1700.000 ;
        RECT 1994.660 1684.710 1994.920 1685.030 ;
        RECT 2018.120 1684.710 2018.380 1685.030 ;
        RECT 2018.180 16.650 2018.320 1684.710 ;
        RECT 2018.120 16.330 2018.380 16.650 ;
        RECT 2054.460 16.330 2054.720 16.650 ;
        RECT 2054.520 2.400 2054.660 16.330 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 772.410 49.200 772.730 49.260 ;
        RECT 1464.250 49.200 1464.570 49.260 ;
        RECT 772.410 49.060 1464.570 49.200 ;
        RECT 772.410 49.000 772.730 49.060 ;
        RECT 1464.250 49.000 1464.570 49.060 ;
      LAYER via ;
        RECT 772.440 49.000 772.700 49.260 ;
        RECT 1464.280 49.000 1464.540 49.260 ;
      LAYER met2 ;
        RECT 1465.585 1700.410 1465.865 1704.000 ;
        RECT 1464.340 1700.270 1465.865 1700.410 ;
        RECT 1464.340 49.290 1464.480 1700.270 ;
        RECT 1465.585 1700.000 1465.865 1700.270 ;
        RECT 772.440 48.970 772.700 49.290 ;
        RECT 1464.280 48.970 1464.540 49.290 ;
        RECT 772.500 17.410 772.640 48.970 ;
        RECT 769.740 17.270 772.640 17.410 ;
        RECT 769.740 2.400 769.880 17.270 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2001.990 1687.660 2002.310 1687.720 ;
        RECT 2031.890 1687.660 2032.210 1687.720 ;
        RECT 2001.990 1687.520 2032.210 1687.660 ;
        RECT 2001.990 1687.460 2002.310 1687.520 ;
        RECT 2031.890 1687.460 2032.210 1687.520 ;
        RECT 2031.890 19.960 2032.210 20.020 ;
        RECT 2072.370 19.960 2072.690 20.020 ;
        RECT 2031.890 19.820 2072.690 19.960 ;
        RECT 2031.890 19.760 2032.210 19.820 ;
        RECT 2072.370 19.760 2072.690 19.820 ;
      LAYER via ;
        RECT 2002.020 1687.460 2002.280 1687.720 ;
        RECT 2031.920 1687.460 2032.180 1687.720 ;
        RECT 2031.920 19.760 2032.180 20.020 ;
        RECT 2072.400 19.760 2072.660 20.020 ;
      LAYER met2 ;
        RECT 2001.945 1700.000 2002.225 1704.000 ;
        RECT 2002.080 1687.750 2002.220 1700.000 ;
        RECT 2002.020 1687.430 2002.280 1687.750 ;
        RECT 2031.920 1687.430 2032.180 1687.750 ;
        RECT 2031.980 20.050 2032.120 1687.430 ;
        RECT 2031.920 19.730 2032.180 20.050 ;
        RECT 2072.400 19.730 2072.660 20.050 ;
        RECT 2072.460 2.400 2072.600 19.730 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2009.350 1689.020 2009.670 1689.080 ;
        RECT 2084.790 1689.020 2085.110 1689.080 ;
        RECT 2009.350 1688.880 2085.110 1689.020 ;
        RECT 2009.350 1688.820 2009.670 1688.880 ;
        RECT 2084.790 1688.820 2085.110 1688.880 ;
      LAYER via ;
        RECT 2009.380 1688.820 2009.640 1689.080 ;
        RECT 2084.820 1688.820 2085.080 1689.080 ;
      LAYER met2 ;
        RECT 2009.305 1700.000 2009.585 1704.000 ;
        RECT 2009.440 1689.110 2009.580 1700.000 ;
        RECT 2009.380 1688.790 2009.640 1689.110 ;
        RECT 2084.820 1688.790 2085.080 1689.110 ;
        RECT 2084.880 16.730 2085.020 1688.790 ;
        RECT 2084.880 16.590 2090.080 16.730 ;
        RECT 2089.940 2.400 2090.080 16.590 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2062.785 1688.185 2062.955 1690.055 ;
        RECT 2067.385 1685.125 2067.555 1688.355 ;
      LAYER mcon ;
        RECT 2062.785 1689.885 2062.955 1690.055 ;
        RECT 2067.385 1688.185 2067.555 1688.355 ;
      LAYER met1 ;
        RECT 2016.710 1690.040 2017.030 1690.100 ;
        RECT 2062.725 1690.040 2063.015 1690.085 ;
        RECT 2016.710 1689.900 2063.015 1690.040 ;
        RECT 2016.710 1689.840 2017.030 1689.900 ;
        RECT 2062.725 1689.855 2063.015 1689.900 ;
        RECT 2062.725 1688.340 2063.015 1688.385 ;
        RECT 2067.325 1688.340 2067.615 1688.385 ;
        RECT 2062.725 1688.200 2067.615 1688.340 ;
        RECT 2062.725 1688.155 2063.015 1688.200 ;
        RECT 2067.325 1688.155 2067.615 1688.200 ;
        RECT 2067.325 1685.280 2067.615 1685.325 ;
        RECT 2105.490 1685.280 2105.810 1685.340 ;
        RECT 2067.325 1685.140 2105.810 1685.280 ;
        RECT 2067.325 1685.095 2067.615 1685.140 ;
        RECT 2105.490 1685.080 2105.810 1685.140 ;
      LAYER via ;
        RECT 2016.740 1689.840 2017.000 1690.100 ;
        RECT 2105.520 1685.080 2105.780 1685.340 ;
      LAYER met2 ;
        RECT 2016.665 1700.000 2016.945 1704.000 ;
        RECT 2016.800 1690.130 2016.940 1700.000 ;
        RECT 2016.740 1689.810 2017.000 1690.130 ;
        RECT 2105.520 1685.050 2105.780 1685.370 ;
        RECT 2105.580 16.730 2105.720 1685.050 ;
        RECT 2105.580 16.590 2108.020 16.730 ;
        RECT 2107.880 2.400 2108.020 16.590 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2077.505 1685.805 2077.675 1688.015 ;
      LAYER mcon ;
        RECT 2077.505 1687.845 2077.675 1688.015 ;
      LAYER met1 ;
        RECT 2024.070 1688.000 2024.390 1688.060 ;
        RECT 2077.445 1688.000 2077.735 1688.045 ;
        RECT 2024.070 1687.860 2077.735 1688.000 ;
        RECT 2024.070 1687.800 2024.390 1687.860 ;
        RECT 2077.445 1687.815 2077.735 1687.860 ;
        RECT 2077.445 1685.960 2077.735 1686.005 ;
        RECT 2121.590 1685.960 2121.910 1686.020 ;
        RECT 2077.445 1685.820 2121.910 1685.960 ;
        RECT 2077.445 1685.775 2077.735 1685.820 ;
        RECT 2121.590 1685.760 2121.910 1685.820 ;
        RECT 2121.590 17.240 2121.910 17.300 ;
        RECT 2125.730 17.240 2126.050 17.300 ;
        RECT 2121.590 17.100 2126.050 17.240 ;
        RECT 2121.590 17.040 2121.910 17.100 ;
        RECT 2125.730 17.040 2126.050 17.100 ;
      LAYER via ;
        RECT 2024.100 1687.800 2024.360 1688.060 ;
        RECT 2121.620 1685.760 2121.880 1686.020 ;
        RECT 2121.620 17.040 2121.880 17.300 ;
        RECT 2125.760 17.040 2126.020 17.300 ;
      LAYER met2 ;
        RECT 2024.025 1700.000 2024.305 1704.000 ;
        RECT 2024.160 1688.090 2024.300 1700.000 ;
        RECT 2024.100 1687.770 2024.360 1688.090 ;
        RECT 2121.620 1685.730 2121.880 1686.050 ;
        RECT 2121.680 17.330 2121.820 1685.730 ;
        RECT 2121.620 17.010 2121.880 17.330 ;
        RECT 2125.760 17.010 2126.020 17.330 ;
        RECT 2125.820 2.400 2125.960 17.010 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2031.430 1685.620 2031.750 1685.680 ;
        RECT 2059.490 1685.620 2059.810 1685.680 ;
        RECT 2031.430 1685.480 2059.810 1685.620 ;
        RECT 2031.430 1685.420 2031.750 1685.480 ;
        RECT 2059.490 1685.420 2059.810 1685.480 ;
        RECT 2059.490 15.540 2059.810 15.600 ;
        RECT 2143.670 15.540 2143.990 15.600 ;
        RECT 2059.490 15.400 2143.990 15.540 ;
        RECT 2059.490 15.340 2059.810 15.400 ;
        RECT 2143.670 15.340 2143.990 15.400 ;
      LAYER via ;
        RECT 2031.460 1685.420 2031.720 1685.680 ;
        RECT 2059.520 1685.420 2059.780 1685.680 ;
        RECT 2059.520 15.340 2059.780 15.600 ;
        RECT 2143.700 15.340 2143.960 15.600 ;
      LAYER met2 ;
        RECT 2031.385 1700.000 2031.665 1704.000 ;
        RECT 2031.520 1685.710 2031.660 1700.000 ;
        RECT 2031.460 1685.390 2031.720 1685.710 ;
        RECT 2059.520 1685.390 2059.780 1685.710 ;
        RECT 2059.580 15.630 2059.720 1685.390 ;
        RECT 2059.520 15.310 2059.780 15.630 ;
        RECT 2143.700 15.310 2143.960 15.630 ;
        RECT 2143.760 2.400 2143.900 15.310 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2038.790 1684.940 2039.110 1685.000 ;
        RECT 2038.790 1684.800 2056.500 1684.940 ;
        RECT 2038.790 1684.740 2039.110 1684.800 ;
        RECT 2056.360 1684.600 2056.500 1684.800 ;
        RECT 2066.390 1684.600 2066.710 1684.660 ;
        RECT 2056.360 1684.460 2066.710 1684.600 ;
        RECT 2066.390 1684.400 2066.710 1684.460 ;
        RECT 2066.390 18.940 2066.710 19.000 ;
        RECT 2067.310 18.940 2067.630 19.000 ;
        RECT 2066.390 18.800 2067.630 18.940 ;
        RECT 2066.390 18.740 2066.710 18.800 ;
        RECT 2067.310 18.740 2067.630 18.800 ;
        RECT 2067.310 14.860 2067.630 14.920 ;
        RECT 2161.610 14.860 2161.930 14.920 ;
        RECT 2067.310 14.720 2161.930 14.860 ;
        RECT 2067.310 14.660 2067.630 14.720 ;
        RECT 2161.610 14.660 2161.930 14.720 ;
      LAYER via ;
        RECT 2038.820 1684.740 2039.080 1685.000 ;
        RECT 2066.420 1684.400 2066.680 1684.660 ;
        RECT 2066.420 18.740 2066.680 19.000 ;
        RECT 2067.340 18.740 2067.600 19.000 ;
        RECT 2067.340 14.660 2067.600 14.920 ;
        RECT 2161.640 14.660 2161.900 14.920 ;
      LAYER met2 ;
        RECT 2038.745 1700.000 2039.025 1704.000 ;
        RECT 2038.880 1685.030 2039.020 1700.000 ;
        RECT 2038.820 1684.710 2039.080 1685.030 ;
        RECT 2066.420 1684.370 2066.680 1684.690 ;
        RECT 2066.480 19.030 2066.620 1684.370 ;
        RECT 2066.420 18.710 2066.680 19.030 ;
        RECT 2067.340 18.710 2067.600 19.030 ;
        RECT 2067.400 14.950 2067.540 18.710 ;
        RECT 2067.340 14.630 2067.600 14.950 ;
        RECT 2161.640 14.630 2161.900 14.950 ;
        RECT 2161.700 2.400 2161.840 14.630 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2140.985 14.025 2141.155 15.215 ;
      LAYER mcon ;
        RECT 2140.985 15.045 2141.155 15.215 ;
      LAYER met1 ;
        RECT 2046.150 1689.700 2046.470 1689.760 ;
        RECT 2080.190 1689.700 2080.510 1689.760 ;
        RECT 2046.150 1689.560 2080.510 1689.700 ;
        RECT 2046.150 1689.500 2046.470 1689.560 ;
        RECT 2080.190 1689.500 2080.510 1689.560 ;
        RECT 2140.925 15.200 2141.215 15.245 ;
        RECT 2179.090 15.200 2179.410 15.260 ;
        RECT 2140.925 15.060 2179.410 15.200 ;
        RECT 2140.925 15.015 2141.215 15.060 ;
        RECT 2179.090 15.000 2179.410 15.060 ;
        RECT 2080.190 14.180 2080.510 14.240 ;
        RECT 2140.925 14.180 2141.215 14.225 ;
        RECT 2080.190 14.040 2141.215 14.180 ;
        RECT 2080.190 13.980 2080.510 14.040 ;
        RECT 2140.925 13.995 2141.215 14.040 ;
      LAYER via ;
        RECT 2046.180 1689.500 2046.440 1689.760 ;
        RECT 2080.220 1689.500 2080.480 1689.760 ;
        RECT 2179.120 15.000 2179.380 15.260 ;
        RECT 2080.220 13.980 2080.480 14.240 ;
      LAYER met2 ;
        RECT 2046.105 1700.000 2046.385 1704.000 ;
        RECT 2046.240 1689.790 2046.380 1700.000 ;
        RECT 2046.180 1689.470 2046.440 1689.790 ;
        RECT 2080.220 1689.470 2080.480 1689.790 ;
        RECT 2080.280 14.270 2080.420 1689.470 ;
        RECT 2179.120 14.970 2179.380 15.290 ;
        RECT 2080.220 13.950 2080.480 14.270 ;
        RECT 2179.180 2.400 2179.320 14.970 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2055.350 20.300 2055.670 20.360 ;
        RECT 2197.030 20.300 2197.350 20.360 ;
        RECT 2055.350 20.160 2197.350 20.300 ;
        RECT 2055.350 20.100 2055.670 20.160 ;
        RECT 2197.030 20.100 2197.350 20.160 ;
      LAYER via ;
        RECT 2055.380 20.100 2055.640 20.360 ;
        RECT 2197.060 20.100 2197.320 20.360 ;
      LAYER met2 ;
        RECT 2053.465 1700.410 2053.745 1704.000 ;
        RECT 2053.465 1700.270 2055.580 1700.410 ;
        RECT 2053.465 1700.000 2053.745 1700.270 ;
        RECT 2055.440 20.390 2055.580 1700.270 ;
        RECT 2055.380 20.070 2055.640 20.390 ;
        RECT 2197.060 20.070 2197.320 20.390 ;
        RECT 2197.120 2.400 2197.260 20.070 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2062.710 19.280 2063.030 19.340 ;
        RECT 2214.970 19.280 2215.290 19.340 ;
        RECT 2062.710 19.140 2215.290 19.280 ;
        RECT 2062.710 19.080 2063.030 19.140 ;
        RECT 2214.970 19.080 2215.290 19.140 ;
      LAYER via ;
        RECT 2062.740 19.080 2063.000 19.340 ;
        RECT 2215.000 19.080 2215.260 19.340 ;
      LAYER met2 ;
        RECT 2060.825 1700.410 2061.105 1704.000 ;
        RECT 2060.825 1700.270 2062.940 1700.410 ;
        RECT 2060.825 1700.000 2061.105 1700.270 ;
        RECT 2062.800 19.370 2062.940 1700.270 ;
        RECT 2062.740 19.050 2063.000 19.370 ;
        RECT 2215.000 19.050 2215.260 19.370 ;
        RECT 2215.060 2.400 2215.200 19.050 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2135.005 18.105 2135.175 19.975 ;
      LAYER mcon ;
        RECT 2135.005 19.805 2135.175 19.975 ;
      LAYER met1 ;
        RECT 2068.230 1689.360 2068.550 1689.420 ;
        RECT 2087.090 1689.360 2087.410 1689.420 ;
        RECT 2068.230 1689.220 2087.410 1689.360 ;
        RECT 2068.230 1689.160 2068.550 1689.220 ;
        RECT 2087.090 1689.160 2087.410 1689.220 ;
        RECT 2134.945 19.960 2135.235 20.005 ;
        RECT 2232.910 19.960 2233.230 20.020 ;
        RECT 2134.945 19.820 2233.230 19.960 ;
        RECT 2134.945 19.775 2135.235 19.820 ;
        RECT 2232.910 19.760 2233.230 19.820 ;
        RECT 2087.090 18.260 2087.410 18.320 ;
        RECT 2134.945 18.260 2135.235 18.305 ;
        RECT 2087.090 18.120 2135.235 18.260 ;
        RECT 2087.090 18.060 2087.410 18.120 ;
        RECT 2134.945 18.075 2135.235 18.120 ;
      LAYER via ;
        RECT 2068.260 1689.160 2068.520 1689.420 ;
        RECT 2087.120 1689.160 2087.380 1689.420 ;
        RECT 2232.940 19.760 2233.200 20.020 ;
        RECT 2087.120 18.060 2087.380 18.320 ;
      LAYER met2 ;
        RECT 2068.185 1700.000 2068.465 1704.000 ;
        RECT 2068.320 1689.450 2068.460 1700.000 ;
        RECT 2068.260 1689.130 2068.520 1689.450 ;
        RECT 2087.120 1689.130 2087.380 1689.450 ;
        RECT 2087.180 18.350 2087.320 1689.130 ;
        RECT 2232.940 19.730 2233.200 20.050 ;
        RECT 2087.120 18.030 2087.380 18.350 ;
        RECT 2233.000 2.400 2233.140 19.730 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 48.860 793.430 48.920 ;
        RECT 1470.230 48.860 1470.550 48.920 ;
        RECT 793.110 48.720 1470.550 48.860 ;
        RECT 793.110 48.660 793.430 48.720 ;
        RECT 1470.230 48.660 1470.550 48.720 ;
      LAYER via ;
        RECT 793.140 48.660 793.400 48.920 ;
        RECT 1470.260 48.660 1470.520 48.920 ;
      LAYER met2 ;
        RECT 1472.945 1700.410 1473.225 1704.000 ;
        RECT 1471.240 1700.270 1473.225 1700.410 ;
        RECT 1471.240 1678.480 1471.380 1700.270 ;
        RECT 1472.945 1700.000 1473.225 1700.270 ;
        RECT 1470.320 1678.340 1471.380 1678.480 ;
        RECT 1470.320 48.950 1470.460 1678.340 ;
        RECT 793.140 48.630 793.400 48.950 ;
        RECT 1470.260 48.630 1470.520 48.950 ;
        RECT 793.200 17.410 793.340 48.630 ;
        RECT 787.680 17.270 793.340 17.410 ;
        RECT 787.680 2.400 787.820 17.270 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2075.590 1690.040 2075.910 1690.100 ;
        RECT 2101.350 1690.040 2101.670 1690.100 ;
        RECT 2075.590 1689.900 2101.670 1690.040 ;
        RECT 2075.590 1689.840 2075.910 1689.900 ;
        RECT 2101.350 1689.840 2101.670 1689.900 ;
        RECT 2101.350 19.620 2101.670 19.680 ;
        RECT 2250.850 19.620 2251.170 19.680 ;
        RECT 2101.350 19.480 2251.170 19.620 ;
        RECT 2101.350 19.420 2101.670 19.480 ;
        RECT 2250.850 19.420 2251.170 19.480 ;
      LAYER via ;
        RECT 2075.620 1689.840 2075.880 1690.100 ;
        RECT 2101.380 1689.840 2101.640 1690.100 ;
        RECT 2101.380 19.420 2101.640 19.680 ;
        RECT 2250.880 19.420 2251.140 19.680 ;
      LAYER met2 ;
        RECT 2075.545 1700.000 2075.825 1704.000 ;
        RECT 2075.680 1690.130 2075.820 1700.000 ;
        RECT 2075.620 1689.810 2075.880 1690.130 ;
        RECT 2101.380 1689.810 2101.640 1690.130 ;
        RECT 2101.440 19.710 2101.580 1689.810 ;
        RECT 2101.380 19.390 2101.640 19.710 ;
        RECT 2250.880 19.390 2251.140 19.710 ;
        RECT 2250.940 2.400 2251.080 19.390 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2111.545 14.365 2111.715 18.615 ;
        RECT 2159.385 13.685 2159.555 18.615 ;
      LAYER mcon ;
        RECT 2111.545 18.445 2111.715 18.615 ;
        RECT 2159.385 18.445 2159.555 18.615 ;
      LAYER met1 ;
        RECT 2082.950 1689.700 2083.270 1689.760 ;
        RECT 2107.790 1689.700 2108.110 1689.760 ;
        RECT 2082.950 1689.560 2108.110 1689.700 ;
        RECT 2082.950 1689.500 2083.270 1689.560 ;
        RECT 2107.790 1689.500 2108.110 1689.560 ;
        RECT 2268.330 19.280 2268.650 19.340 ;
        RECT 2227.480 19.140 2268.650 19.280 ;
        RECT 2107.790 18.600 2108.110 18.660 ;
        RECT 2111.485 18.600 2111.775 18.645 ;
        RECT 2107.790 18.460 2111.775 18.600 ;
        RECT 2107.790 18.400 2108.110 18.460 ;
        RECT 2111.485 18.415 2111.775 18.460 ;
        RECT 2159.325 18.600 2159.615 18.645 ;
        RECT 2227.480 18.600 2227.620 19.140 ;
        RECT 2268.330 19.080 2268.650 19.140 ;
        RECT 2159.325 18.460 2227.620 18.600 ;
        RECT 2159.325 18.415 2159.615 18.460 ;
        RECT 2111.485 14.520 2111.775 14.565 ;
        RECT 2111.485 14.380 2142.060 14.520 ;
        RECT 2111.485 14.335 2111.775 14.380 ;
        RECT 2141.920 13.840 2142.060 14.380 ;
        RECT 2159.325 13.840 2159.615 13.885 ;
        RECT 2141.920 13.700 2159.615 13.840 ;
        RECT 2159.325 13.655 2159.615 13.700 ;
      LAYER via ;
        RECT 2082.980 1689.500 2083.240 1689.760 ;
        RECT 2107.820 1689.500 2108.080 1689.760 ;
        RECT 2107.820 18.400 2108.080 18.660 ;
        RECT 2268.360 19.080 2268.620 19.340 ;
      LAYER met2 ;
        RECT 2082.905 1700.000 2083.185 1704.000 ;
        RECT 2083.040 1689.790 2083.180 1700.000 ;
        RECT 2082.980 1689.470 2083.240 1689.790 ;
        RECT 2107.820 1689.470 2108.080 1689.790 ;
        RECT 2107.880 18.690 2108.020 1689.470 ;
        RECT 2268.360 19.050 2268.620 19.370 ;
        RECT 2107.820 18.370 2108.080 18.690 ;
        RECT 2268.420 2.400 2268.560 19.050 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2090.310 17.580 2090.630 17.640 ;
        RECT 2286.270 17.580 2286.590 17.640 ;
        RECT 2090.310 17.440 2286.590 17.580 ;
        RECT 2090.310 17.380 2090.630 17.440 ;
        RECT 2286.270 17.380 2286.590 17.440 ;
      LAYER via ;
        RECT 2090.340 17.380 2090.600 17.640 ;
        RECT 2286.300 17.380 2286.560 17.640 ;
      LAYER met2 ;
        RECT 2090.265 1700.000 2090.545 1704.000 ;
        RECT 2090.400 17.670 2090.540 1700.000 ;
        RECT 2090.340 17.350 2090.600 17.670 ;
        RECT 2286.300 17.350 2286.560 17.670 ;
        RECT 2286.360 2.400 2286.500 17.350 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2097.670 1688.680 2097.990 1688.740 ;
        RECT 2104.110 1688.680 2104.430 1688.740 ;
        RECT 2097.670 1688.540 2104.430 1688.680 ;
        RECT 2097.670 1688.480 2097.990 1688.540 ;
        RECT 2104.110 1688.480 2104.430 1688.540 ;
        RECT 2104.110 17.920 2104.430 17.980 ;
        RECT 2304.210 17.920 2304.530 17.980 ;
        RECT 2104.110 17.780 2304.530 17.920 ;
        RECT 2104.110 17.720 2104.430 17.780 ;
        RECT 2304.210 17.720 2304.530 17.780 ;
      LAYER via ;
        RECT 2097.700 1688.480 2097.960 1688.740 ;
        RECT 2104.140 1688.480 2104.400 1688.740 ;
        RECT 2104.140 17.720 2104.400 17.980 ;
        RECT 2304.240 17.720 2304.500 17.980 ;
      LAYER met2 ;
        RECT 2097.625 1700.000 2097.905 1704.000 ;
        RECT 2097.760 1688.770 2097.900 1700.000 ;
        RECT 2097.700 1688.450 2097.960 1688.770 ;
        RECT 2104.140 1688.450 2104.400 1688.770 ;
        RECT 2104.200 18.010 2104.340 1688.450 ;
        RECT 2104.140 17.690 2104.400 18.010 ;
        RECT 2304.240 17.690 2304.500 18.010 ;
        RECT 2304.300 2.400 2304.440 17.690 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2295.085 1686.485 2295.255 1689.035 ;
        RECT 2319.005 1352.605 2319.175 1376.575 ;
        RECT 2318.545 1256.045 2318.715 1304.155 ;
        RECT 2319.005 1173.085 2319.175 1207.255 ;
        RECT 2318.545 724.625 2318.715 738.735 ;
        RECT 2319.465 524.365 2319.635 572.475 ;
        RECT 2318.545 427.805 2318.715 470.815 ;
      LAYER mcon ;
        RECT 2295.085 1688.865 2295.255 1689.035 ;
        RECT 2319.005 1376.405 2319.175 1376.575 ;
        RECT 2318.545 1303.985 2318.715 1304.155 ;
        RECT 2319.005 1207.085 2319.175 1207.255 ;
        RECT 2318.545 738.565 2318.715 738.735 ;
        RECT 2319.465 572.305 2319.635 572.475 ;
        RECT 2318.545 470.645 2318.715 470.815 ;
      LAYER met1 ;
        RECT 2295.025 1689.020 2295.315 1689.065 ;
        RECT 2318.930 1689.020 2319.250 1689.080 ;
        RECT 2295.025 1688.880 2319.250 1689.020 ;
        RECT 2295.025 1688.835 2295.315 1688.880 ;
        RECT 2318.930 1688.820 2319.250 1688.880 ;
        RECT 2105.030 1686.640 2105.350 1686.700 ;
        RECT 2295.025 1686.640 2295.315 1686.685 ;
        RECT 2105.030 1686.500 2295.315 1686.640 ;
        RECT 2105.030 1686.440 2105.350 1686.500 ;
        RECT 2295.025 1686.455 2295.315 1686.500 ;
        RECT 2318.470 1531.940 2318.790 1532.000 ;
        RECT 2319.390 1531.940 2319.710 1532.000 ;
        RECT 2318.470 1531.800 2319.710 1531.940 ;
        RECT 2318.470 1531.740 2318.790 1531.800 ;
        RECT 2319.390 1531.740 2319.710 1531.800 ;
        RECT 2318.930 1376.560 2319.250 1376.620 ;
        RECT 2318.735 1376.420 2319.250 1376.560 ;
        RECT 2318.930 1376.360 2319.250 1376.420 ;
        RECT 2318.945 1352.760 2319.235 1352.805 ;
        RECT 2319.390 1352.760 2319.710 1352.820 ;
        RECT 2318.945 1352.620 2319.710 1352.760 ;
        RECT 2318.945 1352.575 2319.235 1352.620 ;
        RECT 2319.390 1352.560 2319.710 1352.620 ;
        RECT 2318.485 1304.140 2318.775 1304.185 ;
        RECT 2318.930 1304.140 2319.250 1304.200 ;
        RECT 2318.485 1304.000 2319.250 1304.140 ;
        RECT 2318.485 1303.955 2318.775 1304.000 ;
        RECT 2318.930 1303.940 2319.250 1304.000 ;
        RECT 2318.470 1256.200 2318.790 1256.260 ;
        RECT 2318.470 1256.060 2318.985 1256.200 ;
        RECT 2318.470 1256.000 2318.790 1256.060 ;
        RECT 2318.930 1207.240 2319.250 1207.300 ;
        RECT 2318.735 1207.100 2319.250 1207.240 ;
        RECT 2318.930 1207.040 2319.250 1207.100 ;
        RECT 2318.945 1173.240 2319.235 1173.285 ;
        RECT 2319.850 1173.240 2320.170 1173.300 ;
        RECT 2318.945 1173.100 2320.170 1173.240 ;
        RECT 2318.945 1173.055 2319.235 1173.100 ;
        RECT 2319.850 1173.040 2320.170 1173.100 ;
        RECT 2318.930 1111.020 2319.250 1111.080 ;
        RECT 2320.310 1111.020 2320.630 1111.080 ;
        RECT 2318.930 1110.880 2320.630 1111.020 ;
        RECT 2318.930 1110.820 2319.250 1110.880 ;
        RECT 2320.310 1110.820 2320.630 1110.880 ;
        RECT 2320.310 1077.020 2320.630 1077.080 ;
        RECT 2319.940 1076.880 2320.630 1077.020 ;
        RECT 2319.940 1076.400 2320.080 1076.880 ;
        RECT 2320.310 1076.820 2320.630 1076.880 ;
        RECT 2319.850 1076.140 2320.170 1076.400 ;
        RECT 2318.930 1014.460 2319.250 1014.520 ;
        RECT 2320.310 1014.460 2320.630 1014.520 ;
        RECT 2318.930 1014.320 2320.630 1014.460 ;
        RECT 2318.930 1014.260 2319.250 1014.320 ;
        RECT 2320.310 1014.260 2320.630 1014.320 ;
        RECT 2320.310 980.460 2320.630 980.520 ;
        RECT 2319.940 980.320 2320.630 980.460 ;
        RECT 2319.940 979.840 2320.080 980.320 ;
        RECT 2320.310 980.260 2320.630 980.320 ;
        RECT 2319.850 979.580 2320.170 979.840 ;
        RECT 2318.930 917.900 2319.250 917.960 ;
        RECT 2320.310 917.900 2320.630 917.960 ;
        RECT 2318.930 917.760 2320.630 917.900 ;
        RECT 2318.930 917.700 2319.250 917.760 ;
        RECT 2320.310 917.700 2320.630 917.760 ;
        RECT 2319.390 869.620 2319.710 869.680 ;
        RECT 2320.310 869.620 2320.630 869.680 ;
        RECT 2319.390 869.480 2320.630 869.620 ;
        RECT 2319.390 869.420 2319.710 869.480 ;
        RECT 2320.310 869.420 2320.630 869.480 ;
        RECT 2318.485 738.720 2318.775 738.765 ;
        RECT 2318.930 738.720 2319.250 738.780 ;
        RECT 2318.485 738.580 2319.250 738.720 ;
        RECT 2318.485 738.535 2318.775 738.580 ;
        RECT 2318.930 738.520 2319.250 738.580 ;
        RECT 2318.470 724.780 2318.790 724.840 ;
        RECT 2318.470 724.640 2318.985 724.780 ;
        RECT 2318.470 724.580 2318.790 724.640 ;
        RECT 2318.470 689.900 2318.790 690.160 ;
        RECT 2318.560 689.760 2318.700 689.900 ;
        RECT 2319.390 689.760 2319.710 689.820 ;
        RECT 2318.560 689.620 2319.710 689.760 ;
        RECT 2319.390 689.560 2319.710 689.620 ;
        RECT 2319.390 652.020 2319.710 652.080 ;
        RECT 2320.310 652.020 2320.630 652.080 ;
        RECT 2319.390 651.880 2320.630 652.020 ;
        RECT 2319.390 651.820 2319.710 651.880 ;
        RECT 2320.310 651.820 2320.630 651.880 ;
        RECT 2319.405 572.460 2319.695 572.505 ;
        RECT 2319.850 572.460 2320.170 572.520 ;
        RECT 2319.405 572.320 2320.170 572.460 ;
        RECT 2319.405 572.275 2319.695 572.320 ;
        RECT 2319.850 572.260 2320.170 572.320 ;
        RECT 2319.390 524.520 2319.710 524.580 ;
        RECT 2319.195 524.380 2319.710 524.520 ;
        RECT 2319.390 524.320 2319.710 524.380 ;
        RECT 2318.470 476.240 2318.790 476.300 ;
        RECT 2319.390 476.240 2319.710 476.300 ;
        RECT 2318.470 476.100 2319.710 476.240 ;
        RECT 2318.470 476.040 2318.790 476.100 ;
        RECT 2319.390 476.040 2319.710 476.100 ;
        RECT 2318.470 470.800 2318.790 470.860 ;
        RECT 2318.275 470.660 2318.790 470.800 ;
        RECT 2318.470 470.600 2318.790 470.660 ;
        RECT 2318.485 427.960 2318.775 428.005 ;
        RECT 2319.390 427.960 2319.710 428.020 ;
        RECT 2318.485 427.820 2319.710 427.960 ;
        RECT 2318.485 427.775 2318.775 427.820 ;
        RECT 2319.390 427.760 2319.710 427.820 ;
        RECT 2318.470 2.960 2318.790 3.020 ;
        RECT 2322.150 2.960 2322.470 3.020 ;
        RECT 2318.470 2.820 2322.470 2.960 ;
        RECT 2318.470 2.760 2318.790 2.820 ;
        RECT 2322.150 2.760 2322.470 2.820 ;
      LAYER via ;
        RECT 2318.960 1688.820 2319.220 1689.080 ;
        RECT 2105.060 1686.440 2105.320 1686.700 ;
        RECT 2318.500 1531.740 2318.760 1532.000 ;
        RECT 2319.420 1531.740 2319.680 1532.000 ;
        RECT 2318.960 1376.360 2319.220 1376.620 ;
        RECT 2319.420 1352.560 2319.680 1352.820 ;
        RECT 2318.960 1303.940 2319.220 1304.200 ;
        RECT 2318.500 1256.000 2318.760 1256.260 ;
        RECT 2318.960 1207.040 2319.220 1207.300 ;
        RECT 2319.880 1173.040 2320.140 1173.300 ;
        RECT 2318.960 1110.820 2319.220 1111.080 ;
        RECT 2320.340 1110.820 2320.600 1111.080 ;
        RECT 2320.340 1076.820 2320.600 1077.080 ;
        RECT 2319.880 1076.140 2320.140 1076.400 ;
        RECT 2318.960 1014.260 2319.220 1014.520 ;
        RECT 2320.340 1014.260 2320.600 1014.520 ;
        RECT 2320.340 980.260 2320.600 980.520 ;
        RECT 2319.880 979.580 2320.140 979.840 ;
        RECT 2318.960 917.700 2319.220 917.960 ;
        RECT 2320.340 917.700 2320.600 917.960 ;
        RECT 2319.420 869.420 2319.680 869.680 ;
        RECT 2320.340 869.420 2320.600 869.680 ;
        RECT 2318.960 738.520 2319.220 738.780 ;
        RECT 2318.500 724.580 2318.760 724.840 ;
        RECT 2318.500 689.900 2318.760 690.160 ;
        RECT 2319.420 689.560 2319.680 689.820 ;
        RECT 2319.420 651.820 2319.680 652.080 ;
        RECT 2320.340 651.820 2320.600 652.080 ;
        RECT 2319.880 572.260 2320.140 572.520 ;
        RECT 2319.420 524.320 2319.680 524.580 ;
        RECT 2318.500 476.040 2318.760 476.300 ;
        RECT 2319.420 476.040 2319.680 476.300 ;
        RECT 2318.500 470.600 2318.760 470.860 ;
        RECT 2319.420 427.760 2319.680 428.020 ;
        RECT 2318.500 2.760 2318.760 3.020 ;
        RECT 2322.180 2.760 2322.440 3.020 ;
      LAYER met2 ;
        RECT 2104.985 1700.000 2105.265 1704.000 ;
        RECT 2105.120 1686.730 2105.260 1700.000 ;
        RECT 2318.960 1688.790 2319.220 1689.110 ;
        RECT 2105.060 1686.410 2105.320 1686.730 ;
        RECT 2319.020 1607.930 2319.160 1688.790 ;
        RECT 2318.560 1607.790 2319.160 1607.930 ;
        RECT 2318.560 1580.050 2318.700 1607.790 ;
        RECT 2318.560 1579.910 2319.620 1580.050 ;
        RECT 2319.480 1532.030 2319.620 1579.910 ;
        RECT 2318.500 1531.710 2318.760 1532.030 ;
        RECT 2319.420 1531.710 2319.680 1532.030 ;
        RECT 2318.560 1510.690 2318.700 1531.710 ;
        RECT 2318.560 1510.550 2319.160 1510.690 ;
        RECT 2319.020 1463.090 2319.160 1510.550 ;
        RECT 2319.020 1462.950 2319.620 1463.090 ;
        RECT 2319.480 1462.410 2319.620 1462.950 ;
        RECT 2319.020 1462.270 2319.620 1462.410 ;
        RECT 2319.020 1414.810 2319.160 1462.270 ;
        RECT 2318.560 1414.670 2319.160 1414.810 ;
        RECT 2318.560 1414.130 2318.700 1414.670 ;
        RECT 2318.560 1413.990 2319.160 1414.130 ;
        RECT 2319.020 1376.650 2319.160 1413.990 ;
        RECT 2318.960 1376.330 2319.220 1376.650 ;
        RECT 2319.420 1352.530 2319.680 1352.850 ;
        RECT 2319.480 1317.570 2319.620 1352.530 ;
        RECT 2319.020 1317.430 2319.620 1317.570 ;
        RECT 2319.020 1304.230 2319.160 1317.430 ;
        RECT 2318.960 1303.910 2319.220 1304.230 ;
        RECT 2318.500 1255.970 2318.760 1256.290 ;
        RECT 2318.560 1221.010 2318.700 1255.970 ;
        RECT 2318.560 1220.870 2319.160 1221.010 ;
        RECT 2319.020 1207.330 2319.160 1220.870 ;
        RECT 2318.960 1207.010 2319.220 1207.330 ;
        RECT 2319.880 1173.010 2320.140 1173.330 ;
        RECT 2319.940 1159.245 2320.080 1173.010 ;
        RECT 2318.950 1158.875 2319.230 1159.245 ;
        RECT 2319.870 1158.875 2320.150 1159.245 ;
        RECT 2319.020 1111.110 2319.160 1158.875 ;
        RECT 2318.960 1110.790 2319.220 1111.110 ;
        RECT 2320.340 1110.790 2320.600 1111.110 ;
        RECT 2320.400 1077.110 2320.540 1110.790 ;
        RECT 2320.340 1076.790 2320.600 1077.110 ;
        RECT 2319.880 1076.110 2320.140 1076.430 ;
        RECT 2319.940 1062.685 2320.080 1076.110 ;
        RECT 2318.950 1062.315 2319.230 1062.685 ;
        RECT 2319.870 1062.315 2320.150 1062.685 ;
        RECT 2319.020 1014.550 2319.160 1062.315 ;
        RECT 2318.960 1014.230 2319.220 1014.550 ;
        RECT 2320.340 1014.230 2320.600 1014.550 ;
        RECT 2320.400 980.550 2320.540 1014.230 ;
        RECT 2320.340 980.230 2320.600 980.550 ;
        RECT 2319.880 979.550 2320.140 979.870 ;
        RECT 2319.940 966.125 2320.080 979.550 ;
        RECT 2318.950 965.755 2319.230 966.125 ;
        RECT 2319.870 965.755 2320.150 966.125 ;
        RECT 2319.020 917.990 2319.160 965.755 ;
        RECT 2318.960 917.670 2319.220 917.990 ;
        RECT 2320.340 917.670 2320.600 917.990 ;
        RECT 2320.400 869.710 2320.540 917.670 ;
        RECT 2319.420 869.390 2319.680 869.710 ;
        RECT 2320.340 869.390 2320.600 869.710 ;
        RECT 2319.480 787.170 2319.620 869.390 ;
        RECT 2318.560 787.030 2319.620 787.170 ;
        RECT 2318.560 786.490 2318.700 787.030 ;
        RECT 2318.560 786.350 2319.160 786.490 ;
        RECT 2319.020 738.810 2319.160 786.350 ;
        RECT 2318.960 738.490 2319.220 738.810 ;
        RECT 2318.500 724.550 2318.760 724.870 ;
        RECT 2318.560 690.190 2318.700 724.550 ;
        RECT 2318.500 689.870 2318.760 690.190 ;
        RECT 2319.420 689.530 2319.680 689.850 ;
        RECT 2319.480 652.110 2319.620 689.530 ;
        RECT 2319.420 651.790 2319.680 652.110 ;
        RECT 2320.340 651.790 2320.600 652.110 ;
        RECT 2320.400 628.165 2320.540 651.790 ;
        RECT 2319.410 627.795 2319.690 628.165 ;
        RECT 2320.330 627.795 2320.610 628.165 ;
        RECT 2319.480 572.970 2319.620 627.795 ;
        RECT 2319.480 572.830 2320.080 572.970 ;
        RECT 2319.940 572.550 2320.080 572.830 ;
        RECT 2319.880 572.230 2320.140 572.550 ;
        RECT 2319.420 524.290 2319.680 524.610 ;
        RECT 2319.480 476.330 2319.620 524.290 ;
        RECT 2318.500 476.010 2318.760 476.330 ;
        RECT 2319.420 476.010 2319.680 476.330 ;
        RECT 2318.560 470.890 2318.700 476.010 ;
        RECT 2318.500 470.570 2318.760 470.890 ;
        RECT 2319.420 427.730 2319.680 428.050 ;
        RECT 2319.480 352.650 2319.620 427.730 ;
        RECT 2319.020 352.510 2319.620 352.650 ;
        RECT 2319.020 351.970 2319.160 352.510 ;
        RECT 2318.560 351.830 2319.160 351.970 ;
        RECT 2318.560 3.050 2318.700 351.830 ;
        RECT 2318.500 2.730 2318.760 3.050 ;
        RECT 2322.180 2.730 2322.440 3.050 ;
        RECT 2322.240 2.400 2322.380 2.730 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
      LAYER via2 ;
        RECT 2318.950 1158.920 2319.230 1159.200 ;
        RECT 2319.870 1158.920 2320.150 1159.200 ;
        RECT 2318.950 1062.360 2319.230 1062.640 ;
        RECT 2319.870 1062.360 2320.150 1062.640 ;
        RECT 2318.950 965.800 2319.230 966.080 ;
        RECT 2319.870 965.800 2320.150 966.080 ;
        RECT 2319.410 627.840 2319.690 628.120 ;
        RECT 2320.330 627.840 2320.610 628.120 ;
      LAYER met3 ;
        RECT 2318.925 1159.210 2319.255 1159.225 ;
        RECT 2319.845 1159.210 2320.175 1159.225 ;
        RECT 2318.925 1158.910 2320.175 1159.210 ;
        RECT 2318.925 1158.895 2319.255 1158.910 ;
        RECT 2319.845 1158.895 2320.175 1158.910 ;
        RECT 2318.925 1062.650 2319.255 1062.665 ;
        RECT 2319.845 1062.650 2320.175 1062.665 ;
        RECT 2318.925 1062.350 2320.175 1062.650 ;
        RECT 2318.925 1062.335 2319.255 1062.350 ;
        RECT 2319.845 1062.335 2320.175 1062.350 ;
        RECT 2318.925 966.090 2319.255 966.105 ;
        RECT 2319.845 966.090 2320.175 966.105 ;
        RECT 2318.925 965.790 2320.175 966.090 ;
        RECT 2318.925 965.775 2319.255 965.790 ;
        RECT 2319.845 965.775 2320.175 965.790 ;
        RECT 2319.385 628.130 2319.715 628.145 ;
        RECT 2320.305 628.130 2320.635 628.145 ;
        RECT 2319.385 627.830 2320.635 628.130 ;
        RECT 2319.385 627.815 2319.715 627.830 ;
        RECT 2320.305 627.815 2320.635 627.830 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2126.265 17.085 2126.435 19.975 ;
      LAYER mcon ;
        RECT 2126.265 19.805 2126.435 19.975 ;
      LAYER met1 ;
        RECT 2112.390 1688.680 2112.710 1688.740 ;
        RECT 2122.050 1688.680 2122.370 1688.740 ;
        RECT 2112.390 1688.540 2122.370 1688.680 ;
        RECT 2112.390 1688.480 2112.710 1688.540 ;
        RECT 2122.050 1688.480 2122.370 1688.540 ;
        RECT 2122.050 19.960 2122.370 20.020 ;
        RECT 2126.205 19.960 2126.495 20.005 ;
        RECT 2122.050 19.820 2126.495 19.960 ;
        RECT 2122.050 19.760 2122.370 19.820 ;
        RECT 2126.205 19.775 2126.495 19.820 ;
        RECT 2126.205 17.240 2126.495 17.285 ;
        RECT 2339.630 17.240 2339.950 17.300 ;
        RECT 2126.205 17.100 2339.950 17.240 ;
        RECT 2126.205 17.055 2126.495 17.100 ;
        RECT 2339.630 17.040 2339.950 17.100 ;
      LAYER via ;
        RECT 2112.420 1688.480 2112.680 1688.740 ;
        RECT 2122.080 1688.480 2122.340 1688.740 ;
        RECT 2122.080 19.760 2122.340 20.020 ;
        RECT 2339.660 17.040 2339.920 17.300 ;
      LAYER met2 ;
        RECT 2112.345 1700.000 2112.625 1704.000 ;
        RECT 2112.480 1688.770 2112.620 1700.000 ;
        RECT 2112.420 1688.450 2112.680 1688.770 ;
        RECT 2122.080 1688.450 2122.340 1688.770 ;
        RECT 2122.140 20.050 2122.280 1688.450 ;
        RECT 2122.080 19.730 2122.340 20.050 ;
        RECT 2339.660 17.010 2339.920 17.330 ;
        RECT 2339.720 2.400 2339.860 17.010 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2139.145 1684.105 2139.315 1685.635 ;
        RECT 2163.525 1685.465 2163.695 1687.675 ;
        RECT 2185.605 1683.085 2185.775 1687.675 ;
        RECT 2221.485 1683.085 2221.655 1684.615 ;
        RECT 2295.545 1684.445 2295.715 1686.655 ;
      LAYER mcon ;
        RECT 2163.525 1687.505 2163.695 1687.675 ;
        RECT 2139.145 1685.465 2139.315 1685.635 ;
        RECT 2185.605 1687.505 2185.775 1687.675 ;
        RECT 2295.545 1686.485 2295.715 1686.655 ;
        RECT 2221.485 1684.445 2221.655 1684.615 ;
      LAYER met1 ;
        RECT 2163.465 1687.660 2163.755 1687.705 ;
        RECT 2185.545 1687.660 2185.835 1687.705 ;
        RECT 2163.465 1687.520 2185.835 1687.660 ;
        RECT 2163.465 1687.475 2163.755 1687.520 ;
        RECT 2185.545 1687.475 2185.835 1687.520 ;
        RECT 2295.485 1686.640 2295.775 1686.685 ;
        RECT 2352.970 1686.640 2353.290 1686.700 ;
        RECT 2295.485 1686.500 2353.290 1686.640 ;
        RECT 2295.485 1686.455 2295.775 1686.500 ;
        RECT 2352.970 1686.440 2353.290 1686.500 ;
        RECT 2139.085 1685.620 2139.375 1685.665 ;
        RECT 2163.465 1685.620 2163.755 1685.665 ;
        RECT 2139.085 1685.480 2163.755 1685.620 ;
        RECT 2139.085 1685.435 2139.375 1685.480 ;
        RECT 2163.465 1685.435 2163.755 1685.480 ;
        RECT 2221.425 1684.600 2221.715 1684.645 ;
        RECT 2221.870 1684.600 2222.190 1684.660 ;
        RECT 2295.485 1684.600 2295.775 1684.645 ;
        RECT 2221.425 1684.460 2222.190 1684.600 ;
        RECT 2221.425 1684.415 2221.715 1684.460 ;
        RECT 2221.870 1684.400 2222.190 1684.460 ;
        RECT 2235.300 1684.460 2295.775 1684.600 ;
        RECT 2119.750 1684.260 2120.070 1684.320 ;
        RECT 2139.085 1684.260 2139.375 1684.305 ;
        RECT 2119.750 1684.120 2139.375 1684.260 ;
        RECT 2119.750 1684.060 2120.070 1684.120 ;
        RECT 2139.085 1684.075 2139.375 1684.120 ;
        RECT 2221.870 1683.920 2222.190 1683.980 ;
        RECT 2235.300 1683.920 2235.440 1684.460 ;
        RECT 2295.485 1684.415 2295.775 1684.460 ;
        RECT 2221.870 1683.780 2235.440 1683.920 ;
        RECT 2221.870 1683.720 2222.190 1683.780 ;
        RECT 2185.545 1683.240 2185.835 1683.285 ;
        RECT 2221.425 1683.240 2221.715 1683.285 ;
        RECT 2185.545 1683.100 2221.715 1683.240 ;
        RECT 2185.545 1683.055 2185.835 1683.100 ;
        RECT 2221.425 1683.055 2221.715 1683.100 ;
      LAYER via ;
        RECT 2353.000 1686.440 2353.260 1686.700 ;
        RECT 2221.900 1684.400 2222.160 1684.660 ;
        RECT 2119.780 1684.060 2120.040 1684.320 ;
        RECT 2221.900 1683.720 2222.160 1683.980 ;
      LAYER met2 ;
        RECT 2119.705 1700.000 2119.985 1704.000 ;
        RECT 2119.840 1684.350 2119.980 1700.000 ;
        RECT 2353.000 1686.410 2353.260 1686.730 ;
        RECT 2221.900 1684.370 2222.160 1684.690 ;
        RECT 2119.780 1684.030 2120.040 1684.350 ;
        RECT 2221.960 1684.010 2222.100 1684.370 ;
        RECT 2221.900 1683.690 2222.160 1684.010 ;
        RECT 2353.060 16.730 2353.200 1686.410 ;
        RECT 2353.060 16.590 2357.800 16.730 ;
        RECT 2357.660 2.400 2357.800 16.590 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2162.605 14.365 2162.775 16.575 ;
        RECT 2179.625 14.365 2179.795 15.215 ;
      LAYER mcon ;
        RECT 2162.605 16.405 2162.775 16.575 ;
        RECT 2179.625 15.045 2179.795 15.215 ;
      LAYER met1 ;
        RECT 2127.110 1688.680 2127.430 1688.740 ;
        RECT 2142.290 1688.680 2142.610 1688.740 ;
        RECT 2127.110 1688.540 2142.610 1688.680 ;
        RECT 2127.110 1688.480 2127.430 1688.540 ;
        RECT 2142.290 1688.480 2142.610 1688.540 ;
        RECT 2142.290 16.560 2142.610 16.620 ;
        RECT 2162.545 16.560 2162.835 16.605 ;
        RECT 2142.290 16.420 2162.835 16.560 ;
        RECT 2142.290 16.360 2142.610 16.420 ;
        RECT 2162.545 16.375 2162.835 16.420 ;
        RECT 2179.565 15.200 2179.855 15.245 ;
        RECT 2375.510 15.200 2375.830 15.260 ;
        RECT 2179.565 15.060 2375.830 15.200 ;
        RECT 2179.565 15.015 2179.855 15.060 ;
        RECT 2375.510 15.000 2375.830 15.060 ;
        RECT 2162.545 14.520 2162.835 14.565 ;
        RECT 2179.565 14.520 2179.855 14.565 ;
        RECT 2162.545 14.380 2179.855 14.520 ;
        RECT 2162.545 14.335 2162.835 14.380 ;
        RECT 2179.565 14.335 2179.855 14.380 ;
      LAYER via ;
        RECT 2127.140 1688.480 2127.400 1688.740 ;
        RECT 2142.320 1688.480 2142.580 1688.740 ;
        RECT 2142.320 16.360 2142.580 16.620 ;
        RECT 2375.540 15.000 2375.800 15.260 ;
      LAYER met2 ;
        RECT 2127.065 1700.000 2127.345 1704.000 ;
        RECT 2127.200 1688.770 2127.340 1700.000 ;
        RECT 2127.140 1688.450 2127.400 1688.770 ;
        RECT 2142.320 1688.450 2142.580 1688.770 ;
        RECT 2142.380 16.650 2142.520 1688.450 ;
        RECT 2142.320 16.330 2142.580 16.650 ;
        RECT 2375.540 14.970 2375.800 15.290 ;
        RECT 2375.600 2.400 2375.740 14.970 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2163.065 1685.125 2163.235 1687.675 ;
      LAYER mcon ;
        RECT 2163.065 1687.505 2163.235 1687.675 ;
      LAYER met1 ;
        RECT 2135.850 1687.660 2136.170 1687.720 ;
        RECT 2163.005 1687.660 2163.295 1687.705 ;
        RECT 2135.850 1687.520 2163.295 1687.660 ;
        RECT 2135.850 1687.460 2136.170 1687.520 ;
        RECT 2163.005 1687.475 2163.295 1687.520 ;
        RECT 2163.005 1685.280 2163.295 1685.325 ;
        RECT 2221.870 1685.280 2222.190 1685.340 ;
        RECT 2163.005 1685.140 2222.190 1685.280 ;
        RECT 2163.005 1685.095 2163.295 1685.140 ;
        RECT 2221.870 1685.080 2222.190 1685.140 ;
        RECT 2223.710 1685.280 2224.030 1685.340 ;
        RECT 2387.930 1685.280 2388.250 1685.340 ;
        RECT 2223.710 1685.140 2388.250 1685.280 ;
        RECT 2223.710 1685.080 2224.030 1685.140 ;
        RECT 2387.930 1685.080 2388.250 1685.140 ;
      LAYER via ;
        RECT 2135.880 1687.460 2136.140 1687.720 ;
        RECT 2221.900 1685.080 2222.160 1685.340 ;
        RECT 2223.740 1685.080 2224.000 1685.340 ;
        RECT 2387.960 1685.080 2388.220 1685.340 ;
      LAYER met2 ;
        RECT 2134.425 1700.410 2134.705 1704.000 ;
        RECT 2134.425 1700.270 2136.080 1700.410 ;
        RECT 2134.425 1700.000 2134.705 1700.270 ;
        RECT 2135.940 1687.750 2136.080 1700.270 ;
        RECT 2135.880 1687.430 2136.140 1687.750 ;
        RECT 2221.960 1685.370 2223.940 1685.450 ;
        RECT 2221.900 1685.310 2224.000 1685.370 ;
        RECT 2221.900 1685.050 2222.160 1685.310 ;
        RECT 2223.740 1685.050 2224.000 1685.310 ;
        RECT 2387.960 1685.050 2388.220 1685.370 ;
        RECT 2388.020 16.730 2388.160 1685.050 ;
        RECT 2388.020 16.590 2393.680 16.730 ;
        RECT 2393.540 2.400 2393.680 16.590 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 2141.830 1684.260 2142.150 1684.320 ;
        RECT 2156.090 1684.260 2156.410 1684.320 ;
        RECT 2141.830 1684.120 2156.410 1684.260 ;
        RECT 2141.830 1684.060 2142.150 1684.120 ;
        RECT 2156.090 1684.060 2156.410 1684.120 ;
        RECT 2156.090 15.540 2156.410 15.600 ;
        RECT 2156.090 15.400 2388.160 15.540 ;
        RECT 2156.090 15.340 2156.410 15.400 ;
        RECT 2388.020 15.200 2388.160 15.400 ;
        RECT 2411.390 15.200 2411.710 15.260 ;
        RECT 2388.020 15.060 2411.710 15.200 ;
        RECT 2411.390 15.000 2411.710 15.060 ;
      LAYER via ;
        RECT 2141.860 1684.060 2142.120 1684.320 ;
        RECT 2156.120 1684.060 2156.380 1684.320 ;
        RECT 2156.120 15.340 2156.380 15.600 ;
        RECT 2411.420 15.000 2411.680 15.260 ;
      LAYER met2 ;
        RECT 2141.785 1700.000 2142.065 1704.000 ;
        RECT 2141.920 1684.350 2142.060 1700.000 ;
        RECT 2141.860 1684.030 2142.120 1684.350 ;
        RECT 2156.120 1684.030 2156.380 1684.350 ;
        RECT 2156.180 15.630 2156.320 1684.030 ;
        RECT 2156.120 15.310 2156.380 15.630 ;
        RECT 2411.420 14.970 2411.680 15.290 ;
        RECT 2411.480 2.400 2411.620 14.970 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 806.910 48.520 807.230 48.580 ;
        RECT 1477.130 48.520 1477.450 48.580 ;
        RECT 806.910 48.380 1477.450 48.520 ;
        RECT 806.910 48.320 807.230 48.380 ;
        RECT 1477.130 48.320 1477.450 48.380 ;
      LAYER via ;
        RECT 806.940 48.320 807.200 48.580 ;
        RECT 1477.160 48.320 1477.420 48.580 ;
      LAYER met2 ;
        RECT 1480.305 1700.410 1480.585 1704.000 ;
        RECT 1478.600 1700.270 1480.585 1700.410 ;
        RECT 1478.600 1678.480 1478.740 1700.270 ;
        RECT 1480.305 1700.000 1480.585 1700.270 ;
        RECT 1477.220 1678.340 1478.740 1678.480 ;
        RECT 1477.220 48.610 1477.360 1678.340 ;
        RECT 806.940 48.290 807.200 48.610 ;
        RECT 1477.160 48.290 1477.420 48.610 ;
        RECT 807.000 17.410 807.140 48.290 ;
        RECT 805.620 17.270 807.140 17.410 ;
        RECT 805.620 2.400 805.760 17.270 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1145.470 24.720 1145.790 24.780 ;
        RECT 1121.640 24.580 1145.790 24.720 ;
        RECT 2.830 24.380 3.150 24.440 ;
        RECT 1121.640 24.380 1121.780 24.580 ;
        RECT 1145.470 24.520 1145.790 24.580 ;
        RECT 2.830 24.240 1121.780 24.380 ;
        RECT 2.830 24.180 3.150 24.240 ;
      LAYER via ;
        RECT 2.860 24.180 3.120 24.440 ;
        RECT 1145.500 24.520 1145.760 24.780 ;
      LAYER met2 ;
        RECT 1150.025 1700.410 1150.305 1704.000 ;
        RECT 1145.560 1700.270 1150.305 1700.410 ;
        RECT 1145.560 24.810 1145.700 1700.270 ;
        RECT 1150.025 1700.000 1150.305 1700.270 ;
        RECT 1145.500 24.490 1145.760 24.810 ;
        RECT 2.860 24.150 3.120 24.470 ;
        RECT 2.920 2.400 3.060 24.150 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1120.705 21.165 1120.875 24.055 ;
      LAYER mcon ;
        RECT 1120.705 23.885 1120.875 24.055 ;
      LAYER met1 ;
        RECT 8.350 24.040 8.670 24.100 ;
        RECT 1120.645 24.040 1120.935 24.085 ;
        RECT 8.350 23.900 1120.935 24.040 ;
        RECT 8.350 23.840 8.670 23.900 ;
        RECT 1120.645 23.855 1120.935 23.900 ;
        RECT 1120.645 21.320 1120.935 21.365 ;
        RECT 1152.370 21.320 1152.690 21.380 ;
        RECT 1120.645 21.180 1152.690 21.320 ;
        RECT 1120.645 21.135 1120.935 21.180 ;
        RECT 1152.370 21.120 1152.690 21.180 ;
      LAYER via ;
        RECT 8.380 23.840 8.640 24.100 ;
        RECT 1152.400 21.120 1152.660 21.380 ;
      LAYER met2 ;
        RECT 1152.325 1700.000 1152.605 1704.000 ;
        RECT 8.380 23.810 8.640 24.130 ;
        RECT 8.440 2.400 8.580 23.810 ;
        RECT 1152.460 21.410 1152.600 1700.000 ;
        RECT 1152.400 21.090 1152.660 21.410 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1121.165 23.885 1121.335 24.735 ;
      LAYER mcon ;
        RECT 1121.165 24.565 1121.335 24.735 ;
      LAYER met1 ;
        RECT 14.330 24.720 14.650 24.780 ;
        RECT 1121.105 24.720 1121.395 24.765 ;
        RECT 14.330 24.580 1121.395 24.720 ;
        RECT 14.330 24.520 14.650 24.580 ;
        RECT 1121.105 24.535 1121.395 24.580 ;
        RECT 1121.105 24.040 1121.395 24.085 ;
        RECT 1152.830 24.040 1153.150 24.100 ;
        RECT 1121.105 23.900 1153.150 24.040 ;
        RECT 1121.105 23.855 1121.395 23.900 ;
        RECT 1152.830 23.840 1153.150 23.900 ;
      LAYER via ;
        RECT 14.360 24.520 14.620 24.780 ;
        RECT 1152.860 23.840 1153.120 24.100 ;
      LAYER met2 ;
        RECT 1154.625 1700.410 1154.905 1704.000 ;
        RECT 1152.920 1700.270 1154.905 1700.410 ;
        RECT 14.360 24.490 14.620 24.810 ;
        RECT 14.420 2.400 14.560 24.490 ;
        RECT 1152.920 24.130 1153.060 1700.270 ;
        RECT 1154.625 1700.000 1154.905 1700.270 ;
        RECT 1152.860 23.810 1153.120 24.130 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1161.645 724.965 1161.815 772.735 ;
        RECT 1161.645 669.545 1161.815 717.655 ;
        RECT 1161.645 572.645 1161.815 620.755 ;
        RECT 1161.645 476.085 1161.815 524.195 ;
        RECT 1161.645 379.525 1161.815 427.635 ;
        RECT 1161.645 282.965 1161.815 330.395 ;
        RECT 1161.185 138.125 1161.355 185.895 ;
        RECT 1160.725 70.465 1160.895 113.815 ;
      LAYER mcon ;
        RECT 1161.645 772.565 1161.815 772.735 ;
        RECT 1161.645 717.485 1161.815 717.655 ;
        RECT 1161.645 620.585 1161.815 620.755 ;
        RECT 1161.645 524.025 1161.815 524.195 ;
        RECT 1161.645 427.465 1161.815 427.635 ;
        RECT 1161.645 330.225 1161.815 330.395 ;
        RECT 1161.185 185.725 1161.355 185.895 ;
        RECT 1160.725 113.645 1160.895 113.815 ;
      LAYER met1 ;
        RECT 1161.110 1607.760 1161.430 1607.820 ;
        RECT 1162.030 1607.760 1162.350 1607.820 ;
        RECT 1161.110 1607.620 1162.350 1607.760 ;
        RECT 1161.110 1607.560 1161.430 1607.620 ;
        RECT 1162.030 1607.560 1162.350 1607.620 ;
        RECT 1162.030 1559.820 1162.350 1559.880 ;
        RECT 1161.660 1559.680 1162.350 1559.820 ;
        RECT 1161.660 1559.200 1161.800 1559.680 ;
        RECT 1162.030 1559.620 1162.350 1559.680 ;
        RECT 1161.570 1558.940 1161.890 1559.200 ;
        RECT 1161.110 979.920 1161.430 980.180 ;
        RECT 1161.200 979.780 1161.340 979.920 ;
        RECT 1161.570 979.780 1161.890 979.840 ;
        RECT 1161.200 979.640 1161.890 979.780 ;
        RECT 1161.570 979.580 1161.890 979.640 ;
        RECT 1161.110 883.360 1161.430 883.620 ;
        RECT 1161.200 883.220 1161.340 883.360 ;
        RECT 1161.570 883.220 1161.890 883.280 ;
        RECT 1161.200 883.080 1161.890 883.220 ;
        RECT 1161.570 883.020 1161.890 883.080 ;
        RECT 1161.585 772.720 1161.875 772.765 ;
        RECT 1162.030 772.720 1162.350 772.780 ;
        RECT 1161.585 772.580 1162.350 772.720 ;
        RECT 1161.585 772.535 1161.875 772.580 ;
        RECT 1162.030 772.520 1162.350 772.580 ;
        RECT 1161.570 725.120 1161.890 725.180 ;
        RECT 1161.375 724.980 1161.890 725.120 ;
        RECT 1161.570 724.920 1161.890 724.980 ;
        RECT 1161.570 717.640 1161.890 717.700 ;
        RECT 1161.375 717.500 1161.890 717.640 ;
        RECT 1161.570 717.440 1161.890 717.500 ;
        RECT 1161.570 669.700 1161.890 669.760 ;
        RECT 1161.375 669.560 1161.890 669.700 ;
        RECT 1161.570 669.500 1161.890 669.560 ;
        RECT 1161.570 620.740 1161.890 620.800 ;
        RECT 1161.375 620.600 1161.890 620.740 ;
        RECT 1161.570 620.540 1161.890 620.600 ;
        RECT 1161.570 572.800 1161.890 572.860 ;
        RECT 1161.375 572.660 1161.890 572.800 ;
        RECT 1161.570 572.600 1161.890 572.660 ;
        RECT 1161.570 524.180 1161.890 524.240 ;
        RECT 1161.375 524.040 1161.890 524.180 ;
        RECT 1161.570 523.980 1161.890 524.040 ;
        RECT 1161.570 476.240 1161.890 476.300 ;
        RECT 1161.375 476.100 1161.890 476.240 ;
        RECT 1161.570 476.040 1161.890 476.100 ;
        RECT 1161.570 427.620 1161.890 427.680 ;
        RECT 1161.375 427.480 1161.890 427.620 ;
        RECT 1161.570 427.420 1161.890 427.480 ;
        RECT 1161.570 379.680 1161.890 379.740 ;
        RECT 1161.375 379.540 1161.890 379.680 ;
        RECT 1161.570 379.480 1161.890 379.540 ;
        RECT 1161.570 330.860 1161.890 331.120 ;
        RECT 1161.660 330.425 1161.800 330.860 ;
        RECT 1161.585 330.195 1161.875 330.425 ;
        RECT 1161.570 283.120 1161.890 283.180 ;
        RECT 1161.375 282.980 1161.890 283.120 ;
        RECT 1161.570 282.920 1161.890 282.980 ;
        RECT 1161.570 255.580 1161.890 255.640 ;
        RECT 1161.200 255.440 1161.890 255.580 ;
        RECT 1161.200 255.300 1161.340 255.440 ;
        RECT 1161.570 255.380 1161.890 255.440 ;
        RECT 1161.110 255.040 1161.430 255.300 ;
        RECT 1161.570 186.900 1161.890 186.960 ;
        RECT 1161.200 186.760 1161.890 186.900 ;
        RECT 1161.200 186.620 1161.340 186.760 ;
        RECT 1161.570 186.700 1161.890 186.760 ;
        RECT 1161.110 186.360 1161.430 186.620 ;
        RECT 1161.110 185.880 1161.430 185.940 ;
        RECT 1160.915 185.740 1161.430 185.880 ;
        RECT 1161.110 185.680 1161.430 185.740 ;
        RECT 1161.125 138.280 1161.415 138.325 ;
        RECT 1161.570 138.280 1161.890 138.340 ;
        RECT 1161.125 138.140 1161.890 138.280 ;
        RECT 1161.125 138.095 1161.415 138.140 ;
        RECT 1161.570 138.080 1161.890 138.140 ;
        RECT 1160.665 113.800 1160.955 113.845 ;
        RECT 1162.030 113.800 1162.350 113.860 ;
        RECT 1160.665 113.660 1162.350 113.800 ;
        RECT 1160.665 113.615 1160.955 113.660 ;
        RECT 1162.030 113.600 1162.350 113.660 ;
        RECT 1160.650 70.620 1160.970 70.680 ;
        RECT 1160.455 70.480 1160.970 70.620 ;
        RECT 1160.650 70.420 1160.970 70.480 ;
        RECT 38.250 25.060 38.570 25.120 ;
        RECT 1160.650 25.060 1160.970 25.120 ;
        RECT 38.250 24.920 1160.970 25.060 ;
        RECT 38.250 24.860 38.570 24.920 ;
        RECT 1160.650 24.860 1160.970 24.920 ;
      LAYER via ;
        RECT 1161.140 1607.560 1161.400 1607.820 ;
        RECT 1162.060 1607.560 1162.320 1607.820 ;
        RECT 1162.060 1559.620 1162.320 1559.880 ;
        RECT 1161.600 1558.940 1161.860 1559.200 ;
        RECT 1161.140 979.920 1161.400 980.180 ;
        RECT 1161.600 979.580 1161.860 979.840 ;
        RECT 1161.140 883.360 1161.400 883.620 ;
        RECT 1161.600 883.020 1161.860 883.280 ;
        RECT 1162.060 772.520 1162.320 772.780 ;
        RECT 1161.600 724.920 1161.860 725.180 ;
        RECT 1161.600 717.440 1161.860 717.700 ;
        RECT 1161.600 669.500 1161.860 669.760 ;
        RECT 1161.600 620.540 1161.860 620.800 ;
        RECT 1161.600 572.600 1161.860 572.860 ;
        RECT 1161.600 523.980 1161.860 524.240 ;
        RECT 1161.600 476.040 1161.860 476.300 ;
        RECT 1161.600 427.420 1161.860 427.680 ;
        RECT 1161.600 379.480 1161.860 379.740 ;
        RECT 1161.600 330.860 1161.860 331.120 ;
        RECT 1161.600 282.920 1161.860 283.180 ;
        RECT 1161.600 255.380 1161.860 255.640 ;
        RECT 1161.140 255.040 1161.400 255.300 ;
        RECT 1161.600 186.700 1161.860 186.960 ;
        RECT 1161.140 186.360 1161.400 186.620 ;
        RECT 1161.140 185.680 1161.400 185.940 ;
        RECT 1161.600 138.080 1161.860 138.340 ;
        RECT 1162.060 113.600 1162.320 113.860 ;
        RECT 1160.680 70.420 1160.940 70.680 ;
        RECT 38.280 24.860 38.540 25.120 ;
        RECT 1160.680 24.860 1160.940 25.120 ;
      LAYER met2 ;
        RECT 1164.285 1701.090 1164.565 1704.000 ;
        RECT 1162.580 1700.950 1164.565 1701.090 ;
        RECT 1162.580 1688.850 1162.720 1700.950 ;
        RECT 1164.285 1700.000 1164.565 1700.950 ;
        RECT 1161.200 1688.710 1162.720 1688.850 ;
        RECT 1161.200 1607.850 1161.340 1688.710 ;
        RECT 1161.140 1607.530 1161.400 1607.850 ;
        RECT 1162.060 1607.530 1162.320 1607.850 ;
        RECT 1162.120 1559.910 1162.260 1607.530 ;
        RECT 1162.060 1559.590 1162.320 1559.910 ;
        RECT 1161.600 1558.910 1161.860 1559.230 ;
        RECT 1161.660 1027.890 1161.800 1558.910 ;
        RECT 1161.200 1027.750 1161.800 1027.890 ;
        RECT 1161.200 980.210 1161.340 1027.750 ;
        RECT 1161.140 979.890 1161.400 980.210 ;
        RECT 1161.600 979.550 1161.860 979.870 ;
        RECT 1161.660 931.330 1161.800 979.550 ;
        RECT 1161.200 931.190 1161.800 931.330 ;
        RECT 1161.200 883.650 1161.340 931.190 ;
        RECT 1161.140 883.330 1161.400 883.650 ;
        RECT 1161.600 882.990 1161.860 883.310 ;
        RECT 1161.660 834.770 1161.800 882.990 ;
        RECT 1161.200 834.630 1161.800 834.770 ;
        RECT 1161.200 796.690 1161.340 834.630 ;
        RECT 1161.200 796.550 1162.260 796.690 ;
        RECT 1162.120 772.810 1162.260 796.550 ;
        RECT 1162.060 772.490 1162.320 772.810 ;
        RECT 1161.600 724.890 1161.860 725.210 ;
        RECT 1161.660 717.730 1161.800 724.890 ;
        RECT 1161.600 717.410 1161.860 717.730 ;
        RECT 1161.600 669.470 1161.860 669.790 ;
        RECT 1161.660 620.830 1161.800 669.470 ;
        RECT 1161.600 620.510 1161.860 620.830 ;
        RECT 1161.600 572.570 1161.860 572.890 ;
        RECT 1161.660 524.270 1161.800 572.570 ;
        RECT 1161.600 523.950 1161.860 524.270 ;
        RECT 1161.600 476.010 1161.860 476.330 ;
        RECT 1161.660 427.710 1161.800 476.010 ;
        RECT 1161.600 427.390 1161.860 427.710 ;
        RECT 1161.600 379.450 1161.860 379.770 ;
        RECT 1161.660 331.150 1161.800 379.450 ;
        RECT 1161.600 330.830 1161.860 331.150 ;
        RECT 1161.600 282.890 1161.860 283.210 ;
        RECT 1161.660 255.670 1161.800 282.890 ;
        RECT 1161.600 255.350 1161.860 255.670 ;
        RECT 1161.140 255.010 1161.400 255.330 ;
        RECT 1161.200 241.130 1161.340 255.010 ;
        RECT 1161.200 240.990 1161.800 241.130 ;
        RECT 1161.660 186.990 1161.800 240.990 ;
        RECT 1161.600 186.670 1161.860 186.990 ;
        RECT 1161.140 186.330 1161.400 186.650 ;
        RECT 1161.200 185.970 1161.340 186.330 ;
        RECT 1161.140 185.650 1161.400 185.970 ;
        RECT 1161.600 138.050 1161.860 138.370 ;
        RECT 1161.660 137.770 1161.800 138.050 ;
        RECT 1161.660 137.630 1162.260 137.770 ;
        RECT 1162.120 113.890 1162.260 137.630 ;
        RECT 1162.060 113.570 1162.320 113.890 ;
        RECT 1160.680 70.390 1160.940 70.710 ;
        RECT 1160.740 25.150 1160.880 70.390 ;
        RECT 38.280 24.830 38.540 25.150 ;
        RECT 1160.680 24.830 1160.940 25.150 ;
        RECT 38.340 2.400 38.480 24.830 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1242.530 1677.460 1242.850 1677.520 ;
        RECT 1245.750 1677.460 1246.070 1677.520 ;
        RECT 1242.530 1677.320 1246.070 1677.460 ;
        RECT 1242.530 1677.260 1242.850 1677.320 ;
        RECT 1245.750 1677.260 1246.070 1677.320 ;
        RECT 240.650 26.080 240.970 26.140 ;
        RECT 1242.530 26.080 1242.850 26.140 ;
        RECT 240.650 25.940 1242.850 26.080 ;
        RECT 240.650 25.880 240.970 25.940 ;
        RECT 1242.530 25.880 1242.850 25.940 ;
      LAYER via ;
        RECT 1242.560 1677.260 1242.820 1677.520 ;
        RECT 1245.780 1677.260 1246.040 1677.520 ;
        RECT 240.680 25.880 240.940 26.140 ;
        RECT 1242.560 25.880 1242.820 26.140 ;
      LAYER met2 ;
        RECT 1247.545 1700.410 1247.825 1704.000 ;
        RECT 1245.840 1700.270 1247.825 1700.410 ;
        RECT 1245.840 1677.550 1245.980 1700.270 ;
        RECT 1247.545 1700.000 1247.825 1700.270 ;
        RECT 1242.560 1677.230 1242.820 1677.550 ;
        RECT 1245.780 1677.230 1246.040 1677.550 ;
        RECT 1242.620 26.170 1242.760 1677.230 ;
        RECT 240.680 25.850 240.940 26.170 ;
        RECT 1242.560 25.850 1242.820 26.170 ;
        RECT 240.740 2.400 240.880 25.850 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1250.885 1635.485 1251.055 1677.815 ;
        RECT 1250.885 1562.725 1251.055 1587.035 ;
        RECT 1250.885 1297.185 1251.055 1321.495 ;
        RECT 1250.885 1207.425 1251.055 1255.875 ;
        RECT 1250.885 1152.345 1251.055 1173.255 ;
        RECT 1250.885 689.605 1251.055 717.655 ;
        RECT 1250.885 269.025 1251.055 283.135 ;
        RECT 1250.425 131.325 1250.595 179.095 ;
        RECT 1249.965 83.045 1250.135 110.755 ;
      LAYER mcon ;
        RECT 1250.885 1677.645 1251.055 1677.815 ;
        RECT 1250.885 1586.865 1251.055 1587.035 ;
        RECT 1250.885 1321.325 1251.055 1321.495 ;
        RECT 1250.885 1255.705 1251.055 1255.875 ;
        RECT 1250.885 1173.085 1251.055 1173.255 ;
        RECT 1250.885 717.485 1251.055 717.655 ;
        RECT 1250.885 282.965 1251.055 283.135 ;
        RECT 1250.425 178.925 1250.595 179.095 ;
        RECT 1249.965 110.585 1250.135 110.755 ;
      LAYER met1 ;
        RECT 1250.825 1677.800 1251.115 1677.845 ;
        RECT 1253.110 1677.800 1253.430 1677.860 ;
        RECT 1250.825 1677.660 1253.430 1677.800 ;
        RECT 1250.825 1677.615 1251.115 1677.660 ;
        RECT 1253.110 1677.600 1253.430 1677.660 ;
        RECT 1250.810 1635.640 1251.130 1635.700 ;
        RECT 1250.615 1635.500 1251.130 1635.640 ;
        RECT 1250.810 1635.440 1251.130 1635.500 ;
        RECT 1250.810 1587.020 1251.130 1587.080 ;
        RECT 1250.615 1586.880 1251.130 1587.020 ;
        RECT 1250.810 1586.820 1251.130 1586.880 ;
        RECT 1250.810 1562.880 1251.130 1562.940 ;
        RECT 1250.615 1562.740 1251.130 1562.880 ;
        RECT 1250.810 1562.680 1251.130 1562.740 ;
        RECT 1250.350 1400.700 1250.670 1400.760 ;
        RECT 1250.810 1400.700 1251.130 1400.760 ;
        RECT 1250.350 1400.560 1251.130 1400.700 ;
        RECT 1250.350 1400.500 1250.670 1400.560 ;
        RECT 1250.810 1400.500 1251.130 1400.560 ;
        RECT 1250.350 1369.760 1250.670 1369.820 ;
        RECT 1251.270 1369.760 1251.590 1369.820 ;
        RECT 1250.350 1369.620 1251.590 1369.760 ;
        RECT 1250.350 1369.560 1250.670 1369.620 ;
        RECT 1251.270 1369.560 1251.590 1369.620 ;
        RECT 1250.810 1321.480 1251.130 1321.540 ;
        RECT 1250.615 1321.340 1251.130 1321.480 ;
        RECT 1250.810 1321.280 1251.130 1321.340 ;
        RECT 1250.810 1297.340 1251.130 1297.400 ;
        RECT 1250.615 1297.200 1251.130 1297.340 ;
        RECT 1250.810 1297.140 1251.130 1297.200 ;
        RECT 1250.810 1255.860 1251.130 1255.920 ;
        RECT 1250.615 1255.720 1251.130 1255.860 ;
        RECT 1250.810 1255.660 1251.130 1255.720 ;
        RECT 1250.810 1207.580 1251.130 1207.640 ;
        RECT 1250.615 1207.440 1251.130 1207.580 ;
        RECT 1250.810 1207.380 1251.130 1207.440 ;
        RECT 1250.350 1173.240 1250.670 1173.300 ;
        RECT 1250.825 1173.240 1251.115 1173.285 ;
        RECT 1250.350 1173.100 1251.115 1173.240 ;
        RECT 1250.350 1173.040 1250.670 1173.100 ;
        RECT 1250.825 1173.055 1251.115 1173.100 ;
        RECT 1250.810 1152.500 1251.130 1152.560 ;
        RECT 1250.615 1152.360 1251.130 1152.500 ;
        RECT 1250.810 1152.300 1251.130 1152.360 ;
        RECT 1250.350 1062.740 1250.670 1062.800 ;
        RECT 1251.270 1062.740 1251.590 1062.800 ;
        RECT 1250.350 1062.600 1251.590 1062.740 ;
        RECT 1250.350 1062.540 1250.670 1062.600 ;
        RECT 1251.270 1062.540 1251.590 1062.600 ;
        RECT 1249.890 1055.600 1250.210 1055.660 ;
        RECT 1250.350 1055.600 1250.670 1055.660 ;
        RECT 1249.890 1055.460 1250.670 1055.600 ;
        RECT 1249.890 1055.400 1250.210 1055.460 ;
        RECT 1250.350 1055.400 1250.670 1055.460 ;
        RECT 1250.350 1007.320 1250.670 1007.380 ;
        RECT 1250.810 1007.320 1251.130 1007.380 ;
        RECT 1250.350 1007.180 1251.130 1007.320 ;
        RECT 1250.350 1007.120 1250.670 1007.180 ;
        RECT 1250.810 1007.120 1251.130 1007.180 ;
        RECT 1250.350 1000.520 1250.670 1000.580 ;
        RECT 1251.270 1000.520 1251.590 1000.580 ;
        RECT 1250.350 1000.380 1251.590 1000.520 ;
        RECT 1250.350 1000.320 1250.670 1000.380 ;
        RECT 1251.270 1000.320 1251.590 1000.380 ;
        RECT 1251.270 883.900 1251.590 883.960 ;
        RECT 1250.440 883.760 1251.590 883.900 ;
        RECT 1250.440 883.620 1250.580 883.760 ;
        RECT 1251.270 883.700 1251.590 883.760 ;
        RECT 1250.350 883.360 1250.670 883.620 ;
        RECT 1250.810 814.200 1251.130 814.260 ;
        RECT 1251.270 814.200 1251.590 814.260 ;
        RECT 1250.810 814.060 1251.590 814.200 ;
        RECT 1250.810 814.000 1251.130 814.060 ;
        RECT 1251.270 814.000 1251.590 814.060 ;
        RECT 1250.810 717.640 1251.130 717.700 ;
        RECT 1250.615 717.500 1251.130 717.640 ;
        RECT 1250.810 717.440 1251.130 717.500 ;
        RECT 1250.810 689.760 1251.130 689.820 ;
        RECT 1250.615 689.620 1251.130 689.760 ;
        RECT 1250.810 689.560 1251.130 689.620 ;
        RECT 1250.810 283.120 1251.130 283.180 ;
        RECT 1250.615 282.980 1251.130 283.120 ;
        RECT 1250.810 282.920 1251.130 282.980 ;
        RECT 1250.810 269.180 1251.130 269.240 ;
        RECT 1250.615 269.040 1251.130 269.180 ;
        RECT 1250.810 268.980 1251.130 269.040 ;
        RECT 1250.810 235.180 1251.130 235.240 ;
        RECT 1250.440 235.040 1251.130 235.180 ;
        RECT 1250.440 234.560 1250.580 235.040 ;
        RECT 1250.810 234.980 1251.130 235.040 ;
        RECT 1250.350 234.300 1250.670 234.560 ;
        RECT 1249.890 179.760 1250.210 179.820 ;
        RECT 1250.350 179.760 1250.670 179.820 ;
        RECT 1249.890 179.620 1250.670 179.760 ;
        RECT 1249.890 179.560 1250.210 179.620 ;
        RECT 1250.350 179.560 1250.670 179.620 ;
        RECT 1250.350 179.080 1250.670 179.140 ;
        RECT 1250.155 178.940 1250.670 179.080 ;
        RECT 1250.350 178.880 1250.670 178.940 ;
        RECT 1250.365 131.480 1250.655 131.525 ;
        RECT 1250.810 131.480 1251.130 131.540 ;
        RECT 1250.365 131.340 1251.130 131.480 ;
        RECT 1250.365 131.295 1250.655 131.340 ;
        RECT 1250.810 131.280 1251.130 131.340 ;
        RECT 1249.905 110.740 1250.195 110.785 ;
        RECT 1250.810 110.740 1251.130 110.800 ;
        RECT 1249.905 110.600 1251.130 110.740 ;
        RECT 1249.905 110.555 1250.195 110.600 ;
        RECT 1250.810 110.540 1251.130 110.600 ;
        RECT 1249.890 83.200 1250.210 83.260 ;
        RECT 1249.695 83.060 1250.210 83.200 ;
        RECT 1249.890 83.000 1250.210 83.060 ;
      LAYER via ;
        RECT 1253.140 1677.600 1253.400 1677.860 ;
        RECT 1250.840 1635.440 1251.100 1635.700 ;
        RECT 1250.840 1586.820 1251.100 1587.080 ;
        RECT 1250.840 1562.680 1251.100 1562.940 ;
        RECT 1250.380 1400.500 1250.640 1400.760 ;
        RECT 1250.840 1400.500 1251.100 1400.760 ;
        RECT 1250.380 1369.560 1250.640 1369.820 ;
        RECT 1251.300 1369.560 1251.560 1369.820 ;
        RECT 1250.840 1321.280 1251.100 1321.540 ;
        RECT 1250.840 1297.140 1251.100 1297.400 ;
        RECT 1250.840 1255.660 1251.100 1255.920 ;
        RECT 1250.840 1207.380 1251.100 1207.640 ;
        RECT 1250.380 1173.040 1250.640 1173.300 ;
        RECT 1250.840 1152.300 1251.100 1152.560 ;
        RECT 1250.380 1062.540 1250.640 1062.800 ;
        RECT 1251.300 1062.540 1251.560 1062.800 ;
        RECT 1249.920 1055.400 1250.180 1055.660 ;
        RECT 1250.380 1055.400 1250.640 1055.660 ;
        RECT 1250.380 1007.120 1250.640 1007.380 ;
        RECT 1250.840 1007.120 1251.100 1007.380 ;
        RECT 1250.380 1000.320 1250.640 1000.580 ;
        RECT 1251.300 1000.320 1251.560 1000.580 ;
        RECT 1251.300 883.700 1251.560 883.960 ;
        RECT 1250.380 883.360 1250.640 883.620 ;
        RECT 1250.840 814.000 1251.100 814.260 ;
        RECT 1251.300 814.000 1251.560 814.260 ;
        RECT 1250.840 717.440 1251.100 717.700 ;
        RECT 1250.840 689.560 1251.100 689.820 ;
        RECT 1250.840 282.920 1251.100 283.180 ;
        RECT 1250.840 268.980 1251.100 269.240 ;
        RECT 1250.840 234.980 1251.100 235.240 ;
        RECT 1250.380 234.300 1250.640 234.560 ;
        RECT 1249.920 179.560 1250.180 179.820 ;
        RECT 1250.380 179.560 1250.640 179.820 ;
        RECT 1250.380 178.880 1250.640 179.140 ;
        RECT 1250.840 131.280 1251.100 131.540 ;
        RECT 1250.840 110.540 1251.100 110.800 ;
        RECT 1249.920 83.000 1250.180 83.260 ;
      LAYER met2 ;
        RECT 1254.905 1700.410 1255.185 1704.000 ;
        RECT 1253.200 1700.270 1255.185 1700.410 ;
        RECT 1253.200 1677.890 1253.340 1700.270 ;
        RECT 1254.905 1700.000 1255.185 1700.270 ;
        RECT 1253.140 1677.570 1253.400 1677.890 ;
        RECT 1250.840 1635.410 1251.100 1635.730 ;
        RECT 1250.900 1587.110 1251.040 1635.410 ;
        RECT 1250.840 1586.790 1251.100 1587.110 ;
        RECT 1250.840 1562.650 1251.100 1562.970 ;
        RECT 1250.900 1400.790 1251.040 1562.650 ;
        RECT 1250.380 1400.470 1250.640 1400.790 ;
        RECT 1250.840 1400.470 1251.100 1400.790 ;
        RECT 1250.440 1369.850 1250.580 1400.470 ;
        RECT 1250.380 1369.530 1250.640 1369.850 ;
        RECT 1251.300 1369.530 1251.560 1369.850 ;
        RECT 1251.360 1345.450 1251.500 1369.530 ;
        RECT 1250.900 1345.310 1251.500 1345.450 ;
        RECT 1250.900 1321.570 1251.040 1345.310 ;
        RECT 1250.840 1321.250 1251.100 1321.570 ;
        RECT 1250.840 1297.110 1251.100 1297.430 ;
        RECT 1250.900 1255.950 1251.040 1297.110 ;
        RECT 1250.840 1255.630 1251.100 1255.950 ;
        RECT 1250.840 1207.350 1251.100 1207.670 ;
        RECT 1250.900 1200.610 1251.040 1207.350 ;
        RECT 1250.440 1200.470 1251.040 1200.610 ;
        RECT 1250.440 1173.330 1250.580 1200.470 ;
        RECT 1250.380 1173.010 1250.640 1173.330 ;
        RECT 1250.840 1152.270 1251.100 1152.590 ;
        RECT 1250.900 1087.050 1251.040 1152.270 ;
        RECT 1250.900 1086.910 1251.500 1087.050 ;
        RECT 1251.360 1062.830 1251.500 1086.910 ;
        RECT 1250.380 1062.510 1250.640 1062.830 ;
        RECT 1251.300 1062.510 1251.560 1062.830 ;
        RECT 1250.440 1055.690 1250.580 1062.510 ;
        RECT 1249.920 1055.370 1250.180 1055.690 ;
        RECT 1250.380 1055.370 1250.640 1055.690 ;
        RECT 1249.980 1007.605 1250.120 1055.370 ;
        RECT 1249.910 1007.235 1250.190 1007.605 ;
        RECT 1250.380 1007.090 1250.640 1007.410 ;
        RECT 1250.830 1007.235 1251.110 1007.605 ;
        RECT 1250.840 1007.090 1251.100 1007.235 ;
        RECT 1250.440 1000.610 1250.580 1007.090 ;
        RECT 1250.380 1000.290 1250.640 1000.610 ;
        RECT 1251.300 1000.290 1251.560 1000.610 ;
        RECT 1251.360 883.990 1251.500 1000.290 ;
        RECT 1251.300 883.670 1251.560 883.990 ;
        RECT 1250.380 883.330 1250.640 883.650 ;
        RECT 1250.440 821.170 1250.580 883.330 ;
        RECT 1250.440 821.030 1251.040 821.170 ;
        RECT 1250.900 814.290 1251.040 821.030 ;
        RECT 1250.840 813.970 1251.100 814.290 ;
        RECT 1251.300 813.970 1251.560 814.290 ;
        RECT 1251.360 747.730 1251.500 813.970 ;
        RECT 1250.900 747.590 1251.500 747.730 ;
        RECT 1250.900 717.730 1251.040 747.590 ;
        RECT 1250.840 717.410 1251.100 717.730 ;
        RECT 1250.840 689.530 1251.100 689.850 ;
        RECT 1250.900 580.565 1251.040 689.530 ;
        RECT 1250.830 580.195 1251.110 580.565 ;
        RECT 1250.370 579.515 1250.650 579.885 ;
        RECT 1250.440 555.290 1250.580 579.515 ;
        RECT 1250.440 555.150 1251.040 555.290 ;
        RECT 1250.900 507.010 1251.040 555.150 ;
        RECT 1250.440 506.870 1251.040 507.010 ;
        RECT 1250.440 362.170 1250.580 506.870 ;
        RECT 1250.440 362.030 1251.040 362.170 ;
        RECT 1250.900 283.210 1251.040 362.030 ;
        RECT 1250.840 282.890 1251.100 283.210 ;
        RECT 1250.840 268.950 1251.100 269.270 ;
        RECT 1250.900 235.270 1251.040 268.950 ;
        RECT 1250.840 234.950 1251.100 235.270 ;
        RECT 1250.380 234.270 1250.640 234.590 ;
        RECT 1250.440 227.530 1250.580 234.270 ;
        RECT 1249.980 227.390 1250.580 227.530 ;
        RECT 1249.980 179.850 1250.120 227.390 ;
        RECT 1249.920 179.530 1250.180 179.850 ;
        RECT 1250.380 179.530 1250.640 179.850 ;
        RECT 1250.440 179.170 1250.580 179.530 ;
        RECT 1250.380 178.850 1250.640 179.170 ;
        RECT 1250.840 131.250 1251.100 131.570 ;
        RECT 1250.900 110.830 1251.040 131.250 ;
        RECT 1250.840 110.510 1251.100 110.830 ;
        RECT 1249.920 82.970 1250.180 83.290 ;
        RECT 1249.980 31.125 1250.120 82.970 ;
        RECT 258.150 30.755 258.430 31.125 ;
        RECT 1249.910 30.755 1250.190 31.125 ;
        RECT 258.220 2.400 258.360 30.755 ;
        RECT 258.010 -4.800 258.570 2.400 ;
      LAYER via2 ;
        RECT 1249.910 1007.280 1250.190 1007.560 ;
        RECT 1250.830 1007.280 1251.110 1007.560 ;
        RECT 1250.830 580.240 1251.110 580.520 ;
        RECT 1250.370 579.560 1250.650 579.840 ;
        RECT 258.150 30.800 258.430 31.080 ;
        RECT 1249.910 30.800 1250.190 31.080 ;
      LAYER met3 ;
        RECT 1249.885 1007.570 1250.215 1007.585 ;
        RECT 1250.805 1007.570 1251.135 1007.585 ;
        RECT 1249.885 1007.270 1251.135 1007.570 ;
        RECT 1249.885 1007.255 1250.215 1007.270 ;
        RECT 1250.805 1007.255 1251.135 1007.270 ;
        RECT 1250.805 580.530 1251.135 580.545 ;
        RECT 1250.590 580.215 1251.135 580.530 ;
        RECT 1250.590 579.865 1250.890 580.215 ;
        RECT 1250.345 579.550 1250.890 579.865 ;
        RECT 1250.345 579.535 1250.675 579.550 ;
        RECT 258.125 31.090 258.455 31.105 ;
        RECT 1249.885 31.090 1250.215 31.105 ;
        RECT 258.125 30.790 1250.215 31.090 ;
        RECT 258.125 30.775 258.455 30.790 ;
        RECT 1249.885 30.775 1250.215 30.790 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1257.785 1538.925 1257.955 1587.035 ;
        RECT 1256.865 1442.025 1257.035 1490.475 ;
        RECT 1256.865 662.405 1257.035 710.515 ;
        RECT 1256.865 565.845 1257.035 613.955 ;
        RECT 1256.865 324.445 1257.035 386.155 ;
        RECT 1256.865 179.605 1257.035 227.715 ;
      LAYER mcon ;
        RECT 1257.785 1586.865 1257.955 1587.035 ;
        RECT 1256.865 1490.305 1257.035 1490.475 ;
        RECT 1256.865 710.345 1257.035 710.515 ;
        RECT 1256.865 613.785 1257.035 613.955 ;
        RECT 1256.865 385.985 1257.035 386.155 ;
        RECT 1256.865 227.545 1257.035 227.715 ;
      LAYER met1 ;
        RECT 1257.710 1587.020 1258.030 1587.080 ;
        RECT 1257.515 1586.880 1258.030 1587.020 ;
        RECT 1257.710 1586.820 1258.030 1586.880 ;
        RECT 1257.710 1539.080 1258.030 1539.140 ;
        RECT 1257.515 1538.940 1258.030 1539.080 ;
        RECT 1257.710 1538.880 1258.030 1538.940 ;
        RECT 1256.805 1490.460 1257.095 1490.505 ;
        RECT 1257.710 1490.460 1258.030 1490.520 ;
        RECT 1256.805 1490.320 1258.030 1490.460 ;
        RECT 1256.805 1490.275 1257.095 1490.320 ;
        RECT 1257.710 1490.260 1258.030 1490.320 ;
        RECT 1256.790 1442.180 1257.110 1442.240 ;
        RECT 1256.595 1442.040 1257.110 1442.180 ;
        RECT 1256.790 1441.980 1257.110 1442.040 ;
        RECT 1255.870 1352.760 1256.190 1352.820 ;
        RECT 1257.250 1352.760 1257.570 1352.820 ;
        RECT 1255.870 1352.620 1257.570 1352.760 ;
        RECT 1255.870 1352.560 1256.190 1352.620 ;
        RECT 1257.250 1352.560 1257.570 1352.620 ;
        RECT 1255.870 1256.200 1256.190 1256.260 ;
        RECT 1257.250 1256.200 1257.570 1256.260 ;
        RECT 1255.870 1256.060 1257.570 1256.200 ;
        RECT 1255.870 1256.000 1256.190 1256.060 ;
        RECT 1257.250 1256.000 1257.570 1256.060 ;
        RECT 1255.870 1200.780 1256.190 1200.840 ;
        RECT 1256.790 1200.780 1257.110 1200.840 ;
        RECT 1255.870 1200.640 1257.110 1200.780 ;
        RECT 1255.870 1200.580 1256.190 1200.640 ;
        RECT 1256.790 1200.580 1257.110 1200.640 ;
        RECT 1255.410 1152.500 1255.730 1152.560 ;
        RECT 1256.790 1152.500 1257.110 1152.560 ;
        RECT 1255.410 1152.360 1257.110 1152.500 ;
        RECT 1255.410 1152.300 1255.730 1152.360 ;
        RECT 1256.790 1152.300 1257.110 1152.360 ;
        RECT 1257.710 1104.220 1258.030 1104.280 ;
        RECT 1258.170 1104.220 1258.490 1104.280 ;
        RECT 1257.710 1104.080 1258.490 1104.220 ;
        RECT 1257.710 1104.020 1258.030 1104.080 ;
        RECT 1258.170 1104.020 1258.490 1104.080 ;
        RECT 1256.790 931.640 1257.110 931.900 ;
        RECT 1256.880 931.220 1257.020 931.640 ;
        RECT 1256.790 930.960 1257.110 931.220 ;
        RECT 1256.790 917.560 1257.110 917.620 ;
        RECT 1257.710 917.560 1258.030 917.620 ;
        RECT 1256.790 917.420 1258.030 917.560 ;
        RECT 1256.790 917.360 1257.110 917.420 ;
        RECT 1257.710 917.360 1258.030 917.420 ;
        RECT 1255.870 862.820 1256.190 862.880 ;
        RECT 1257.710 862.820 1258.030 862.880 ;
        RECT 1255.870 862.680 1258.030 862.820 ;
        RECT 1255.870 862.620 1256.190 862.680 ;
        RECT 1257.710 862.620 1258.030 862.680 ;
        RECT 1255.870 821.140 1256.190 821.400 ;
        RECT 1255.960 820.660 1256.100 821.140 ;
        RECT 1256.790 820.660 1257.110 820.720 ;
        RECT 1255.960 820.520 1257.110 820.660 ;
        RECT 1256.790 820.460 1257.110 820.520 ;
        RECT 1256.790 814.200 1257.110 814.260 ;
        RECT 1258.170 814.200 1258.490 814.260 ;
        RECT 1256.790 814.060 1258.490 814.200 ;
        RECT 1256.790 814.000 1257.110 814.060 ;
        RECT 1258.170 814.000 1258.490 814.060 ;
        RECT 1256.790 718.320 1257.110 718.380 ;
        RECT 1257.710 718.320 1258.030 718.380 ;
        RECT 1256.790 718.180 1258.030 718.320 ;
        RECT 1256.790 718.120 1257.110 718.180 ;
        RECT 1257.710 718.120 1258.030 718.180 ;
        RECT 1256.790 710.500 1257.110 710.560 ;
        RECT 1256.595 710.360 1257.110 710.500 ;
        RECT 1256.790 710.300 1257.110 710.360 ;
        RECT 1256.805 662.560 1257.095 662.605 ;
        RECT 1257.250 662.560 1257.570 662.620 ;
        RECT 1256.805 662.420 1257.570 662.560 ;
        RECT 1256.805 662.375 1257.095 662.420 ;
        RECT 1257.250 662.360 1257.570 662.420 ;
        RECT 1256.790 613.940 1257.110 614.000 ;
        RECT 1256.595 613.800 1257.110 613.940 ;
        RECT 1256.790 613.740 1257.110 613.800 ;
        RECT 1256.805 566.000 1257.095 566.045 ;
        RECT 1257.250 566.000 1257.570 566.060 ;
        RECT 1256.805 565.860 1257.570 566.000 ;
        RECT 1256.805 565.815 1257.095 565.860 ;
        RECT 1257.250 565.800 1257.570 565.860 ;
        RECT 1256.805 386.140 1257.095 386.185 ;
        RECT 1257.250 386.140 1257.570 386.200 ;
        RECT 1256.805 386.000 1257.570 386.140 ;
        RECT 1256.805 385.955 1257.095 386.000 ;
        RECT 1257.250 385.940 1257.570 386.000 ;
        RECT 1256.790 324.600 1257.110 324.660 ;
        RECT 1256.595 324.460 1257.110 324.600 ;
        RECT 1256.790 324.400 1257.110 324.460 ;
        RECT 1256.790 227.700 1257.110 227.760 ;
        RECT 1256.595 227.560 1257.110 227.700 ;
        RECT 1256.790 227.500 1257.110 227.560 ;
        RECT 1256.805 179.760 1257.095 179.805 ;
        RECT 1257.250 179.760 1257.570 179.820 ;
        RECT 1256.805 179.620 1257.570 179.760 ;
        RECT 1256.805 179.575 1257.095 179.620 ;
        RECT 1257.250 179.560 1257.570 179.620 ;
        RECT 1256.790 96.800 1257.110 96.860 ;
        RECT 1257.710 96.800 1258.030 96.860 ;
        RECT 1256.790 96.660 1258.030 96.800 ;
        RECT 1256.790 96.600 1257.110 96.660 ;
        RECT 1257.710 96.600 1258.030 96.660 ;
        RECT 276.070 30.840 276.390 30.900 ;
        RECT 1257.250 30.840 1257.570 30.900 ;
        RECT 276.070 30.700 1257.570 30.840 ;
        RECT 276.070 30.640 276.390 30.700 ;
        RECT 1257.250 30.640 1257.570 30.700 ;
      LAYER via ;
        RECT 1257.740 1586.820 1258.000 1587.080 ;
        RECT 1257.740 1538.880 1258.000 1539.140 ;
        RECT 1257.740 1490.260 1258.000 1490.520 ;
        RECT 1256.820 1441.980 1257.080 1442.240 ;
        RECT 1255.900 1352.560 1256.160 1352.820 ;
        RECT 1257.280 1352.560 1257.540 1352.820 ;
        RECT 1255.900 1256.000 1256.160 1256.260 ;
        RECT 1257.280 1256.000 1257.540 1256.260 ;
        RECT 1255.900 1200.580 1256.160 1200.840 ;
        RECT 1256.820 1200.580 1257.080 1200.840 ;
        RECT 1255.440 1152.300 1255.700 1152.560 ;
        RECT 1256.820 1152.300 1257.080 1152.560 ;
        RECT 1257.740 1104.020 1258.000 1104.280 ;
        RECT 1258.200 1104.020 1258.460 1104.280 ;
        RECT 1256.820 931.640 1257.080 931.900 ;
        RECT 1256.820 930.960 1257.080 931.220 ;
        RECT 1256.820 917.360 1257.080 917.620 ;
        RECT 1257.740 917.360 1258.000 917.620 ;
        RECT 1255.900 862.620 1256.160 862.880 ;
        RECT 1257.740 862.620 1258.000 862.880 ;
        RECT 1255.900 821.140 1256.160 821.400 ;
        RECT 1256.820 820.460 1257.080 820.720 ;
        RECT 1256.820 814.000 1257.080 814.260 ;
        RECT 1258.200 814.000 1258.460 814.260 ;
        RECT 1256.820 718.120 1257.080 718.380 ;
        RECT 1257.740 718.120 1258.000 718.380 ;
        RECT 1256.820 710.300 1257.080 710.560 ;
        RECT 1257.280 662.360 1257.540 662.620 ;
        RECT 1256.820 613.740 1257.080 614.000 ;
        RECT 1257.280 565.800 1257.540 566.060 ;
        RECT 1257.280 385.940 1257.540 386.200 ;
        RECT 1256.820 324.400 1257.080 324.660 ;
        RECT 1256.820 227.500 1257.080 227.760 ;
        RECT 1257.280 179.560 1257.540 179.820 ;
        RECT 1256.820 96.600 1257.080 96.860 ;
        RECT 1257.740 96.600 1258.000 96.860 ;
        RECT 276.100 30.640 276.360 30.900 ;
        RECT 1257.280 30.640 1257.540 30.900 ;
      LAYER met2 ;
        RECT 1262.265 1700.410 1262.545 1704.000 ;
        RECT 1260.560 1700.270 1262.545 1700.410 ;
        RECT 1260.560 1678.650 1260.700 1700.270 ;
        RECT 1262.265 1700.000 1262.545 1700.270 ;
        RECT 1257.340 1678.510 1260.700 1678.650 ;
        RECT 1257.340 1618.130 1257.480 1678.510 ;
        RECT 1257.340 1617.990 1257.940 1618.130 ;
        RECT 1257.800 1587.110 1257.940 1617.990 ;
        RECT 1257.740 1586.790 1258.000 1587.110 ;
        RECT 1257.740 1538.850 1258.000 1539.170 ;
        RECT 1257.800 1538.685 1257.940 1538.850 ;
        RECT 1257.730 1538.315 1258.010 1538.685 ;
        RECT 1257.730 1490.715 1258.010 1491.085 ;
        RECT 1257.800 1490.550 1257.940 1490.715 ;
        RECT 1257.740 1490.230 1258.000 1490.550 ;
        RECT 1256.820 1441.950 1257.080 1442.270 ;
        RECT 1256.880 1400.645 1257.020 1441.950 ;
        RECT 1255.890 1400.275 1256.170 1400.645 ;
        RECT 1256.810 1400.275 1257.090 1400.645 ;
        RECT 1255.960 1352.850 1256.100 1400.275 ;
        RECT 1255.900 1352.530 1256.160 1352.850 ;
        RECT 1257.280 1352.530 1257.540 1352.850 ;
        RECT 1257.340 1328.450 1257.480 1352.530 ;
        RECT 1257.340 1328.310 1257.940 1328.450 ;
        RECT 1257.800 1317.570 1257.940 1328.310 ;
        RECT 1256.880 1317.430 1257.940 1317.570 ;
        RECT 1256.880 1304.085 1257.020 1317.430 ;
        RECT 1255.890 1303.715 1256.170 1304.085 ;
        RECT 1256.810 1303.715 1257.090 1304.085 ;
        RECT 1255.960 1256.290 1256.100 1303.715 ;
        RECT 1255.900 1255.970 1256.160 1256.290 ;
        RECT 1257.280 1255.970 1257.540 1256.290 ;
        RECT 1257.340 1249.005 1257.480 1255.970 ;
        RECT 1255.890 1248.635 1256.170 1249.005 ;
        RECT 1257.270 1248.635 1257.550 1249.005 ;
        RECT 1255.960 1200.870 1256.100 1248.635 ;
        RECT 1255.430 1200.355 1255.710 1200.725 ;
        RECT 1255.900 1200.550 1256.160 1200.870 ;
        RECT 1256.820 1200.725 1257.080 1200.870 ;
        RECT 1256.810 1200.355 1257.090 1200.725 ;
        RECT 1255.500 1152.590 1255.640 1200.355 ;
        RECT 1255.440 1152.270 1255.700 1152.590 ;
        RECT 1256.820 1152.445 1257.080 1152.590 ;
        RECT 1256.810 1152.075 1257.090 1152.445 ;
        RECT 1257.730 1152.075 1258.010 1152.445 ;
        RECT 1257.800 1104.310 1257.940 1152.075 ;
        RECT 1257.740 1103.990 1258.000 1104.310 ;
        RECT 1258.200 1103.990 1258.460 1104.310 ;
        RECT 1258.260 1062.570 1258.400 1103.990 ;
        RECT 1257.800 1062.430 1258.400 1062.570 ;
        RECT 1257.800 1027.890 1257.940 1062.430 ;
        RECT 1257.340 1027.750 1257.940 1027.890 ;
        RECT 1257.340 1013.610 1257.480 1027.750 ;
        RECT 1257.340 1013.470 1257.940 1013.610 ;
        RECT 1257.800 966.125 1257.940 1013.470 ;
        RECT 1256.810 965.755 1257.090 966.125 ;
        RECT 1257.730 965.755 1258.010 966.125 ;
        RECT 1256.880 931.930 1257.020 965.755 ;
        RECT 1256.820 931.610 1257.080 931.930 ;
        RECT 1256.820 930.930 1257.080 931.250 ;
        RECT 1256.880 917.650 1257.020 930.930 ;
        RECT 1256.820 917.330 1257.080 917.650 ;
        RECT 1257.740 917.330 1258.000 917.650 ;
        RECT 1257.800 862.910 1257.940 917.330 ;
        RECT 1255.900 862.590 1256.160 862.910 ;
        RECT 1257.740 862.590 1258.000 862.910 ;
        RECT 1255.960 821.430 1256.100 862.590 ;
        RECT 1255.900 821.110 1256.160 821.430 ;
        RECT 1256.820 820.430 1257.080 820.750 ;
        RECT 1256.880 814.290 1257.020 820.430 ;
        RECT 1256.820 813.970 1257.080 814.290 ;
        RECT 1258.200 813.970 1258.460 814.290 ;
        RECT 1258.260 772.210 1258.400 813.970 ;
        RECT 1257.800 772.070 1258.400 772.210 ;
        RECT 1257.800 718.410 1257.940 772.070 ;
        RECT 1256.820 718.090 1257.080 718.410 ;
        RECT 1257.740 718.090 1258.000 718.410 ;
        RECT 1256.880 710.590 1257.020 718.090 ;
        RECT 1256.820 710.270 1257.080 710.590 ;
        RECT 1257.280 662.330 1257.540 662.650 ;
        RECT 1257.340 621.250 1257.480 662.330 ;
        RECT 1256.880 621.110 1257.480 621.250 ;
        RECT 1256.880 614.030 1257.020 621.110 ;
        RECT 1256.820 613.710 1257.080 614.030 ;
        RECT 1257.280 565.770 1257.540 566.090 ;
        RECT 1257.340 388.010 1257.480 565.770 ;
        RECT 1257.340 387.870 1258.400 388.010 ;
        RECT 1258.260 386.765 1258.400 387.870 ;
        RECT 1257.270 386.395 1257.550 386.765 ;
        RECT 1258.190 386.395 1258.470 386.765 ;
        RECT 1257.340 386.230 1257.480 386.395 ;
        RECT 1257.280 385.910 1257.540 386.230 ;
        RECT 1256.820 324.370 1257.080 324.690 ;
        RECT 1256.880 227.790 1257.020 324.370 ;
        RECT 1256.820 227.470 1257.080 227.790 ;
        RECT 1257.280 179.530 1257.540 179.850 ;
        RECT 1257.340 144.570 1257.480 179.530 ;
        RECT 1257.340 144.430 1257.940 144.570 ;
        RECT 1257.800 96.890 1257.940 144.430 ;
        RECT 1256.820 96.570 1257.080 96.890 ;
        RECT 1257.740 96.570 1258.000 96.890 ;
        RECT 1256.880 96.405 1257.020 96.570 ;
        RECT 1256.810 96.035 1257.090 96.405 ;
        RECT 1258.190 95.355 1258.470 95.725 ;
        RECT 1258.260 48.805 1258.400 95.355 ;
        RECT 1257.270 48.435 1257.550 48.805 ;
        RECT 1258.190 48.435 1258.470 48.805 ;
        RECT 1257.340 30.930 1257.480 48.435 ;
        RECT 276.100 30.610 276.360 30.930 ;
        RECT 1257.280 30.610 1257.540 30.930 ;
        RECT 276.160 2.400 276.300 30.610 ;
        RECT 275.950 -4.800 276.510 2.400 ;
      LAYER via2 ;
        RECT 1257.730 1538.360 1258.010 1538.640 ;
        RECT 1257.730 1490.760 1258.010 1491.040 ;
        RECT 1255.890 1400.320 1256.170 1400.600 ;
        RECT 1256.810 1400.320 1257.090 1400.600 ;
        RECT 1255.890 1303.760 1256.170 1304.040 ;
        RECT 1256.810 1303.760 1257.090 1304.040 ;
        RECT 1255.890 1248.680 1256.170 1248.960 ;
        RECT 1257.270 1248.680 1257.550 1248.960 ;
        RECT 1255.430 1200.400 1255.710 1200.680 ;
        RECT 1256.810 1200.400 1257.090 1200.680 ;
        RECT 1256.810 1152.120 1257.090 1152.400 ;
        RECT 1257.730 1152.120 1258.010 1152.400 ;
        RECT 1256.810 965.800 1257.090 966.080 ;
        RECT 1257.730 965.800 1258.010 966.080 ;
        RECT 1257.270 386.440 1257.550 386.720 ;
        RECT 1258.190 386.440 1258.470 386.720 ;
        RECT 1256.810 96.080 1257.090 96.360 ;
        RECT 1258.190 95.400 1258.470 95.680 ;
        RECT 1257.270 48.480 1257.550 48.760 ;
        RECT 1258.190 48.480 1258.470 48.760 ;
      LAYER met3 ;
        RECT 1256.990 1538.650 1257.370 1538.660 ;
        RECT 1257.705 1538.650 1258.035 1538.665 ;
        RECT 1256.990 1538.350 1258.035 1538.650 ;
        RECT 1256.990 1538.340 1257.370 1538.350 ;
        RECT 1257.705 1538.335 1258.035 1538.350 ;
        RECT 1256.990 1491.050 1257.370 1491.060 ;
        RECT 1257.705 1491.050 1258.035 1491.065 ;
        RECT 1256.990 1490.750 1258.035 1491.050 ;
        RECT 1256.990 1490.740 1257.370 1490.750 ;
        RECT 1257.705 1490.735 1258.035 1490.750 ;
        RECT 1255.865 1400.610 1256.195 1400.625 ;
        RECT 1256.785 1400.610 1257.115 1400.625 ;
        RECT 1255.865 1400.310 1257.115 1400.610 ;
        RECT 1255.865 1400.295 1256.195 1400.310 ;
        RECT 1256.785 1400.295 1257.115 1400.310 ;
        RECT 1255.865 1304.050 1256.195 1304.065 ;
        RECT 1256.785 1304.050 1257.115 1304.065 ;
        RECT 1255.865 1303.750 1257.115 1304.050 ;
        RECT 1255.865 1303.735 1256.195 1303.750 ;
        RECT 1256.785 1303.735 1257.115 1303.750 ;
        RECT 1255.865 1248.970 1256.195 1248.985 ;
        RECT 1257.245 1248.970 1257.575 1248.985 ;
        RECT 1255.865 1248.670 1257.575 1248.970 ;
        RECT 1255.865 1248.655 1256.195 1248.670 ;
        RECT 1257.245 1248.655 1257.575 1248.670 ;
        RECT 1255.405 1200.690 1255.735 1200.705 ;
        RECT 1256.785 1200.690 1257.115 1200.705 ;
        RECT 1255.405 1200.390 1257.115 1200.690 ;
        RECT 1255.405 1200.375 1255.735 1200.390 ;
        RECT 1256.785 1200.375 1257.115 1200.390 ;
        RECT 1256.785 1152.410 1257.115 1152.425 ;
        RECT 1257.705 1152.410 1258.035 1152.425 ;
        RECT 1256.785 1152.110 1258.035 1152.410 ;
        RECT 1256.785 1152.095 1257.115 1152.110 ;
        RECT 1257.705 1152.095 1258.035 1152.110 ;
        RECT 1256.785 966.090 1257.115 966.105 ;
        RECT 1257.705 966.090 1258.035 966.105 ;
        RECT 1256.785 965.790 1258.035 966.090 ;
        RECT 1256.785 965.775 1257.115 965.790 ;
        RECT 1257.705 965.775 1258.035 965.790 ;
        RECT 1257.245 386.730 1257.575 386.745 ;
        RECT 1258.165 386.730 1258.495 386.745 ;
        RECT 1257.245 386.430 1258.495 386.730 ;
        RECT 1257.245 386.415 1257.575 386.430 ;
        RECT 1258.165 386.415 1258.495 386.430 ;
        RECT 1256.785 96.370 1257.115 96.385 ;
        RECT 1256.110 96.070 1257.115 96.370 ;
        RECT 1256.110 95.690 1256.410 96.070 ;
        RECT 1256.785 96.055 1257.115 96.070 ;
        RECT 1258.165 95.690 1258.495 95.705 ;
        RECT 1256.110 95.390 1258.495 95.690 ;
        RECT 1258.165 95.375 1258.495 95.390 ;
        RECT 1257.245 48.770 1257.575 48.785 ;
        RECT 1258.165 48.770 1258.495 48.785 ;
        RECT 1257.245 48.470 1258.495 48.770 ;
        RECT 1257.245 48.455 1257.575 48.470 ;
        RECT 1258.165 48.455 1258.495 48.470 ;
      LAYER via3 ;
        RECT 1257.020 1538.340 1257.340 1538.660 ;
        RECT 1257.020 1490.740 1257.340 1491.060 ;
      LAYER met4 ;
        RECT 1257.015 1538.335 1257.345 1538.665 ;
        RECT 1257.030 1491.065 1257.330 1538.335 ;
        RECT 1257.015 1490.735 1257.345 1491.065 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 294.010 31.180 294.330 31.240 ;
        RECT 1269.670 31.180 1269.990 31.240 ;
        RECT 294.010 31.040 1269.990 31.180 ;
        RECT 294.010 30.980 294.330 31.040 ;
        RECT 1269.670 30.980 1269.990 31.040 ;
      LAYER via ;
        RECT 294.040 30.980 294.300 31.240 ;
        RECT 1269.700 30.980 1269.960 31.240 ;
      LAYER met2 ;
        RECT 1269.625 1700.000 1269.905 1704.000 ;
        RECT 1269.760 31.270 1269.900 1700.000 ;
        RECT 294.040 30.950 294.300 31.270 ;
        RECT 1269.700 30.950 1269.960 31.270 ;
        RECT 294.100 2.400 294.240 30.950 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 311.950 31.520 312.270 31.580 ;
        RECT 1277.490 31.520 1277.810 31.580 ;
        RECT 311.950 31.380 1277.810 31.520 ;
        RECT 311.950 31.320 312.270 31.380 ;
        RECT 1277.490 31.320 1277.810 31.380 ;
      LAYER via ;
        RECT 311.980 31.320 312.240 31.580 ;
        RECT 1277.520 31.320 1277.780 31.580 ;
      LAYER met2 ;
        RECT 1276.985 1700.410 1277.265 1704.000 ;
        RECT 1276.985 1700.270 1277.720 1700.410 ;
        RECT 1276.985 1700.000 1277.265 1700.270 ;
        RECT 1277.580 31.610 1277.720 1700.270 ;
        RECT 311.980 31.290 312.240 31.610 ;
        RECT 1277.520 31.290 1277.780 31.610 ;
        RECT 312.040 2.400 312.180 31.290 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 31.860 330.210 31.920 ;
        RECT 1283.930 31.860 1284.250 31.920 ;
        RECT 329.890 31.720 1284.250 31.860 ;
        RECT 329.890 31.660 330.210 31.720 ;
        RECT 1283.930 31.660 1284.250 31.720 ;
      LAYER via ;
        RECT 329.920 31.660 330.180 31.920 ;
        RECT 1283.960 31.660 1284.220 31.920 ;
      LAYER met2 ;
        RECT 1284.345 1700.410 1284.625 1704.000 ;
        RECT 1284.020 1700.270 1284.625 1700.410 ;
        RECT 1284.020 31.950 1284.160 1700.270 ;
        RECT 1284.345 1700.000 1284.625 1700.270 ;
        RECT 329.920 31.630 330.180 31.950 ;
        RECT 1283.960 31.630 1284.220 31.950 ;
        RECT 329.980 2.400 330.120 31.630 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 32.200 347.690 32.260 ;
        RECT 1291.290 32.200 1291.610 32.260 ;
        RECT 347.370 32.060 1291.610 32.200 ;
        RECT 347.370 32.000 347.690 32.060 ;
        RECT 1291.290 32.000 1291.610 32.060 ;
      LAYER via ;
        RECT 347.400 32.000 347.660 32.260 ;
        RECT 1291.320 32.000 1291.580 32.260 ;
      LAYER met2 ;
        RECT 1291.705 1700.410 1291.985 1704.000 ;
        RECT 1291.380 1700.270 1291.985 1700.410 ;
        RECT 1291.380 32.290 1291.520 1700.270 ;
        RECT 1291.705 1700.000 1291.985 1700.270 ;
        RECT 347.400 31.970 347.660 32.290 ;
        RECT 1291.320 31.970 1291.580 32.290 ;
        RECT 347.460 2.400 347.600 31.970 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 365.310 32.540 365.630 32.600 ;
        RECT 1297.270 32.540 1297.590 32.600 ;
        RECT 365.310 32.400 1297.590 32.540 ;
        RECT 365.310 32.340 365.630 32.400 ;
        RECT 1297.270 32.340 1297.590 32.400 ;
      LAYER via ;
        RECT 365.340 32.340 365.600 32.600 ;
        RECT 1297.300 32.340 1297.560 32.600 ;
      LAYER met2 ;
        RECT 1299.065 1700.410 1299.345 1704.000 ;
        RECT 1297.360 1700.270 1299.345 1700.410 ;
        RECT 1297.360 32.630 1297.500 1700.270 ;
        RECT 1299.065 1700.000 1299.345 1700.270 ;
        RECT 365.340 32.310 365.600 32.630 ;
        RECT 1297.300 32.310 1297.560 32.630 ;
        RECT 365.400 2.400 365.540 32.310 ;
        RECT 365.190 -4.800 365.750 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 32.880 383.570 32.940 ;
        RECT 1305.090 32.880 1305.410 32.940 ;
        RECT 383.250 32.740 1305.410 32.880 ;
        RECT 383.250 32.680 383.570 32.740 ;
        RECT 1305.090 32.680 1305.410 32.740 ;
      LAYER via ;
        RECT 383.280 32.680 383.540 32.940 ;
        RECT 1305.120 32.680 1305.380 32.940 ;
      LAYER met2 ;
        RECT 1306.425 1700.410 1306.705 1704.000 ;
        RECT 1305.180 1700.270 1306.705 1700.410 ;
        RECT 1305.180 32.970 1305.320 1700.270 ;
        RECT 1306.425 1700.000 1306.705 1700.270 ;
        RECT 383.280 32.650 383.540 32.970 ;
        RECT 1305.120 32.650 1305.380 32.970 ;
        RECT 383.340 2.400 383.480 32.650 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 401.190 40.700 401.510 40.760 ;
        RECT 1311.990 40.700 1312.310 40.760 ;
        RECT 401.190 40.560 1312.310 40.700 ;
        RECT 401.190 40.500 401.510 40.560 ;
        RECT 1311.990 40.500 1312.310 40.560 ;
      LAYER via ;
        RECT 401.220 40.500 401.480 40.760 ;
        RECT 1312.020 40.500 1312.280 40.760 ;
      LAYER met2 ;
        RECT 1313.785 1700.410 1314.065 1704.000 ;
        RECT 1312.080 1700.270 1314.065 1700.410 ;
        RECT 1312.080 40.790 1312.220 1700.270 ;
        RECT 1313.785 1700.000 1314.065 1700.270 ;
        RECT 401.220 40.470 401.480 40.790 ;
        RECT 1312.020 40.470 1312.280 40.790 ;
        RECT 401.280 2.400 401.420 40.470 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 62.170 25.400 62.490 25.460 ;
        RECT 1173.530 25.400 1173.850 25.460 ;
        RECT 62.170 25.260 1173.850 25.400 ;
        RECT 62.170 25.200 62.490 25.260 ;
        RECT 1173.530 25.200 1173.850 25.260 ;
      LAYER via ;
        RECT 62.200 25.200 62.460 25.460 ;
        RECT 1173.560 25.200 1173.820 25.460 ;
      LAYER met2 ;
        RECT 1174.405 1700.410 1174.685 1704.000 ;
        RECT 1173.620 1700.270 1174.685 1700.410 ;
        RECT 1173.620 25.490 1173.760 1700.270 ;
        RECT 1174.405 1700.000 1174.685 1700.270 ;
        RECT 62.200 25.170 62.460 25.490 ;
        RECT 1173.560 25.170 1173.820 25.490 ;
        RECT 62.260 2.400 62.400 25.170 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 41.040 419.450 41.100 ;
        RECT 1319.350 41.040 1319.670 41.100 ;
        RECT 419.130 40.900 1319.670 41.040 ;
        RECT 419.130 40.840 419.450 40.900 ;
        RECT 1319.350 40.840 1319.670 40.900 ;
      LAYER via ;
        RECT 419.160 40.840 419.420 41.100 ;
        RECT 1319.380 40.840 1319.640 41.100 ;
      LAYER met2 ;
        RECT 1321.145 1700.410 1321.425 1704.000 ;
        RECT 1319.440 1700.270 1321.425 1700.410 ;
        RECT 1319.440 41.130 1319.580 1700.270 ;
        RECT 1321.145 1700.000 1321.425 1700.270 ;
        RECT 419.160 40.810 419.420 41.130 ;
        RECT 1319.380 40.810 1319.640 41.130 ;
        RECT 419.220 2.400 419.360 40.810 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1326.325 1587.205 1326.495 1635.315 ;
        RECT 1326.325 1500.505 1326.495 1545.555 ;
        RECT 1326.785 752.165 1326.955 800.275 ;
        RECT 1326.325 462.485 1326.495 476.595 ;
        RECT 1326.325 254.405 1326.495 331.075 ;
        RECT 1325.865 186.405 1326.035 234.515 ;
        RECT 1326.325 90.185 1326.495 137.955 ;
      LAYER mcon ;
        RECT 1326.325 1635.145 1326.495 1635.315 ;
        RECT 1326.325 1545.385 1326.495 1545.555 ;
        RECT 1326.785 800.105 1326.955 800.275 ;
        RECT 1326.325 476.425 1326.495 476.595 ;
        RECT 1326.325 330.905 1326.495 331.075 ;
        RECT 1325.865 234.345 1326.035 234.515 ;
        RECT 1326.325 137.785 1326.495 137.955 ;
      LAYER met1 ;
        RECT 1326.250 1642.100 1326.570 1642.160 ;
        RECT 1326.710 1642.100 1327.030 1642.160 ;
        RECT 1326.250 1641.960 1327.030 1642.100 ;
        RECT 1326.250 1641.900 1326.570 1641.960 ;
        RECT 1326.710 1641.900 1327.030 1641.960 ;
        RECT 1326.265 1635.300 1326.555 1635.345 ;
        RECT 1326.710 1635.300 1327.030 1635.360 ;
        RECT 1326.265 1635.160 1327.030 1635.300 ;
        RECT 1326.265 1635.115 1326.555 1635.160 ;
        RECT 1326.710 1635.100 1327.030 1635.160 ;
        RECT 1326.250 1587.360 1326.570 1587.420 ;
        RECT 1326.055 1587.220 1326.570 1587.360 ;
        RECT 1326.250 1587.160 1326.570 1587.220 ;
        RECT 1326.250 1545.540 1326.570 1545.600 ;
        RECT 1326.055 1545.400 1326.570 1545.540 ;
        RECT 1326.250 1545.340 1326.570 1545.400 ;
        RECT 1326.265 1500.660 1326.555 1500.705 ;
        RECT 1326.710 1500.660 1327.030 1500.720 ;
        RECT 1326.265 1500.520 1327.030 1500.660 ;
        RECT 1326.265 1500.475 1326.555 1500.520 ;
        RECT 1326.710 1500.460 1327.030 1500.520 ;
        RECT 1326.710 1469.720 1327.030 1469.780 ;
        RECT 1327.630 1469.720 1327.950 1469.780 ;
        RECT 1326.710 1469.580 1327.950 1469.720 ;
        RECT 1326.710 1469.520 1327.030 1469.580 ;
        RECT 1327.630 1469.520 1327.950 1469.580 ;
        RECT 1326.250 1345.420 1326.570 1345.680 ;
        RECT 1325.790 1345.280 1326.110 1345.340 ;
        RECT 1326.340 1345.280 1326.480 1345.420 ;
        RECT 1325.790 1345.140 1326.480 1345.280 ;
        RECT 1325.790 1345.080 1326.110 1345.140 ;
        RECT 1325.790 1111.020 1326.110 1111.080 ;
        RECT 1326.710 1111.020 1327.030 1111.080 ;
        RECT 1325.790 1110.880 1327.030 1111.020 ;
        RECT 1325.790 1110.820 1326.110 1110.880 ;
        RECT 1326.710 1110.820 1327.030 1110.880 ;
        RECT 1326.250 966.180 1326.570 966.240 ;
        RECT 1326.710 966.180 1327.030 966.240 ;
        RECT 1326.250 966.040 1327.030 966.180 ;
        RECT 1326.250 965.980 1326.570 966.040 ;
        RECT 1326.710 965.980 1327.030 966.040 ;
        RECT 1324.870 917.900 1325.190 917.960 ;
        RECT 1325.790 917.900 1326.110 917.960 ;
        RECT 1324.870 917.760 1326.110 917.900 ;
        RECT 1324.870 917.700 1325.190 917.760 ;
        RECT 1325.790 917.700 1326.110 917.760 ;
        RECT 1326.250 869.620 1326.570 869.680 ;
        RECT 1326.710 869.620 1327.030 869.680 ;
        RECT 1326.250 869.480 1327.030 869.620 ;
        RECT 1326.250 869.420 1326.570 869.480 ;
        RECT 1326.710 869.420 1327.030 869.480 ;
        RECT 1325.790 807.400 1326.110 807.460 ;
        RECT 1326.250 807.400 1326.570 807.460 ;
        RECT 1325.790 807.260 1326.570 807.400 ;
        RECT 1325.790 807.200 1326.110 807.260 ;
        RECT 1326.250 807.200 1326.570 807.260 ;
        RECT 1325.790 800.260 1326.110 800.320 ;
        RECT 1326.725 800.260 1327.015 800.305 ;
        RECT 1325.790 800.120 1327.015 800.260 ;
        RECT 1325.790 800.060 1326.110 800.120 ;
        RECT 1326.725 800.075 1327.015 800.120 ;
        RECT 1326.710 752.320 1327.030 752.380 ;
        RECT 1326.515 752.180 1327.030 752.320 ;
        RECT 1326.710 752.120 1327.030 752.180 ;
        RECT 1325.790 572.800 1326.110 572.860 ;
        RECT 1326.250 572.800 1326.570 572.860 ;
        RECT 1325.790 572.660 1326.570 572.800 ;
        RECT 1325.790 572.600 1326.110 572.660 ;
        RECT 1326.250 572.600 1326.570 572.660 ;
        RECT 1325.790 545.060 1326.110 545.320 ;
        RECT 1325.880 544.920 1326.020 545.060 ;
        RECT 1326.250 544.920 1326.570 544.980 ;
        RECT 1325.880 544.780 1326.570 544.920 ;
        RECT 1326.250 544.720 1326.570 544.780 ;
        RECT 1326.250 476.580 1326.570 476.640 ;
        RECT 1326.055 476.440 1326.570 476.580 ;
        RECT 1326.250 476.380 1326.570 476.440 ;
        RECT 1326.250 462.640 1326.570 462.700 ;
        RECT 1326.055 462.500 1326.570 462.640 ;
        RECT 1326.250 462.440 1326.570 462.500 ;
        RECT 1325.790 338.200 1326.110 338.260 ;
        RECT 1326.250 338.200 1326.570 338.260 ;
        RECT 1325.790 338.060 1326.570 338.200 ;
        RECT 1325.790 338.000 1326.110 338.060 ;
        RECT 1326.250 338.000 1326.570 338.060 ;
        RECT 1325.790 331.060 1326.110 331.120 ;
        RECT 1326.265 331.060 1326.555 331.105 ;
        RECT 1325.790 330.920 1326.555 331.060 ;
        RECT 1325.790 330.860 1326.110 330.920 ;
        RECT 1326.265 330.875 1326.555 330.920 ;
        RECT 1325.790 254.560 1326.110 254.620 ;
        RECT 1326.265 254.560 1326.555 254.605 ;
        RECT 1325.790 254.420 1326.555 254.560 ;
        RECT 1325.790 254.360 1326.110 254.420 ;
        RECT 1326.265 254.375 1326.555 254.420 ;
        RECT 1325.790 234.500 1326.110 234.560 ;
        RECT 1325.595 234.360 1326.110 234.500 ;
        RECT 1325.790 234.300 1326.110 234.360 ;
        RECT 1325.790 186.560 1326.110 186.620 ;
        RECT 1325.595 186.420 1326.110 186.560 ;
        RECT 1325.790 186.360 1326.110 186.420 ;
        RECT 1325.790 145.080 1326.110 145.140 ;
        RECT 1326.250 145.080 1326.570 145.140 ;
        RECT 1325.790 144.940 1326.570 145.080 ;
        RECT 1325.790 144.880 1326.110 144.940 ;
        RECT 1326.250 144.880 1326.570 144.940 ;
        RECT 1326.250 137.940 1326.570 138.000 ;
        RECT 1326.055 137.800 1326.570 137.940 ;
        RECT 1326.250 137.740 1326.570 137.800 ;
        RECT 1326.265 90.155 1326.555 90.385 ;
        RECT 1324.870 89.660 1325.190 89.720 ;
        RECT 1326.340 89.660 1326.480 90.155 ;
        RECT 1324.870 89.520 1326.480 89.660 ;
        RECT 1324.870 89.460 1325.190 89.520 ;
        RECT 436.610 41.380 436.930 41.440 ;
        RECT 1325.790 41.380 1326.110 41.440 ;
        RECT 436.610 41.240 1326.110 41.380 ;
        RECT 436.610 41.180 436.930 41.240 ;
        RECT 1325.790 41.180 1326.110 41.240 ;
      LAYER via ;
        RECT 1326.280 1641.900 1326.540 1642.160 ;
        RECT 1326.740 1641.900 1327.000 1642.160 ;
        RECT 1326.740 1635.100 1327.000 1635.360 ;
        RECT 1326.280 1587.160 1326.540 1587.420 ;
        RECT 1326.280 1545.340 1326.540 1545.600 ;
        RECT 1326.740 1500.460 1327.000 1500.720 ;
        RECT 1326.740 1469.520 1327.000 1469.780 ;
        RECT 1327.660 1469.520 1327.920 1469.780 ;
        RECT 1326.280 1345.420 1326.540 1345.680 ;
        RECT 1325.820 1345.080 1326.080 1345.340 ;
        RECT 1325.820 1110.820 1326.080 1111.080 ;
        RECT 1326.740 1110.820 1327.000 1111.080 ;
        RECT 1326.280 965.980 1326.540 966.240 ;
        RECT 1326.740 965.980 1327.000 966.240 ;
        RECT 1324.900 917.700 1325.160 917.960 ;
        RECT 1325.820 917.700 1326.080 917.960 ;
        RECT 1326.280 869.420 1326.540 869.680 ;
        RECT 1326.740 869.420 1327.000 869.680 ;
        RECT 1325.820 807.200 1326.080 807.460 ;
        RECT 1326.280 807.200 1326.540 807.460 ;
        RECT 1325.820 800.060 1326.080 800.320 ;
        RECT 1326.740 752.120 1327.000 752.380 ;
        RECT 1325.820 572.600 1326.080 572.860 ;
        RECT 1326.280 572.600 1326.540 572.860 ;
        RECT 1325.820 545.060 1326.080 545.320 ;
        RECT 1326.280 544.720 1326.540 544.980 ;
        RECT 1326.280 476.380 1326.540 476.640 ;
        RECT 1326.280 462.440 1326.540 462.700 ;
        RECT 1325.820 338.000 1326.080 338.260 ;
        RECT 1326.280 338.000 1326.540 338.260 ;
        RECT 1325.820 330.860 1326.080 331.120 ;
        RECT 1325.820 254.360 1326.080 254.620 ;
        RECT 1325.820 234.300 1326.080 234.560 ;
        RECT 1325.820 186.360 1326.080 186.620 ;
        RECT 1325.820 144.880 1326.080 145.140 ;
        RECT 1326.280 144.880 1326.540 145.140 ;
        RECT 1326.280 137.740 1326.540 138.000 ;
        RECT 1324.900 89.460 1325.160 89.720 ;
        RECT 436.640 41.180 436.900 41.440 ;
        RECT 1325.820 41.180 1326.080 41.440 ;
      LAYER met2 ;
        RECT 1328.505 1700.410 1328.785 1704.000 ;
        RECT 1327.260 1700.270 1328.785 1700.410 ;
        RECT 1327.260 1677.970 1327.400 1700.270 ;
        RECT 1328.505 1700.000 1328.785 1700.270 ;
        RECT 1326.340 1677.830 1327.400 1677.970 ;
        RECT 1326.340 1642.190 1326.480 1677.830 ;
        RECT 1326.280 1641.870 1326.540 1642.190 ;
        RECT 1326.740 1641.870 1327.000 1642.190 ;
        RECT 1326.800 1635.390 1326.940 1641.870 ;
        RECT 1326.740 1635.070 1327.000 1635.390 ;
        RECT 1326.280 1587.130 1326.540 1587.450 ;
        RECT 1326.340 1545.630 1326.480 1587.130 ;
        RECT 1326.280 1545.310 1326.540 1545.630 ;
        RECT 1326.740 1500.430 1327.000 1500.750 ;
        RECT 1326.800 1469.810 1326.940 1500.430 ;
        RECT 1326.740 1469.490 1327.000 1469.810 ;
        RECT 1327.660 1469.490 1327.920 1469.810 ;
        RECT 1327.720 1380.245 1327.860 1469.490 ;
        RECT 1326.270 1379.875 1326.550 1380.245 ;
        RECT 1327.650 1379.875 1327.930 1380.245 ;
        RECT 1326.340 1345.710 1326.480 1379.875 ;
        RECT 1326.280 1345.390 1326.540 1345.710 ;
        RECT 1325.820 1345.050 1326.080 1345.370 ;
        RECT 1325.880 1331.965 1326.020 1345.050 ;
        RECT 1325.810 1331.595 1326.090 1331.965 ;
        RECT 1326.730 1331.595 1327.010 1331.965 ;
        RECT 1326.800 1297.170 1326.940 1331.595 ;
        RECT 1326.340 1297.030 1326.940 1297.170 ;
        RECT 1326.340 1242.090 1326.480 1297.030 ;
        RECT 1325.880 1241.950 1326.480 1242.090 ;
        RECT 1325.880 1172.050 1326.020 1241.950 ;
        RECT 1325.880 1171.910 1326.480 1172.050 ;
        RECT 1326.340 1136.010 1326.480 1171.910 ;
        RECT 1326.340 1135.870 1326.940 1136.010 ;
        RECT 1326.800 1111.110 1326.940 1135.870 ;
        RECT 1325.820 1110.965 1326.080 1111.110 ;
        RECT 1326.740 1110.965 1327.000 1111.110 ;
        RECT 1325.810 1110.595 1326.090 1110.965 ;
        RECT 1326.730 1110.595 1327.010 1110.965 ;
        RECT 1326.800 1062.740 1326.940 1110.595 ;
        RECT 1326.340 1062.600 1326.940 1062.740 ;
        RECT 1326.340 1062.570 1326.480 1062.600 ;
        RECT 1325.880 1062.430 1326.480 1062.570 ;
        RECT 1325.880 1014.405 1326.020 1062.430 ;
        RECT 1325.810 1014.035 1326.090 1014.405 ;
        RECT 1326.730 1014.035 1327.010 1014.405 ;
        RECT 1326.800 966.270 1326.940 1014.035 ;
        RECT 1326.280 966.125 1326.540 966.270 ;
        RECT 1324.890 965.755 1325.170 966.125 ;
        RECT 1326.270 965.755 1326.550 966.125 ;
        RECT 1326.740 965.950 1327.000 966.270 ;
        RECT 1324.960 917.990 1325.100 965.755 ;
        RECT 1324.900 917.670 1325.160 917.990 ;
        RECT 1325.820 917.845 1326.080 917.990 ;
        RECT 1325.810 917.475 1326.090 917.845 ;
        RECT 1326.730 917.475 1327.010 917.845 ;
        RECT 1326.800 869.710 1326.940 917.475 ;
        RECT 1326.280 869.390 1326.540 869.710 ;
        RECT 1326.740 869.390 1327.000 869.710 ;
        RECT 1326.340 807.490 1326.480 869.390 ;
        RECT 1325.820 807.170 1326.080 807.490 ;
        RECT 1326.280 807.170 1326.540 807.490 ;
        RECT 1325.880 800.350 1326.020 807.170 ;
        RECT 1325.820 800.030 1326.080 800.350 ;
        RECT 1326.740 752.090 1327.000 752.410 ;
        RECT 1326.800 688.570 1326.940 752.090 ;
        RECT 1326.340 688.430 1326.940 688.570 ;
        RECT 1326.340 628.845 1326.480 688.430 ;
        RECT 1326.270 628.475 1326.550 628.845 ;
        RECT 1326.270 627.795 1326.550 628.165 ;
        RECT 1326.340 572.890 1326.480 627.795 ;
        RECT 1325.820 572.570 1326.080 572.890 ;
        RECT 1326.280 572.570 1326.540 572.890 ;
        RECT 1325.880 545.350 1326.020 572.570 ;
        RECT 1325.820 545.030 1326.080 545.350 ;
        RECT 1326.280 544.690 1326.540 545.010 ;
        RECT 1326.340 476.670 1326.480 544.690 ;
        RECT 1326.280 476.350 1326.540 476.670 ;
        RECT 1326.280 462.410 1326.540 462.730 ;
        RECT 1326.340 338.290 1326.480 462.410 ;
        RECT 1325.820 337.970 1326.080 338.290 ;
        RECT 1326.280 337.970 1326.540 338.290 ;
        RECT 1325.880 331.150 1326.020 337.970 ;
        RECT 1325.820 330.830 1326.080 331.150 ;
        RECT 1325.820 254.330 1326.080 254.650 ;
        RECT 1325.880 234.590 1326.020 254.330 ;
        RECT 1325.820 234.270 1326.080 234.590 ;
        RECT 1325.820 186.330 1326.080 186.650 ;
        RECT 1325.880 145.170 1326.020 186.330 ;
        RECT 1325.820 144.850 1326.080 145.170 ;
        RECT 1326.280 144.850 1326.540 145.170 ;
        RECT 1326.340 138.030 1326.480 144.850 ;
        RECT 1326.280 137.710 1326.540 138.030 ;
        RECT 1324.900 89.430 1325.160 89.750 ;
        RECT 1324.960 42.005 1325.100 89.430 ;
        RECT 1324.890 41.635 1325.170 42.005 ;
        RECT 1325.810 41.635 1326.090 42.005 ;
        RECT 1325.880 41.470 1326.020 41.635 ;
        RECT 436.640 41.150 436.900 41.470 ;
        RECT 1325.820 41.150 1326.080 41.470 ;
        RECT 436.700 2.400 436.840 41.150 ;
        RECT 436.490 -4.800 437.050 2.400 ;
      LAYER via2 ;
        RECT 1326.270 1379.920 1326.550 1380.200 ;
        RECT 1327.650 1379.920 1327.930 1380.200 ;
        RECT 1325.810 1331.640 1326.090 1331.920 ;
        RECT 1326.730 1331.640 1327.010 1331.920 ;
        RECT 1325.810 1110.640 1326.090 1110.920 ;
        RECT 1326.730 1110.640 1327.010 1110.920 ;
        RECT 1325.810 1014.080 1326.090 1014.360 ;
        RECT 1326.730 1014.080 1327.010 1014.360 ;
        RECT 1324.890 965.800 1325.170 966.080 ;
        RECT 1326.270 965.800 1326.550 966.080 ;
        RECT 1325.810 917.520 1326.090 917.800 ;
        RECT 1326.730 917.520 1327.010 917.800 ;
        RECT 1326.270 628.520 1326.550 628.800 ;
        RECT 1326.270 627.840 1326.550 628.120 ;
        RECT 1324.890 41.680 1325.170 41.960 ;
        RECT 1325.810 41.680 1326.090 41.960 ;
      LAYER met3 ;
        RECT 1326.245 1380.210 1326.575 1380.225 ;
        RECT 1327.625 1380.210 1327.955 1380.225 ;
        RECT 1326.245 1379.910 1327.955 1380.210 ;
        RECT 1326.245 1379.895 1326.575 1379.910 ;
        RECT 1327.625 1379.895 1327.955 1379.910 ;
        RECT 1325.785 1331.930 1326.115 1331.945 ;
        RECT 1326.705 1331.930 1327.035 1331.945 ;
        RECT 1325.785 1331.630 1327.035 1331.930 ;
        RECT 1325.785 1331.615 1326.115 1331.630 ;
        RECT 1326.705 1331.615 1327.035 1331.630 ;
        RECT 1325.785 1110.930 1326.115 1110.945 ;
        RECT 1326.705 1110.930 1327.035 1110.945 ;
        RECT 1325.785 1110.630 1327.035 1110.930 ;
        RECT 1325.785 1110.615 1326.115 1110.630 ;
        RECT 1326.705 1110.615 1327.035 1110.630 ;
        RECT 1325.785 1014.370 1326.115 1014.385 ;
        RECT 1326.705 1014.370 1327.035 1014.385 ;
        RECT 1325.785 1014.070 1327.035 1014.370 ;
        RECT 1325.785 1014.055 1326.115 1014.070 ;
        RECT 1326.705 1014.055 1327.035 1014.070 ;
        RECT 1324.865 966.090 1325.195 966.105 ;
        RECT 1326.245 966.090 1326.575 966.105 ;
        RECT 1324.865 965.790 1326.575 966.090 ;
        RECT 1324.865 965.775 1325.195 965.790 ;
        RECT 1326.245 965.775 1326.575 965.790 ;
        RECT 1325.785 917.810 1326.115 917.825 ;
        RECT 1326.705 917.810 1327.035 917.825 ;
        RECT 1325.785 917.510 1327.035 917.810 ;
        RECT 1325.785 917.495 1326.115 917.510 ;
        RECT 1326.705 917.495 1327.035 917.510 ;
        RECT 1326.245 628.810 1326.575 628.825 ;
        RECT 1326.030 628.495 1326.575 628.810 ;
        RECT 1326.030 628.145 1326.330 628.495 ;
        RECT 1326.030 627.830 1326.575 628.145 ;
        RECT 1326.245 627.815 1326.575 627.830 ;
        RECT 1324.865 41.970 1325.195 41.985 ;
        RECT 1325.785 41.970 1326.115 41.985 ;
        RECT 1324.865 41.670 1326.115 41.970 ;
        RECT 1324.865 41.655 1325.195 41.670 ;
        RECT 1325.785 41.655 1326.115 41.670 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1333.225 1594.005 1333.395 1608.115 ;
        RECT 1333.225 1524.985 1333.395 1546.235 ;
        RECT 1333.685 1442.025 1333.855 1490.475 ;
        RECT 1333.685 1297.185 1333.855 1318.095 ;
        RECT 1333.225 807.245 1333.395 855.355 ;
        RECT 1333.685 186.405 1333.855 234.515 ;
      LAYER mcon ;
        RECT 1333.225 1607.945 1333.395 1608.115 ;
        RECT 1333.225 1546.065 1333.395 1546.235 ;
        RECT 1333.685 1490.305 1333.855 1490.475 ;
        RECT 1333.685 1317.925 1333.855 1318.095 ;
        RECT 1333.225 855.185 1333.395 855.355 ;
        RECT 1333.685 234.345 1333.855 234.515 ;
      LAYER met1 ;
        RECT 1333.165 1608.100 1333.455 1608.145 ;
        RECT 1333.610 1608.100 1333.930 1608.160 ;
        RECT 1333.165 1607.960 1333.930 1608.100 ;
        RECT 1333.165 1607.915 1333.455 1607.960 ;
        RECT 1333.610 1607.900 1333.930 1607.960 ;
        RECT 1333.150 1594.160 1333.470 1594.220 ;
        RECT 1332.955 1594.020 1333.470 1594.160 ;
        RECT 1333.150 1593.960 1333.470 1594.020 ;
        RECT 1333.150 1546.220 1333.470 1546.280 ;
        RECT 1332.955 1546.080 1333.470 1546.220 ;
        RECT 1333.150 1546.020 1333.470 1546.080 ;
        RECT 1333.150 1525.140 1333.470 1525.200 ;
        RECT 1332.955 1525.000 1333.470 1525.140 ;
        RECT 1333.150 1524.940 1333.470 1525.000 ;
        RECT 1333.150 1497.600 1333.470 1497.660 ;
        RECT 1333.610 1497.600 1333.930 1497.660 ;
        RECT 1333.150 1497.460 1333.930 1497.600 ;
        RECT 1333.150 1497.400 1333.470 1497.460 ;
        RECT 1333.610 1497.400 1333.930 1497.460 ;
        RECT 1333.610 1490.460 1333.930 1490.520 ;
        RECT 1333.415 1490.320 1333.930 1490.460 ;
        RECT 1333.610 1490.260 1333.930 1490.320 ;
        RECT 1333.625 1442.180 1333.915 1442.225 ;
        RECT 1334.070 1442.180 1334.390 1442.240 ;
        RECT 1333.625 1442.040 1334.390 1442.180 ;
        RECT 1333.625 1441.995 1333.915 1442.040 ;
        RECT 1334.070 1441.980 1334.390 1442.040 ;
        RECT 1333.610 1401.040 1333.930 1401.100 ;
        RECT 1334.070 1401.040 1334.390 1401.100 ;
        RECT 1333.610 1400.900 1334.390 1401.040 ;
        RECT 1333.610 1400.840 1333.930 1400.900 ;
        RECT 1334.070 1400.840 1334.390 1400.900 ;
        RECT 1333.610 1318.080 1333.930 1318.140 ;
        RECT 1333.415 1317.940 1333.930 1318.080 ;
        RECT 1333.610 1317.880 1333.930 1317.940 ;
        RECT 1333.610 1297.340 1333.930 1297.400 ;
        RECT 1333.415 1297.200 1333.930 1297.340 ;
        RECT 1333.610 1297.140 1333.930 1297.200 ;
        RECT 1333.150 1207.580 1333.470 1207.640 ;
        RECT 1333.610 1207.580 1333.930 1207.640 ;
        RECT 1333.150 1207.440 1333.930 1207.580 ;
        RECT 1333.150 1207.380 1333.470 1207.440 ;
        RECT 1333.610 1207.380 1333.930 1207.440 ;
        RECT 1333.610 990.460 1333.930 990.720 ;
        RECT 1333.700 990.040 1333.840 990.460 ;
        RECT 1333.610 989.780 1333.930 990.040 ;
        RECT 1333.150 931.640 1333.470 931.900 ;
        RECT 1333.240 931.160 1333.380 931.640 ;
        RECT 1333.610 931.160 1333.930 931.220 ;
        RECT 1333.240 931.020 1333.930 931.160 ;
        RECT 1333.610 930.960 1333.930 931.020 ;
        RECT 1333.610 893.900 1333.930 894.160 ;
        RECT 1333.700 893.480 1333.840 893.900 ;
        RECT 1333.610 893.220 1333.930 893.480 ;
        RECT 1333.150 855.340 1333.470 855.400 ;
        RECT 1332.955 855.200 1333.470 855.340 ;
        RECT 1333.150 855.140 1333.470 855.200 ;
        RECT 1333.165 807.400 1333.455 807.445 ;
        RECT 1334.070 807.400 1334.390 807.460 ;
        RECT 1333.165 807.260 1334.390 807.400 ;
        RECT 1333.165 807.215 1333.455 807.260 ;
        RECT 1334.070 807.200 1334.390 807.260 ;
        RECT 1334.070 758.920 1334.390 759.180 ;
        RECT 1334.160 758.500 1334.300 758.920 ;
        RECT 1334.070 758.240 1334.390 758.500 ;
        RECT 1333.150 386.480 1333.470 386.540 ;
        RECT 1333.610 386.480 1333.930 386.540 ;
        RECT 1333.150 386.340 1333.930 386.480 ;
        RECT 1333.150 386.280 1333.470 386.340 ;
        RECT 1333.610 386.280 1333.930 386.340 ;
        RECT 1333.150 303.660 1333.470 303.920 ;
        RECT 1333.240 303.180 1333.380 303.660 ;
        RECT 1333.610 303.180 1333.930 303.240 ;
        RECT 1333.240 303.040 1333.930 303.180 ;
        RECT 1333.610 302.980 1333.930 303.040 ;
        RECT 1333.610 234.500 1333.930 234.560 ;
        RECT 1333.415 234.360 1333.930 234.500 ;
        RECT 1333.610 234.300 1333.930 234.360 ;
        RECT 1333.610 186.560 1333.930 186.620 ;
        RECT 1333.415 186.420 1333.930 186.560 ;
        RECT 1333.610 186.360 1333.930 186.420 ;
        RECT 1333.610 97.140 1333.930 97.200 ;
        RECT 1333.240 97.000 1333.930 97.140 ;
        RECT 1333.240 96.520 1333.380 97.000 ;
        RECT 1333.610 96.940 1333.930 97.000 ;
        RECT 1333.150 96.260 1333.470 96.520 ;
        RECT 455.010 52.940 455.330 53.000 ;
        RECT 1333.150 52.940 1333.470 53.000 ;
        RECT 455.010 52.800 1333.470 52.940 ;
        RECT 455.010 52.740 455.330 52.800 ;
        RECT 1333.150 52.740 1333.470 52.800 ;
      LAYER via ;
        RECT 1333.640 1607.900 1333.900 1608.160 ;
        RECT 1333.180 1593.960 1333.440 1594.220 ;
        RECT 1333.180 1546.020 1333.440 1546.280 ;
        RECT 1333.180 1524.940 1333.440 1525.200 ;
        RECT 1333.180 1497.400 1333.440 1497.660 ;
        RECT 1333.640 1497.400 1333.900 1497.660 ;
        RECT 1333.640 1490.260 1333.900 1490.520 ;
        RECT 1334.100 1441.980 1334.360 1442.240 ;
        RECT 1333.640 1400.840 1333.900 1401.100 ;
        RECT 1334.100 1400.840 1334.360 1401.100 ;
        RECT 1333.640 1317.880 1333.900 1318.140 ;
        RECT 1333.640 1297.140 1333.900 1297.400 ;
        RECT 1333.180 1207.380 1333.440 1207.640 ;
        RECT 1333.640 1207.380 1333.900 1207.640 ;
        RECT 1333.640 990.460 1333.900 990.720 ;
        RECT 1333.640 989.780 1333.900 990.040 ;
        RECT 1333.180 931.640 1333.440 931.900 ;
        RECT 1333.640 930.960 1333.900 931.220 ;
        RECT 1333.640 893.900 1333.900 894.160 ;
        RECT 1333.640 893.220 1333.900 893.480 ;
        RECT 1333.180 855.140 1333.440 855.400 ;
        RECT 1334.100 807.200 1334.360 807.460 ;
        RECT 1334.100 758.920 1334.360 759.180 ;
        RECT 1334.100 758.240 1334.360 758.500 ;
        RECT 1333.180 386.280 1333.440 386.540 ;
        RECT 1333.640 386.280 1333.900 386.540 ;
        RECT 1333.180 303.660 1333.440 303.920 ;
        RECT 1333.640 302.980 1333.900 303.240 ;
        RECT 1333.640 234.300 1333.900 234.560 ;
        RECT 1333.640 186.360 1333.900 186.620 ;
        RECT 1333.640 96.940 1333.900 97.200 ;
        RECT 1333.180 96.260 1333.440 96.520 ;
        RECT 455.040 52.740 455.300 53.000 ;
        RECT 1333.180 52.740 1333.440 53.000 ;
      LAYER met2 ;
        RECT 1335.865 1700.410 1336.145 1704.000 ;
        RECT 1334.620 1700.270 1336.145 1700.410 ;
        RECT 1334.620 1677.970 1334.760 1700.270 ;
        RECT 1335.865 1700.000 1336.145 1700.270 ;
        RECT 1333.700 1677.830 1334.760 1677.970 ;
        RECT 1333.700 1608.190 1333.840 1677.830 ;
        RECT 1333.640 1607.870 1333.900 1608.190 ;
        RECT 1333.180 1593.930 1333.440 1594.250 ;
        RECT 1333.240 1546.310 1333.380 1593.930 ;
        RECT 1333.180 1545.990 1333.440 1546.310 ;
        RECT 1333.180 1524.910 1333.440 1525.230 ;
        RECT 1333.240 1497.690 1333.380 1524.910 ;
        RECT 1333.180 1497.370 1333.440 1497.690 ;
        RECT 1333.640 1497.370 1333.900 1497.690 ;
        RECT 1333.700 1490.550 1333.840 1497.370 ;
        RECT 1333.640 1490.230 1333.900 1490.550 ;
        RECT 1334.100 1441.950 1334.360 1442.270 ;
        RECT 1334.160 1401.130 1334.300 1441.950 ;
        RECT 1333.640 1400.810 1333.900 1401.130 ;
        RECT 1334.100 1400.810 1334.360 1401.130 ;
        RECT 1333.700 1318.170 1333.840 1400.810 ;
        RECT 1333.640 1317.850 1333.900 1318.170 ;
        RECT 1333.700 1297.430 1333.840 1297.585 ;
        RECT 1333.640 1297.170 1333.900 1297.430 ;
        RECT 1333.240 1297.110 1333.900 1297.170 ;
        RECT 1333.240 1297.030 1333.840 1297.110 ;
        RECT 1333.240 1207.670 1333.380 1297.030 ;
        RECT 1333.180 1207.350 1333.440 1207.670 ;
        RECT 1333.640 1207.350 1333.900 1207.670 ;
        RECT 1333.700 1176.810 1333.840 1207.350 ;
        RECT 1333.700 1176.670 1334.300 1176.810 ;
        RECT 1334.160 1104.165 1334.300 1176.670 ;
        RECT 1333.170 1103.795 1333.450 1104.165 ;
        RECT 1334.090 1103.795 1334.370 1104.165 ;
        RECT 1333.240 1079.570 1333.380 1103.795 ;
        RECT 1333.240 1079.430 1333.840 1079.570 ;
        RECT 1333.700 990.750 1333.840 1079.430 ;
        RECT 1333.640 990.430 1333.900 990.750 ;
        RECT 1333.640 989.750 1333.900 990.070 ;
        RECT 1333.700 966.180 1333.840 989.750 ;
        RECT 1333.240 966.040 1333.840 966.180 ;
        RECT 1333.240 931.930 1333.380 966.040 ;
        RECT 1333.180 931.610 1333.440 931.930 ;
        RECT 1333.640 930.930 1333.900 931.250 ;
        RECT 1333.700 894.190 1333.840 930.930 ;
        RECT 1333.640 893.870 1333.900 894.190 ;
        RECT 1333.640 893.190 1333.900 893.510 ;
        RECT 1333.700 869.620 1333.840 893.190 ;
        RECT 1333.240 869.480 1333.840 869.620 ;
        RECT 1333.240 855.430 1333.380 869.480 ;
        RECT 1333.180 855.110 1333.440 855.430 ;
        RECT 1334.100 807.170 1334.360 807.490 ;
        RECT 1334.160 759.210 1334.300 807.170 ;
        RECT 1334.100 758.890 1334.360 759.210 ;
        RECT 1334.100 758.210 1334.360 758.530 ;
        RECT 1334.160 699.450 1334.300 758.210 ;
        RECT 1333.700 699.310 1334.300 699.450 ;
        RECT 1333.700 628.845 1333.840 699.310 ;
        RECT 1333.630 628.475 1333.910 628.845 ;
        RECT 1333.170 627.795 1333.450 628.165 ;
        RECT 1333.240 386.570 1333.380 627.795 ;
        RECT 1333.180 386.250 1333.440 386.570 ;
        RECT 1333.640 386.250 1333.900 386.570 ;
        RECT 1333.700 338.370 1333.840 386.250 ;
        RECT 1333.240 338.230 1333.840 338.370 ;
        RECT 1333.240 303.950 1333.380 338.230 ;
        RECT 1333.180 303.630 1333.440 303.950 ;
        RECT 1333.640 302.950 1333.900 303.270 ;
        RECT 1333.700 234.590 1333.840 302.950 ;
        RECT 1333.640 234.270 1333.900 234.590 ;
        RECT 1333.640 186.330 1333.900 186.650 ;
        RECT 1333.700 97.230 1333.840 186.330 ;
        RECT 1333.640 96.910 1333.900 97.230 ;
        RECT 1333.180 96.230 1333.440 96.550 ;
        RECT 1333.240 53.030 1333.380 96.230 ;
        RECT 455.040 52.710 455.300 53.030 ;
        RECT 1333.180 52.710 1333.440 53.030 ;
        RECT 455.100 17.410 455.240 52.710 ;
        RECT 454.640 17.270 455.240 17.410 ;
        RECT 454.640 2.400 454.780 17.270 ;
        RECT 454.430 -4.800 454.990 2.400 ;
      LAYER via2 ;
        RECT 1333.170 1103.840 1333.450 1104.120 ;
        RECT 1334.090 1103.840 1334.370 1104.120 ;
        RECT 1333.630 628.520 1333.910 628.800 ;
        RECT 1333.170 627.840 1333.450 628.120 ;
      LAYER met3 ;
        RECT 1333.145 1104.130 1333.475 1104.145 ;
        RECT 1334.065 1104.130 1334.395 1104.145 ;
        RECT 1333.145 1103.830 1334.395 1104.130 ;
        RECT 1333.145 1103.815 1333.475 1103.830 ;
        RECT 1334.065 1103.815 1334.395 1103.830 ;
        RECT 1333.605 628.810 1333.935 628.825 ;
        RECT 1333.390 628.495 1333.935 628.810 ;
        RECT 1333.390 628.145 1333.690 628.495 ;
        RECT 1333.145 627.830 1333.690 628.145 ;
        RECT 1333.145 627.815 1333.475 627.830 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1338.745 1594.005 1338.915 1608.115 ;
        RECT 1338.745 1555.585 1338.915 1579.895 ;
        RECT 1339.205 1435.225 1339.375 1482.995 ;
        RECT 1339.205 848.725 1339.375 896.835 ;
        RECT 1339.205 365.925 1339.375 414.035 ;
        RECT 1338.745 53.125 1338.915 113.135 ;
      LAYER mcon ;
        RECT 1338.745 1607.945 1338.915 1608.115 ;
        RECT 1338.745 1579.725 1338.915 1579.895 ;
        RECT 1339.205 1482.825 1339.375 1482.995 ;
        RECT 1339.205 896.665 1339.375 896.835 ;
        RECT 1339.205 413.865 1339.375 414.035 ;
        RECT 1338.745 112.965 1338.915 113.135 ;
      LAYER met1 ;
        RECT 1338.685 1608.100 1338.975 1608.145 ;
        RECT 1339.130 1608.100 1339.450 1608.160 ;
        RECT 1338.685 1607.960 1339.450 1608.100 ;
        RECT 1338.685 1607.915 1338.975 1607.960 ;
        RECT 1339.130 1607.900 1339.450 1607.960 ;
        RECT 1338.670 1594.160 1338.990 1594.220 ;
        RECT 1338.475 1594.020 1338.990 1594.160 ;
        RECT 1338.670 1593.960 1338.990 1594.020 ;
        RECT 1338.670 1579.880 1338.990 1579.940 ;
        RECT 1338.670 1579.740 1339.185 1579.880 ;
        RECT 1338.670 1579.680 1338.990 1579.740 ;
        RECT 1338.685 1555.740 1338.975 1555.785 ;
        RECT 1339.130 1555.740 1339.450 1555.800 ;
        RECT 1338.685 1555.600 1339.450 1555.740 ;
        RECT 1338.685 1555.555 1338.975 1555.600 ;
        RECT 1339.130 1555.540 1339.450 1555.600 ;
        RECT 1338.670 1483.660 1338.990 1483.720 ;
        RECT 1340.050 1483.660 1340.370 1483.720 ;
        RECT 1338.670 1483.520 1340.370 1483.660 ;
        RECT 1338.670 1483.460 1338.990 1483.520 ;
        RECT 1340.050 1483.460 1340.370 1483.520 ;
        RECT 1338.670 1482.980 1338.990 1483.040 ;
        RECT 1339.145 1482.980 1339.435 1483.025 ;
        RECT 1338.670 1482.840 1339.435 1482.980 ;
        RECT 1338.670 1482.780 1338.990 1482.840 ;
        RECT 1339.145 1482.795 1339.435 1482.840 ;
        RECT 1338.670 1435.380 1338.990 1435.440 ;
        RECT 1339.145 1435.380 1339.435 1435.425 ;
        RECT 1338.670 1435.240 1339.435 1435.380 ;
        RECT 1338.670 1435.180 1338.990 1435.240 ;
        RECT 1339.145 1435.195 1339.435 1435.240 ;
        RECT 1338.670 1200.780 1338.990 1200.840 ;
        RECT 1339.130 1200.780 1339.450 1200.840 ;
        RECT 1338.670 1200.640 1339.450 1200.780 ;
        RECT 1338.670 1200.580 1338.990 1200.640 ;
        RECT 1339.130 1200.580 1339.450 1200.640 ;
        RECT 1338.670 1173.380 1338.990 1173.640 ;
        RECT 1338.760 1172.960 1338.900 1173.380 ;
        RECT 1338.670 1172.700 1338.990 1172.960 ;
        RECT 1339.130 966.180 1339.450 966.240 ;
        RECT 1339.590 966.180 1339.910 966.240 ;
        RECT 1339.130 966.040 1339.910 966.180 ;
        RECT 1339.130 965.980 1339.450 966.040 ;
        RECT 1339.590 965.980 1339.910 966.040 ;
        RECT 1338.670 952.240 1338.990 952.300 ;
        RECT 1339.130 952.240 1339.450 952.300 ;
        RECT 1338.670 952.100 1339.450 952.240 ;
        RECT 1338.670 952.040 1338.990 952.100 ;
        RECT 1339.130 952.040 1339.450 952.100 ;
        RECT 1339.130 903.960 1339.450 904.020 ;
        RECT 1339.590 903.960 1339.910 904.020 ;
        RECT 1339.130 903.820 1339.910 903.960 ;
        RECT 1339.130 903.760 1339.450 903.820 ;
        RECT 1339.590 903.760 1339.910 903.820 ;
        RECT 1339.130 896.820 1339.450 896.880 ;
        RECT 1338.935 896.680 1339.450 896.820 ;
        RECT 1339.130 896.620 1339.450 896.680 ;
        RECT 1339.130 848.880 1339.450 848.940 ;
        RECT 1338.935 848.740 1339.450 848.880 ;
        RECT 1339.130 848.680 1339.450 848.740 ;
        RECT 1338.670 787.140 1338.990 787.400 ;
        RECT 1338.760 786.720 1338.900 787.140 ;
        RECT 1338.670 786.460 1338.990 786.720 ;
        RECT 1338.670 724.440 1338.990 724.500 ;
        RECT 1339.590 724.440 1339.910 724.500 ;
        RECT 1338.670 724.300 1339.910 724.440 ;
        RECT 1338.670 724.240 1338.990 724.300 ;
        RECT 1339.590 724.240 1339.910 724.300 ;
        RECT 1338.670 524.520 1338.990 524.580 ;
        RECT 1339.130 524.520 1339.450 524.580 ;
        RECT 1338.670 524.380 1339.450 524.520 ;
        RECT 1338.670 524.320 1338.990 524.380 ;
        RECT 1339.130 524.320 1339.450 524.380 ;
        RECT 1339.130 497.320 1339.450 497.380 ;
        RECT 1338.760 497.180 1339.450 497.320 ;
        RECT 1338.760 496.700 1338.900 497.180 ;
        RECT 1339.130 497.120 1339.450 497.180 ;
        RECT 1338.670 496.440 1338.990 496.700 ;
        RECT 1338.670 427.760 1338.990 428.020 ;
        RECT 1338.760 427.280 1338.900 427.760 ;
        RECT 1339.130 427.280 1339.450 427.340 ;
        RECT 1338.760 427.140 1339.450 427.280 ;
        RECT 1339.130 427.080 1339.450 427.140 ;
        RECT 1339.130 414.020 1339.450 414.080 ;
        RECT 1338.935 413.880 1339.450 414.020 ;
        RECT 1339.130 413.820 1339.450 413.880 ;
        RECT 1339.145 366.080 1339.435 366.125 ;
        RECT 1339.590 366.080 1339.910 366.140 ;
        RECT 1339.145 365.940 1339.910 366.080 ;
        RECT 1339.145 365.895 1339.435 365.940 ;
        RECT 1339.590 365.880 1339.910 365.940 ;
        RECT 1339.590 324.940 1339.910 325.000 ;
        RECT 1338.760 324.800 1339.910 324.940 ;
        RECT 1338.760 324.660 1338.900 324.800 ;
        RECT 1339.590 324.740 1339.910 324.800 ;
        RECT 1338.670 324.400 1338.990 324.660 ;
        RECT 1338.670 304.000 1338.990 304.260 ;
        RECT 1338.760 303.580 1338.900 304.000 ;
        RECT 1338.670 303.320 1338.990 303.580 ;
        RECT 1339.590 193.500 1339.910 193.760 ;
        RECT 1339.680 193.080 1339.820 193.500 ;
        RECT 1339.590 192.820 1339.910 193.080 ;
        RECT 1339.130 145.080 1339.450 145.140 ;
        RECT 1339.590 145.080 1339.910 145.140 ;
        RECT 1339.130 144.940 1339.910 145.080 ;
        RECT 1339.130 144.880 1339.450 144.940 ;
        RECT 1339.590 144.880 1339.910 144.940 ;
        RECT 1338.685 113.120 1338.975 113.165 ;
        RECT 1339.130 113.120 1339.450 113.180 ;
        RECT 1338.685 112.980 1339.450 113.120 ;
        RECT 1338.685 112.935 1338.975 112.980 ;
        RECT 1339.130 112.920 1339.450 112.980 ;
        RECT 475.710 53.280 476.030 53.340 ;
        RECT 1338.685 53.280 1338.975 53.325 ;
        RECT 475.710 53.140 1338.975 53.280 ;
        RECT 475.710 53.080 476.030 53.140 ;
        RECT 1338.685 53.095 1338.975 53.140 ;
        RECT 472.490 15.540 472.810 15.600 ;
        RECT 475.710 15.540 476.030 15.600 ;
        RECT 472.490 15.400 476.030 15.540 ;
        RECT 472.490 15.340 472.810 15.400 ;
        RECT 475.710 15.340 476.030 15.400 ;
      LAYER via ;
        RECT 1339.160 1607.900 1339.420 1608.160 ;
        RECT 1338.700 1593.960 1338.960 1594.220 ;
        RECT 1338.700 1579.680 1338.960 1579.940 ;
        RECT 1339.160 1555.540 1339.420 1555.800 ;
        RECT 1338.700 1483.460 1338.960 1483.720 ;
        RECT 1340.080 1483.460 1340.340 1483.720 ;
        RECT 1338.700 1482.780 1338.960 1483.040 ;
        RECT 1338.700 1435.180 1338.960 1435.440 ;
        RECT 1338.700 1200.580 1338.960 1200.840 ;
        RECT 1339.160 1200.580 1339.420 1200.840 ;
        RECT 1338.700 1173.380 1338.960 1173.640 ;
        RECT 1338.700 1172.700 1338.960 1172.960 ;
        RECT 1339.160 965.980 1339.420 966.240 ;
        RECT 1339.620 965.980 1339.880 966.240 ;
        RECT 1338.700 952.040 1338.960 952.300 ;
        RECT 1339.160 952.040 1339.420 952.300 ;
        RECT 1339.160 903.760 1339.420 904.020 ;
        RECT 1339.620 903.760 1339.880 904.020 ;
        RECT 1339.160 896.620 1339.420 896.880 ;
        RECT 1339.160 848.680 1339.420 848.940 ;
        RECT 1338.700 787.140 1338.960 787.400 ;
        RECT 1338.700 786.460 1338.960 786.720 ;
        RECT 1338.700 724.240 1338.960 724.500 ;
        RECT 1339.620 724.240 1339.880 724.500 ;
        RECT 1338.700 524.320 1338.960 524.580 ;
        RECT 1339.160 524.320 1339.420 524.580 ;
        RECT 1339.160 497.120 1339.420 497.380 ;
        RECT 1338.700 496.440 1338.960 496.700 ;
        RECT 1338.700 427.760 1338.960 428.020 ;
        RECT 1339.160 427.080 1339.420 427.340 ;
        RECT 1339.160 413.820 1339.420 414.080 ;
        RECT 1339.620 365.880 1339.880 366.140 ;
        RECT 1339.620 324.740 1339.880 325.000 ;
        RECT 1338.700 324.400 1338.960 324.660 ;
        RECT 1338.700 304.000 1338.960 304.260 ;
        RECT 1338.700 303.320 1338.960 303.580 ;
        RECT 1339.620 193.500 1339.880 193.760 ;
        RECT 1339.620 192.820 1339.880 193.080 ;
        RECT 1339.160 144.880 1339.420 145.140 ;
        RECT 1339.620 144.880 1339.880 145.140 ;
        RECT 1339.160 112.920 1339.420 113.180 ;
        RECT 475.740 53.080 476.000 53.340 ;
        RECT 472.520 15.340 472.780 15.600 ;
        RECT 475.740 15.340 476.000 15.600 ;
      LAYER met2 ;
        RECT 1343.225 1700.410 1343.505 1704.000 ;
        RECT 1341.980 1700.270 1343.505 1700.410 ;
        RECT 1341.980 1677.970 1342.120 1700.270 ;
        RECT 1343.225 1700.000 1343.505 1700.270 ;
        RECT 1339.220 1677.830 1342.120 1677.970 ;
        RECT 1339.220 1608.190 1339.360 1677.830 ;
        RECT 1339.160 1607.870 1339.420 1608.190 ;
        RECT 1338.700 1593.930 1338.960 1594.250 ;
        RECT 1338.760 1579.970 1338.900 1593.930 ;
        RECT 1338.700 1579.650 1338.960 1579.970 ;
        RECT 1339.160 1555.510 1339.420 1555.830 ;
        RECT 1339.220 1531.885 1339.360 1555.510 ;
        RECT 1339.150 1531.515 1339.430 1531.885 ;
        RECT 1340.070 1531.515 1340.350 1531.885 ;
        RECT 1340.140 1483.750 1340.280 1531.515 ;
        RECT 1338.700 1483.430 1338.960 1483.750 ;
        RECT 1340.080 1483.430 1340.340 1483.750 ;
        RECT 1338.760 1483.070 1338.900 1483.430 ;
        RECT 1338.700 1482.750 1338.960 1483.070 ;
        RECT 1338.700 1435.150 1338.960 1435.470 ;
        RECT 1338.760 1345.565 1338.900 1435.150 ;
        RECT 1338.690 1345.195 1338.970 1345.565 ;
        RECT 1339.150 1344.515 1339.430 1344.885 ;
        RECT 1339.220 1200.870 1339.360 1344.515 ;
        RECT 1338.700 1200.550 1338.960 1200.870 ;
        RECT 1339.160 1200.550 1339.420 1200.870 ;
        RECT 1338.760 1173.670 1338.900 1200.550 ;
        RECT 1338.700 1173.350 1338.960 1173.670 ;
        RECT 1338.700 1172.670 1338.960 1172.990 ;
        RECT 1338.760 1110.965 1338.900 1172.670 ;
        RECT 1338.690 1110.595 1338.970 1110.965 ;
        RECT 1338.690 1109.915 1338.970 1110.285 ;
        RECT 1338.760 1062.740 1338.900 1109.915 ;
        RECT 1338.760 1062.600 1339.360 1062.740 ;
        RECT 1339.220 1014.460 1339.360 1062.600 ;
        RECT 1338.760 1014.405 1339.360 1014.460 ;
        RECT 1338.690 1014.320 1339.360 1014.405 ;
        RECT 1338.690 1014.035 1338.970 1014.320 ;
        RECT 1339.610 1014.035 1339.890 1014.405 ;
        RECT 1339.680 966.270 1339.820 1014.035 ;
        RECT 1339.160 965.950 1339.420 966.270 ;
        RECT 1339.620 965.950 1339.880 966.270 ;
        RECT 1339.220 952.330 1339.360 965.950 ;
        RECT 1338.700 952.010 1338.960 952.330 ;
        RECT 1339.160 952.010 1339.420 952.330 ;
        RECT 1338.760 904.245 1338.900 952.010 ;
        RECT 1338.690 903.875 1338.970 904.245 ;
        RECT 1339.160 903.730 1339.420 904.050 ;
        RECT 1339.610 903.875 1339.890 904.245 ;
        RECT 1339.620 903.730 1339.880 903.875 ;
        RECT 1339.220 896.910 1339.360 903.730 ;
        RECT 1339.160 896.590 1339.420 896.910 ;
        RECT 1339.160 848.650 1339.420 848.970 ;
        RECT 1339.220 807.570 1339.360 848.650 ;
        RECT 1338.760 807.430 1339.360 807.570 ;
        RECT 1338.760 787.430 1338.900 807.430 ;
        RECT 1338.700 787.110 1338.960 787.430 ;
        RECT 1338.700 786.430 1338.960 786.750 ;
        RECT 1338.760 724.530 1338.900 786.430 ;
        RECT 1338.700 724.210 1338.960 724.530 ;
        RECT 1339.620 724.210 1339.880 724.530 ;
        RECT 1339.680 699.450 1339.820 724.210 ;
        RECT 1339.220 699.310 1339.820 699.450 ;
        RECT 1339.220 628.845 1339.360 699.310 ;
        RECT 1339.150 628.475 1339.430 628.845 ;
        RECT 1338.690 627.795 1338.970 628.165 ;
        RECT 1338.760 524.610 1338.900 627.795 ;
        RECT 1338.700 524.290 1338.960 524.610 ;
        RECT 1339.160 524.290 1339.420 524.610 ;
        RECT 1339.220 497.410 1339.360 524.290 ;
        RECT 1339.160 497.090 1339.420 497.410 ;
        RECT 1338.700 496.410 1338.960 496.730 ;
        RECT 1338.760 428.050 1338.900 496.410 ;
        RECT 1338.700 427.730 1338.960 428.050 ;
        RECT 1339.160 427.050 1339.420 427.370 ;
        RECT 1339.220 414.110 1339.360 427.050 ;
        RECT 1339.160 413.790 1339.420 414.110 ;
        RECT 1339.620 365.850 1339.880 366.170 ;
        RECT 1339.680 325.030 1339.820 365.850 ;
        RECT 1339.620 324.710 1339.880 325.030 ;
        RECT 1338.700 324.370 1338.960 324.690 ;
        RECT 1338.760 304.290 1338.900 324.370 ;
        RECT 1338.700 303.970 1338.960 304.290 ;
        RECT 1338.700 303.290 1338.960 303.610 ;
        RECT 1338.760 241.925 1338.900 303.290 ;
        RECT 1338.690 241.555 1338.970 241.925 ;
        RECT 1339.610 240.875 1339.890 241.245 ;
        RECT 1339.680 193.790 1339.820 240.875 ;
        RECT 1339.620 193.470 1339.880 193.790 ;
        RECT 1339.620 192.790 1339.880 193.110 ;
        RECT 1339.680 145.170 1339.820 192.790 ;
        RECT 1339.160 144.850 1339.420 145.170 ;
        RECT 1339.620 144.850 1339.880 145.170 ;
        RECT 1339.220 113.210 1339.360 144.850 ;
        RECT 1339.160 112.890 1339.420 113.210 ;
        RECT 475.740 53.050 476.000 53.370 ;
        RECT 475.800 15.630 475.940 53.050 ;
        RECT 472.520 15.310 472.780 15.630 ;
        RECT 475.740 15.310 476.000 15.630 ;
        RECT 472.580 2.400 472.720 15.310 ;
        RECT 472.370 -4.800 472.930 2.400 ;
      LAYER via2 ;
        RECT 1339.150 1531.560 1339.430 1531.840 ;
        RECT 1340.070 1531.560 1340.350 1531.840 ;
        RECT 1338.690 1345.240 1338.970 1345.520 ;
        RECT 1339.150 1344.560 1339.430 1344.840 ;
        RECT 1338.690 1110.640 1338.970 1110.920 ;
        RECT 1338.690 1109.960 1338.970 1110.240 ;
        RECT 1338.690 1014.080 1338.970 1014.360 ;
        RECT 1339.610 1014.080 1339.890 1014.360 ;
        RECT 1338.690 903.920 1338.970 904.200 ;
        RECT 1339.610 903.920 1339.890 904.200 ;
        RECT 1339.150 628.520 1339.430 628.800 ;
        RECT 1338.690 627.840 1338.970 628.120 ;
        RECT 1338.690 241.600 1338.970 241.880 ;
        RECT 1339.610 240.920 1339.890 241.200 ;
      LAYER met3 ;
        RECT 1339.125 1531.850 1339.455 1531.865 ;
        RECT 1340.045 1531.850 1340.375 1531.865 ;
        RECT 1339.125 1531.550 1340.375 1531.850 ;
        RECT 1339.125 1531.535 1339.455 1531.550 ;
        RECT 1340.045 1531.535 1340.375 1531.550 ;
        RECT 1338.665 1345.530 1338.995 1345.545 ;
        RECT 1338.665 1345.215 1339.210 1345.530 ;
        RECT 1338.910 1344.865 1339.210 1345.215 ;
        RECT 1338.910 1344.550 1339.455 1344.865 ;
        RECT 1339.125 1344.535 1339.455 1344.550 ;
        RECT 1338.665 1110.930 1338.995 1110.945 ;
        RECT 1338.665 1110.615 1339.210 1110.930 ;
        RECT 1338.910 1110.265 1339.210 1110.615 ;
        RECT 1338.665 1109.950 1339.210 1110.265 ;
        RECT 1338.665 1109.935 1338.995 1109.950 ;
        RECT 1338.665 1014.370 1338.995 1014.385 ;
        RECT 1339.585 1014.370 1339.915 1014.385 ;
        RECT 1338.665 1014.070 1339.915 1014.370 ;
        RECT 1338.665 1014.055 1338.995 1014.070 ;
        RECT 1339.585 1014.055 1339.915 1014.070 ;
        RECT 1338.665 904.210 1338.995 904.225 ;
        RECT 1339.585 904.210 1339.915 904.225 ;
        RECT 1338.665 903.910 1339.915 904.210 ;
        RECT 1338.665 903.895 1338.995 903.910 ;
        RECT 1339.585 903.895 1339.915 903.910 ;
        RECT 1339.125 628.810 1339.455 628.825 ;
        RECT 1338.910 628.495 1339.455 628.810 ;
        RECT 1338.910 628.145 1339.210 628.495 ;
        RECT 1338.665 627.830 1339.210 628.145 ;
        RECT 1338.665 627.815 1338.995 627.830 ;
        RECT 1338.665 241.890 1338.995 241.905 ;
        RECT 1338.665 241.575 1339.210 241.890 ;
        RECT 1338.910 241.210 1339.210 241.575 ;
        RECT 1339.585 241.210 1339.915 241.225 ;
        RECT 1338.910 240.910 1339.915 241.210 ;
        RECT 1339.585 240.895 1339.915 240.910 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 495.950 53.620 496.270 53.680 ;
        RECT 1346.490 53.620 1346.810 53.680 ;
        RECT 495.950 53.480 1346.810 53.620 ;
        RECT 495.950 53.420 496.270 53.480 ;
        RECT 1346.490 53.420 1346.810 53.480 ;
        RECT 490.430 15.540 490.750 15.600 ;
        RECT 495.950 15.540 496.270 15.600 ;
        RECT 490.430 15.400 496.270 15.540 ;
        RECT 490.430 15.340 490.750 15.400 ;
        RECT 495.950 15.340 496.270 15.400 ;
      LAYER via ;
        RECT 495.980 53.420 496.240 53.680 ;
        RECT 1346.520 53.420 1346.780 53.680 ;
        RECT 490.460 15.340 490.720 15.600 ;
        RECT 495.980 15.340 496.240 15.600 ;
      LAYER met2 ;
        RECT 1350.585 1700.410 1350.865 1704.000 ;
        RECT 1349.340 1700.270 1350.865 1700.410 ;
        RECT 1349.340 1677.970 1349.480 1700.270 ;
        RECT 1350.585 1700.000 1350.865 1700.270 ;
        RECT 1346.580 1677.830 1349.480 1677.970 ;
        RECT 1346.580 53.710 1346.720 1677.830 ;
        RECT 495.980 53.390 496.240 53.710 ;
        RECT 1346.520 53.390 1346.780 53.710 ;
        RECT 496.040 15.630 496.180 53.390 ;
        RECT 490.460 15.310 490.720 15.630 ;
        RECT 495.980 15.310 496.240 15.630 ;
        RECT 490.520 2.400 490.660 15.310 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1353.925 1538.925 1354.095 1587.035 ;
        RECT 1353.925 1449.165 1354.095 1497.275 ;
        RECT 1353.465 1376.405 1353.635 1400.715 ;
        RECT 1353.465 1279.845 1353.635 1304.155 ;
        RECT 1353.465 1062.585 1353.635 1110.695 ;
        RECT 1353.925 565.845 1354.095 613.955 ;
        RECT 1353.465 386.325 1353.635 452.115 ;
        RECT 1353.925 131.325 1354.095 179.435 ;
      LAYER mcon ;
        RECT 1353.925 1586.865 1354.095 1587.035 ;
        RECT 1353.925 1497.105 1354.095 1497.275 ;
        RECT 1353.465 1400.545 1353.635 1400.715 ;
        RECT 1353.465 1303.985 1353.635 1304.155 ;
        RECT 1353.465 1110.525 1353.635 1110.695 ;
        RECT 1353.925 613.785 1354.095 613.955 ;
        RECT 1353.465 451.945 1353.635 452.115 ;
        RECT 1353.925 179.265 1354.095 179.435 ;
      LAYER met1 ;
        RECT 1353.850 1671.680 1354.170 1671.740 ;
        RECT 1356.150 1671.680 1356.470 1671.740 ;
        RECT 1353.850 1671.540 1356.470 1671.680 ;
        RECT 1353.850 1671.480 1354.170 1671.540 ;
        RECT 1356.150 1671.480 1356.470 1671.540 ;
        RECT 1353.850 1587.020 1354.170 1587.080 ;
        RECT 1353.655 1586.880 1354.170 1587.020 ;
        RECT 1353.850 1586.820 1354.170 1586.880 ;
        RECT 1353.850 1539.080 1354.170 1539.140 ;
        RECT 1353.655 1538.940 1354.170 1539.080 ;
        RECT 1353.850 1538.880 1354.170 1538.940 ;
        RECT 1353.850 1497.260 1354.170 1497.320 ;
        RECT 1353.655 1497.120 1354.170 1497.260 ;
        RECT 1353.850 1497.060 1354.170 1497.120 ;
        RECT 1353.850 1449.320 1354.170 1449.380 ;
        RECT 1353.655 1449.180 1354.170 1449.320 ;
        RECT 1353.850 1449.120 1354.170 1449.180 ;
        RECT 1353.850 1414.980 1354.170 1415.040 ;
        RECT 1353.480 1414.840 1354.170 1414.980 ;
        RECT 1353.480 1414.360 1353.620 1414.840 ;
        RECT 1353.850 1414.780 1354.170 1414.840 ;
        RECT 1353.390 1414.100 1353.710 1414.360 ;
        RECT 1353.390 1400.700 1353.710 1400.760 ;
        RECT 1353.195 1400.560 1353.710 1400.700 ;
        RECT 1353.390 1400.500 1353.710 1400.560 ;
        RECT 1353.390 1376.560 1353.710 1376.620 ;
        RECT 1353.195 1376.420 1353.710 1376.560 ;
        RECT 1353.390 1376.360 1353.710 1376.420 ;
        RECT 1353.390 1317.880 1353.710 1318.140 ;
        RECT 1353.480 1317.460 1353.620 1317.880 ;
        RECT 1353.390 1317.200 1353.710 1317.460 ;
        RECT 1353.390 1304.140 1353.710 1304.200 ;
        RECT 1353.195 1304.000 1353.710 1304.140 ;
        RECT 1353.390 1303.940 1353.710 1304.000 ;
        RECT 1353.390 1280.000 1353.710 1280.060 ;
        RECT 1353.195 1279.860 1353.710 1280.000 ;
        RECT 1353.390 1279.800 1353.710 1279.860 ;
        RECT 1353.390 1207.240 1353.710 1207.300 ;
        RECT 1354.310 1207.240 1354.630 1207.300 ;
        RECT 1353.390 1207.100 1354.630 1207.240 ;
        RECT 1353.390 1207.040 1353.710 1207.100 ;
        RECT 1354.310 1207.040 1354.630 1207.100 ;
        RECT 1353.390 1152.500 1353.710 1152.560 ;
        RECT 1353.850 1152.500 1354.170 1152.560 ;
        RECT 1353.390 1152.360 1354.170 1152.500 ;
        RECT 1353.390 1152.300 1353.710 1152.360 ;
        RECT 1353.850 1152.300 1354.170 1152.360 ;
        RECT 1353.390 1124.760 1353.710 1125.020 ;
        RECT 1353.480 1124.340 1353.620 1124.760 ;
        RECT 1353.390 1124.080 1353.710 1124.340 ;
        RECT 1353.390 1110.680 1353.710 1110.740 ;
        RECT 1353.195 1110.540 1353.710 1110.680 ;
        RECT 1353.390 1110.480 1353.710 1110.540 ;
        RECT 1353.405 1062.740 1353.695 1062.785 ;
        RECT 1353.850 1062.740 1354.170 1062.800 ;
        RECT 1353.405 1062.600 1354.170 1062.740 ;
        RECT 1353.405 1062.555 1353.695 1062.600 ;
        RECT 1353.850 1062.540 1354.170 1062.600 ;
        RECT 1352.470 1014.460 1352.790 1014.520 ;
        RECT 1353.390 1014.460 1353.710 1014.520 ;
        RECT 1352.470 1014.320 1353.710 1014.460 ;
        RECT 1352.470 1014.260 1352.790 1014.320 ;
        RECT 1353.390 1014.260 1353.710 1014.320 ;
        RECT 1352.470 966.180 1352.790 966.240 ;
        RECT 1353.850 966.180 1354.170 966.240 ;
        RECT 1352.470 966.040 1354.170 966.180 ;
        RECT 1352.470 965.980 1352.790 966.040 ;
        RECT 1353.850 965.980 1354.170 966.040 ;
        RECT 1352.470 917.900 1352.790 917.960 ;
        RECT 1353.390 917.900 1353.710 917.960 ;
        RECT 1352.470 917.760 1353.710 917.900 ;
        RECT 1352.470 917.700 1352.790 917.760 ;
        RECT 1353.390 917.700 1353.710 917.760 ;
        RECT 1352.470 869.620 1352.790 869.680 ;
        RECT 1353.850 869.620 1354.170 869.680 ;
        RECT 1352.470 869.480 1354.170 869.620 ;
        RECT 1352.470 869.420 1352.790 869.480 ;
        RECT 1353.850 869.420 1354.170 869.480 ;
        RECT 1353.390 820.800 1353.710 821.060 ;
        RECT 1353.480 820.660 1353.620 820.800 ;
        RECT 1353.850 820.660 1354.170 820.720 ;
        RECT 1353.480 820.520 1354.170 820.660 ;
        RECT 1353.850 820.460 1354.170 820.520 ;
        RECT 1353.850 765.920 1354.170 765.980 ;
        RECT 1354.310 765.920 1354.630 765.980 ;
        RECT 1353.850 765.780 1354.630 765.920 ;
        RECT 1353.850 765.720 1354.170 765.780 ;
        RECT 1354.310 765.720 1354.630 765.780 ;
        RECT 1353.850 669.360 1354.170 669.420 ;
        RECT 1355.230 669.360 1355.550 669.420 ;
        RECT 1353.850 669.220 1355.550 669.360 ;
        RECT 1353.850 669.160 1354.170 669.220 ;
        RECT 1355.230 669.160 1355.550 669.220 ;
        RECT 1353.865 613.940 1354.155 613.985 ;
        RECT 1354.310 613.940 1354.630 614.000 ;
        RECT 1353.865 613.800 1354.630 613.940 ;
        RECT 1353.865 613.755 1354.155 613.800 ;
        RECT 1354.310 613.740 1354.630 613.800 ;
        RECT 1353.850 566.000 1354.170 566.060 ;
        RECT 1353.655 565.860 1354.170 566.000 ;
        RECT 1353.850 565.800 1354.170 565.860 ;
        RECT 1353.390 524.520 1353.710 524.580 ;
        RECT 1353.850 524.520 1354.170 524.580 ;
        RECT 1353.390 524.380 1354.170 524.520 ;
        RECT 1353.390 524.320 1353.710 524.380 ;
        RECT 1353.850 524.320 1354.170 524.380 ;
        RECT 1353.390 476.240 1353.710 476.300 ;
        RECT 1353.850 476.240 1354.170 476.300 ;
        RECT 1353.390 476.100 1354.170 476.240 ;
        RECT 1353.390 476.040 1353.710 476.100 ;
        RECT 1353.850 476.040 1354.170 476.100 ;
        RECT 1353.405 452.100 1353.695 452.145 ;
        RECT 1353.850 452.100 1354.170 452.160 ;
        RECT 1353.405 451.960 1354.170 452.100 ;
        RECT 1353.405 451.915 1353.695 451.960 ;
        RECT 1353.850 451.900 1354.170 451.960 ;
        RECT 1353.405 386.480 1353.695 386.525 ;
        RECT 1353.850 386.480 1354.170 386.540 ;
        RECT 1353.405 386.340 1354.170 386.480 ;
        RECT 1353.405 386.295 1353.695 386.340 ;
        RECT 1353.850 386.280 1354.170 386.340 ;
        RECT 1353.850 352.480 1354.170 352.540 ;
        RECT 1353.480 352.340 1354.170 352.480 ;
        RECT 1353.480 351.860 1353.620 352.340 ;
        RECT 1353.850 352.280 1354.170 352.340 ;
        RECT 1353.390 351.600 1353.710 351.860 ;
        RECT 1353.390 290.060 1353.710 290.320 ;
        RECT 1353.480 289.640 1353.620 290.060 ;
        RECT 1353.390 289.380 1353.710 289.640 ;
        RECT 1353.390 193.360 1353.710 193.420 ;
        RECT 1353.850 193.360 1354.170 193.420 ;
        RECT 1353.390 193.220 1354.170 193.360 ;
        RECT 1353.390 193.160 1353.710 193.220 ;
        RECT 1353.850 193.160 1354.170 193.220 ;
        RECT 1353.850 186.220 1354.170 186.280 ;
        RECT 1354.310 186.220 1354.630 186.280 ;
        RECT 1353.850 186.080 1354.630 186.220 ;
        RECT 1353.850 186.020 1354.170 186.080 ;
        RECT 1354.310 186.020 1354.630 186.080 ;
        RECT 1353.865 179.420 1354.155 179.465 ;
        RECT 1354.310 179.420 1354.630 179.480 ;
        RECT 1353.865 179.280 1354.630 179.420 ;
        RECT 1353.865 179.235 1354.155 179.280 ;
        RECT 1354.310 179.220 1354.630 179.280 ;
        RECT 1353.850 131.480 1354.170 131.540 ;
        RECT 1353.655 131.340 1354.170 131.480 ;
        RECT 1353.850 131.280 1354.170 131.340 ;
        RECT 1349.250 110.740 1349.570 110.800 ;
        RECT 1353.390 110.740 1353.710 110.800 ;
        RECT 1349.250 110.600 1353.710 110.740 ;
        RECT 1349.250 110.540 1349.570 110.600 ;
        RECT 1353.390 110.540 1353.710 110.600 ;
        RECT 510.210 53.960 510.530 54.020 ;
        RECT 1349.250 53.960 1349.570 54.020 ;
        RECT 510.210 53.820 1349.570 53.960 ;
        RECT 510.210 53.760 510.530 53.820 ;
        RECT 1349.250 53.760 1349.570 53.820 ;
        RECT 507.910 15.540 508.230 15.600 ;
        RECT 510.210 15.540 510.530 15.600 ;
        RECT 507.910 15.400 510.530 15.540 ;
        RECT 507.910 15.340 508.230 15.400 ;
        RECT 510.210 15.340 510.530 15.400 ;
      LAYER via ;
        RECT 1353.880 1671.480 1354.140 1671.740 ;
        RECT 1356.180 1671.480 1356.440 1671.740 ;
        RECT 1353.880 1586.820 1354.140 1587.080 ;
        RECT 1353.880 1538.880 1354.140 1539.140 ;
        RECT 1353.880 1497.060 1354.140 1497.320 ;
        RECT 1353.880 1449.120 1354.140 1449.380 ;
        RECT 1353.880 1414.780 1354.140 1415.040 ;
        RECT 1353.420 1414.100 1353.680 1414.360 ;
        RECT 1353.420 1400.500 1353.680 1400.760 ;
        RECT 1353.420 1376.360 1353.680 1376.620 ;
        RECT 1353.420 1317.880 1353.680 1318.140 ;
        RECT 1353.420 1317.200 1353.680 1317.460 ;
        RECT 1353.420 1303.940 1353.680 1304.200 ;
        RECT 1353.420 1279.800 1353.680 1280.060 ;
        RECT 1353.420 1207.040 1353.680 1207.300 ;
        RECT 1354.340 1207.040 1354.600 1207.300 ;
        RECT 1353.420 1152.300 1353.680 1152.560 ;
        RECT 1353.880 1152.300 1354.140 1152.560 ;
        RECT 1353.420 1124.760 1353.680 1125.020 ;
        RECT 1353.420 1124.080 1353.680 1124.340 ;
        RECT 1353.420 1110.480 1353.680 1110.740 ;
        RECT 1353.880 1062.540 1354.140 1062.800 ;
        RECT 1352.500 1014.260 1352.760 1014.520 ;
        RECT 1353.420 1014.260 1353.680 1014.520 ;
        RECT 1352.500 965.980 1352.760 966.240 ;
        RECT 1353.880 965.980 1354.140 966.240 ;
        RECT 1352.500 917.700 1352.760 917.960 ;
        RECT 1353.420 917.700 1353.680 917.960 ;
        RECT 1352.500 869.420 1352.760 869.680 ;
        RECT 1353.880 869.420 1354.140 869.680 ;
        RECT 1353.420 820.800 1353.680 821.060 ;
        RECT 1353.880 820.460 1354.140 820.720 ;
        RECT 1353.880 765.720 1354.140 765.980 ;
        RECT 1354.340 765.720 1354.600 765.980 ;
        RECT 1353.880 669.160 1354.140 669.420 ;
        RECT 1355.260 669.160 1355.520 669.420 ;
        RECT 1354.340 613.740 1354.600 614.000 ;
        RECT 1353.880 565.800 1354.140 566.060 ;
        RECT 1353.420 524.320 1353.680 524.580 ;
        RECT 1353.880 524.320 1354.140 524.580 ;
        RECT 1353.420 476.040 1353.680 476.300 ;
        RECT 1353.880 476.040 1354.140 476.300 ;
        RECT 1353.880 451.900 1354.140 452.160 ;
        RECT 1353.880 386.280 1354.140 386.540 ;
        RECT 1353.880 352.280 1354.140 352.540 ;
        RECT 1353.420 351.600 1353.680 351.860 ;
        RECT 1353.420 290.060 1353.680 290.320 ;
        RECT 1353.420 289.380 1353.680 289.640 ;
        RECT 1353.420 193.160 1353.680 193.420 ;
        RECT 1353.880 193.160 1354.140 193.420 ;
        RECT 1353.880 186.020 1354.140 186.280 ;
        RECT 1354.340 186.020 1354.600 186.280 ;
        RECT 1354.340 179.220 1354.600 179.480 ;
        RECT 1353.880 131.280 1354.140 131.540 ;
        RECT 1349.280 110.540 1349.540 110.800 ;
        RECT 1353.420 110.540 1353.680 110.800 ;
        RECT 510.240 53.760 510.500 54.020 ;
        RECT 1349.280 53.760 1349.540 54.020 ;
        RECT 507.940 15.340 508.200 15.600 ;
        RECT 510.240 15.340 510.500 15.600 ;
      LAYER met2 ;
        RECT 1357.945 1700.410 1358.225 1704.000 ;
        RECT 1356.240 1700.270 1358.225 1700.410 ;
        RECT 1356.240 1671.770 1356.380 1700.270 ;
        RECT 1357.945 1700.000 1358.225 1700.270 ;
        RECT 1353.880 1671.450 1354.140 1671.770 ;
        RECT 1356.180 1671.450 1356.440 1671.770 ;
        RECT 1353.940 1587.110 1354.080 1671.450 ;
        RECT 1353.880 1586.790 1354.140 1587.110 ;
        RECT 1353.880 1538.850 1354.140 1539.170 ;
        RECT 1353.940 1497.350 1354.080 1538.850 ;
        RECT 1353.880 1497.030 1354.140 1497.350 ;
        RECT 1353.880 1449.090 1354.140 1449.410 ;
        RECT 1353.940 1415.070 1354.080 1449.090 ;
        RECT 1353.880 1414.750 1354.140 1415.070 ;
        RECT 1353.420 1414.070 1353.680 1414.390 ;
        RECT 1353.480 1400.790 1353.620 1414.070 ;
        RECT 1353.420 1400.470 1353.680 1400.790 ;
        RECT 1353.420 1376.330 1353.680 1376.650 ;
        RECT 1353.480 1318.170 1353.620 1376.330 ;
        RECT 1353.420 1317.850 1353.680 1318.170 ;
        RECT 1353.420 1317.170 1353.680 1317.490 ;
        RECT 1353.480 1304.230 1353.620 1317.170 ;
        RECT 1353.420 1303.910 1353.680 1304.230 ;
        RECT 1353.420 1279.770 1353.680 1280.090 ;
        RECT 1353.480 1207.330 1353.620 1279.770 ;
        RECT 1353.420 1207.010 1353.680 1207.330 ;
        RECT 1354.340 1207.010 1354.600 1207.330 ;
        RECT 1354.400 1200.610 1354.540 1207.010 ;
        RECT 1353.940 1200.470 1354.540 1200.610 ;
        RECT 1353.940 1152.590 1354.080 1200.470 ;
        RECT 1353.420 1152.270 1353.680 1152.590 ;
        RECT 1353.880 1152.270 1354.140 1152.590 ;
        RECT 1353.480 1125.050 1353.620 1152.270 ;
        RECT 1353.420 1124.730 1353.680 1125.050 ;
        RECT 1353.420 1124.050 1353.680 1124.370 ;
        RECT 1353.480 1110.770 1353.620 1124.050 ;
        RECT 1353.420 1110.450 1353.680 1110.770 ;
        RECT 1353.880 1062.685 1354.140 1062.830 ;
        RECT 1352.490 1062.315 1352.770 1062.685 ;
        RECT 1353.870 1062.315 1354.150 1062.685 ;
        RECT 1352.560 1014.550 1352.700 1062.315 ;
        RECT 1352.500 1014.405 1352.760 1014.550 ;
        RECT 1353.420 1014.405 1353.680 1014.550 ;
        RECT 1352.490 1014.035 1352.770 1014.405 ;
        RECT 1353.410 1014.035 1353.690 1014.405 ;
        RECT 1352.560 966.270 1352.700 1014.035 ;
        RECT 1352.500 966.125 1352.760 966.270 ;
        RECT 1353.880 966.125 1354.140 966.270 ;
        RECT 1352.490 965.755 1352.770 966.125 ;
        RECT 1353.870 965.755 1354.150 966.125 ;
        RECT 1352.560 917.990 1352.700 965.755 ;
        RECT 1352.500 917.845 1352.760 917.990 ;
        RECT 1353.420 917.845 1353.680 917.990 ;
        RECT 1352.490 917.475 1352.770 917.845 ;
        RECT 1353.410 917.475 1353.690 917.845 ;
        RECT 1352.560 869.710 1352.700 917.475 ;
        RECT 1352.500 869.390 1352.760 869.710 ;
        RECT 1353.880 869.390 1354.140 869.710 ;
        RECT 1353.940 845.650 1354.080 869.390 ;
        RECT 1353.480 845.510 1354.080 845.650 ;
        RECT 1353.480 821.090 1353.620 845.510 ;
        RECT 1353.420 820.770 1353.680 821.090 ;
        RECT 1353.880 820.430 1354.140 820.750 ;
        RECT 1353.940 766.010 1354.080 820.430 ;
        RECT 1353.880 765.690 1354.140 766.010 ;
        RECT 1354.340 765.690 1354.600 766.010 ;
        RECT 1354.400 689.250 1354.540 765.690 ;
        RECT 1353.940 689.110 1354.540 689.250 ;
        RECT 1353.940 669.450 1354.080 689.110 ;
        RECT 1353.880 669.130 1354.140 669.450 ;
        RECT 1355.260 669.130 1355.520 669.450 ;
        RECT 1355.320 621.250 1355.460 669.130 ;
        RECT 1354.400 621.110 1355.460 621.250 ;
        RECT 1354.400 614.030 1354.540 621.110 ;
        RECT 1354.340 613.710 1354.600 614.030 ;
        RECT 1353.880 565.770 1354.140 566.090 ;
        RECT 1353.940 524.610 1354.080 565.770 ;
        RECT 1353.420 524.290 1353.680 524.610 ;
        RECT 1353.880 524.290 1354.140 524.610 ;
        RECT 1353.480 476.330 1353.620 524.290 ;
        RECT 1353.420 476.010 1353.680 476.330 ;
        RECT 1353.880 476.010 1354.140 476.330 ;
        RECT 1353.940 452.190 1354.080 476.010 ;
        RECT 1353.880 451.870 1354.140 452.190 ;
        RECT 1353.880 386.250 1354.140 386.570 ;
        RECT 1353.940 352.570 1354.080 386.250 ;
        RECT 1353.880 352.250 1354.140 352.570 ;
        RECT 1353.420 351.570 1353.680 351.890 ;
        RECT 1353.480 290.350 1353.620 351.570 ;
        RECT 1353.420 290.030 1353.680 290.350 ;
        RECT 1353.420 289.350 1353.680 289.670 ;
        RECT 1353.480 193.450 1353.620 289.350 ;
        RECT 1353.420 193.130 1353.680 193.450 ;
        RECT 1353.880 193.130 1354.140 193.450 ;
        RECT 1353.940 186.310 1354.080 193.130 ;
        RECT 1353.880 185.990 1354.140 186.310 ;
        RECT 1354.340 185.990 1354.600 186.310 ;
        RECT 1354.400 179.510 1354.540 185.990 ;
        RECT 1354.340 179.190 1354.600 179.510 ;
        RECT 1353.880 131.250 1354.140 131.570 ;
        RECT 1353.940 130.970 1354.080 131.250 ;
        RECT 1353.480 130.830 1354.080 130.970 ;
        RECT 1353.480 110.830 1353.620 130.830 ;
        RECT 1349.280 110.510 1349.540 110.830 ;
        RECT 1353.420 110.510 1353.680 110.830 ;
        RECT 1349.340 54.050 1349.480 110.510 ;
        RECT 510.240 53.730 510.500 54.050 ;
        RECT 1349.280 53.730 1349.540 54.050 ;
        RECT 510.300 15.630 510.440 53.730 ;
        RECT 507.940 15.310 508.200 15.630 ;
        RECT 510.240 15.310 510.500 15.630 ;
        RECT 508.000 2.400 508.140 15.310 ;
        RECT 507.790 -4.800 508.350 2.400 ;
      LAYER via2 ;
        RECT 1352.490 1062.360 1352.770 1062.640 ;
        RECT 1353.870 1062.360 1354.150 1062.640 ;
        RECT 1352.490 1014.080 1352.770 1014.360 ;
        RECT 1353.410 1014.080 1353.690 1014.360 ;
        RECT 1352.490 965.800 1352.770 966.080 ;
        RECT 1353.870 965.800 1354.150 966.080 ;
        RECT 1352.490 917.520 1352.770 917.800 ;
        RECT 1353.410 917.520 1353.690 917.800 ;
      LAYER met3 ;
        RECT 1352.465 1062.650 1352.795 1062.665 ;
        RECT 1353.845 1062.650 1354.175 1062.665 ;
        RECT 1352.465 1062.350 1354.175 1062.650 ;
        RECT 1352.465 1062.335 1352.795 1062.350 ;
        RECT 1353.845 1062.335 1354.175 1062.350 ;
        RECT 1352.465 1014.370 1352.795 1014.385 ;
        RECT 1353.385 1014.370 1353.715 1014.385 ;
        RECT 1352.465 1014.070 1353.715 1014.370 ;
        RECT 1352.465 1014.055 1352.795 1014.070 ;
        RECT 1353.385 1014.055 1353.715 1014.070 ;
        RECT 1352.465 966.090 1352.795 966.105 ;
        RECT 1353.845 966.090 1354.175 966.105 ;
        RECT 1352.465 965.790 1354.175 966.090 ;
        RECT 1352.465 965.775 1352.795 965.790 ;
        RECT 1353.845 965.775 1354.175 965.790 ;
        RECT 1352.465 917.810 1352.795 917.825 ;
        RECT 1353.385 917.810 1353.715 917.825 ;
        RECT 1352.465 917.510 1353.715 917.810 ;
        RECT 1352.465 917.495 1352.795 917.510 ;
        RECT 1353.385 917.495 1353.715 917.510 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1361.285 1538.925 1361.455 1587.035 ;
        RECT 1361.285 1446.445 1361.455 1497.275 ;
        RECT 1361.745 741.285 1361.915 800.275 ;
        RECT 1360.825 386.325 1360.995 452.115 ;
        RECT 1360.825 338.045 1360.995 352.835 ;
        RECT 1360.365 54.145 1360.535 131.155 ;
      LAYER mcon ;
        RECT 1361.285 1586.865 1361.455 1587.035 ;
        RECT 1361.285 1497.105 1361.455 1497.275 ;
        RECT 1361.745 800.105 1361.915 800.275 ;
        RECT 1360.825 451.945 1360.995 452.115 ;
        RECT 1360.825 352.665 1360.995 352.835 ;
        RECT 1360.365 130.985 1360.535 131.155 ;
      LAYER met1 ;
        RECT 1361.210 1671.680 1361.530 1671.740 ;
        RECT 1363.510 1671.680 1363.830 1671.740 ;
        RECT 1361.210 1671.540 1363.830 1671.680 ;
        RECT 1361.210 1671.480 1361.530 1671.540 ;
        RECT 1363.510 1671.480 1363.830 1671.540 ;
        RECT 1361.210 1587.020 1361.530 1587.080 ;
        RECT 1361.015 1586.880 1361.530 1587.020 ;
        RECT 1361.210 1586.820 1361.530 1586.880 ;
        RECT 1361.210 1539.080 1361.530 1539.140 ;
        RECT 1361.015 1538.940 1361.530 1539.080 ;
        RECT 1361.210 1538.880 1361.530 1538.940 ;
        RECT 1361.210 1497.260 1361.530 1497.320 ;
        RECT 1361.015 1497.120 1361.530 1497.260 ;
        RECT 1361.210 1497.060 1361.530 1497.120 ;
        RECT 1361.210 1446.600 1361.530 1446.660 ;
        RECT 1361.015 1446.460 1361.530 1446.600 ;
        RECT 1361.210 1446.400 1361.530 1446.460 ;
        RECT 1361.210 1441.840 1361.530 1441.900 ;
        RECT 1361.670 1441.840 1361.990 1441.900 ;
        RECT 1361.210 1441.700 1361.990 1441.840 ;
        RECT 1361.210 1441.640 1361.530 1441.700 ;
        RECT 1361.670 1441.640 1361.990 1441.700 ;
        RECT 1361.670 1304.820 1361.990 1304.880 ;
        RECT 1360.840 1304.680 1361.990 1304.820 ;
        RECT 1360.840 1303.860 1360.980 1304.680 ;
        RECT 1361.670 1304.620 1361.990 1304.680 ;
        RECT 1360.750 1303.600 1361.070 1303.860 ;
        RECT 1360.750 1207.240 1361.070 1207.300 ;
        RECT 1361.670 1207.240 1361.990 1207.300 ;
        RECT 1360.750 1207.100 1361.990 1207.240 ;
        RECT 1360.750 1207.040 1361.070 1207.100 ;
        RECT 1361.670 1207.040 1361.990 1207.100 ;
        RECT 1360.750 1110.680 1361.070 1110.740 ;
        RECT 1361.210 1110.680 1361.530 1110.740 ;
        RECT 1360.750 1110.540 1361.530 1110.680 ;
        RECT 1360.750 1110.480 1361.070 1110.540 ;
        RECT 1361.210 1110.480 1361.530 1110.540 ;
        RECT 1360.290 910.760 1360.610 910.820 ;
        RECT 1361.670 910.760 1361.990 910.820 ;
        RECT 1360.290 910.620 1361.990 910.760 ;
        RECT 1360.290 910.560 1360.610 910.620 ;
        RECT 1361.670 910.560 1361.990 910.620 ;
        RECT 1360.750 800.260 1361.070 800.320 ;
        RECT 1361.685 800.260 1361.975 800.305 ;
        RECT 1360.750 800.120 1361.975 800.260 ;
        RECT 1360.750 800.060 1361.070 800.120 ;
        RECT 1361.685 800.075 1361.975 800.120 ;
        RECT 1361.670 741.440 1361.990 741.500 ;
        RECT 1361.475 741.300 1361.990 741.440 ;
        RECT 1361.670 741.240 1361.990 741.300 ;
        RECT 1361.210 572.460 1361.530 572.520 ;
        RECT 1361.670 572.460 1361.990 572.520 ;
        RECT 1361.210 572.320 1361.990 572.460 ;
        RECT 1361.210 572.260 1361.530 572.320 ;
        RECT 1361.670 572.260 1361.990 572.320 ;
        RECT 1361.670 476.380 1361.990 476.640 ;
        RECT 1361.210 476.240 1361.530 476.300 ;
        RECT 1361.760 476.240 1361.900 476.380 ;
        RECT 1361.210 476.100 1361.900 476.240 ;
        RECT 1361.210 476.040 1361.530 476.100 ;
        RECT 1360.765 452.100 1361.055 452.145 ;
        RECT 1361.210 452.100 1361.530 452.160 ;
        RECT 1360.765 451.960 1361.530 452.100 ;
        RECT 1360.765 451.915 1361.055 451.960 ;
        RECT 1361.210 451.900 1361.530 451.960 ;
        RECT 1360.765 386.480 1361.055 386.525 ;
        RECT 1361.210 386.480 1361.530 386.540 ;
        RECT 1360.765 386.340 1361.530 386.480 ;
        RECT 1360.765 386.295 1361.055 386.340 ;
        RECT 1361.210 386.280 1361.530 386.340 ;
        RECT 1360.765 352.820 1361.055 352.865 ;
        RECT 1361.210 352.820 1361.530 352.880 ;
        RECT 1360.765 352.680 1361.530 352.820 ;
        RECT 1360.765 352.635 1361.055 352.680 ;
        RECT 1361.210 352.620 1361.530 352.680 ;
        RECT 1360.750 338.200 1361.070 338.260 ;
        RECT 1360.555 338.060 1361.070 338.200 ;
        RECT 1360.750 338.000 1361.070 338.060 ;
        RECT 1360.750 289.920 1361.070 289.980 ;
        RECT 1361.210 289.920 1361.530 289.980 ;
        RECT 1360.750 289.780 1361.530 289.920 ;
        RECT 1360.750 289.720 1361.070 289.780 ;
        RECT 1361.210 289.720 1361.530 289.780 ;
        RECT 1360.750 193.360 1361.070 193.420 ;
        RECT 1361.210 193.360 1361.530 193.420 ;
        RECT 1360.750 193.220 1361.530 193.360 ;
        RECT 1360.750 193.160 1361.070 193.220 ;
        RECT 1361.210 193.160 1361.530 193.220 ;
        RECT 1360.305 131.140 1360.595 131.185 ;
        RECT 1361.210 131.140 1361.530 131.200 ;
        RECT 1360.305 131.000 1361.530 131.140 ;
        RECT 1360.305 130.955 1360.595 131.000 ;
        RECT 1361.210 130.940 1361.530 131.000 ;
        RECT 530.910 54.300 531.230 54.360 ;
        RECT 1360.305 54.300 1360.595 54.345 ;
        RECT 530.910 54.160 1360.595 54.300 ;
        RECT 530.910 54.100 531.230 54.160 ;
        RECT 1360.305 54.115 1360.595 54.160 ;
        RECT 525.850 15.540 526.170 15.600 ;
        RECT 530.910 15.540 531.230 15.600 ;
        RECT 525.850 15.400 531.230 15.540 ;
        RECT 525.850 15.340 526.170 15.400 ;
        RECT 530.910 15.340 531.230 15.400 ;
      LAYER via ;
        RECT 1361.240 1671.480 1361.500 1671.740 ;
        RECT 1363.540 1671.480 1363.800 1671.740 ;
        RECT 1361.240 1586.820 1361.500 1587.080 ;
        RECT 1361.240 1538.880 1361.500 1539.140 ;
        RECT 1361.240 1497.060 1361.500 1497.320 ;
        RECT 1361.240 1446.400 1361.500 1446.660 ;
        RECT 1361.240 1441.640 1361.500 1441.900 ;
        RECT 1361.700 1441.640 1361.960 1441.900 ;
        RECT 1361.700 1304.620 1361.960 1304.880 ;
        RECT 1360.780 1303.600 1361.040 1303.860 ;
        RECT 1360.780 1207.040 1361.040 1207.300 ;
        RECT 1361.700 1207.040 1361.960 1207.300 ;
        RECT 1360.780 1110.480 1361.040 1110.740 ;
        RECT 1361.240 1110.480 1361.500 1110.740 ;
        RECT 1360.320 910.560 1360.580 910.820 ;
        RECT 1361.700 910.560 1361.960 910.820 ;
        RECT 1360.780 800.060 1361.040 800.320 ;
        RECT 1361.700 741.240 1361.960 741.500 ;
        RECT 1361.240 572.260 1361.500 572.520 ;
        RECT 1361.700 572.260 1361.960 572.520 ;
        RECT 1361.700 476.380 1361.960 476.640 ;
        RECT 1361.240 476.040 1361.500 476.300 ;
        RECT 1361.240 451.900 1361.500 452.160 ;
        RECT 1361.240 386.280 1361.500 386.540 ;
        RECT 1361.240 352.620 1361.500 352.880 ;
        RECT 1360.780 338.000 1361.040 338.260 ;
        RECT 1360.780 289.720 1361.040 289.980 ;
        RECT 1361.240 289.720 1361.500 289.980 ;
        RECT 1360.780 193.160 1361.040 193.420 ;
        RECT 1361.240 193.160 1361.500 193.420 ;
        RECT 1361.240 130.940 1361.500 131.200 ;
        RECT 530.940 54.100 531.200 54.360 ;
        RECT 525.880 15.340 526.140 15.600 ;
        RECT 530.940 15.340 531.200 15.600 ;
      LAYER met2 ;
        RECT 1365.305 1700.410 1365.585 1704.000 ;
        RECT 1363.600 1700.270 1365.585 1700.410 ;
        RECT 1363.600 1671.770 1363.740 1700.270 ;
        RECT 1365.305 1700.000 1365.585 1700.270 ;
        RECT 1361.240 1671.450 1361.500 1671.770 ;
        RECT 1363.540 1671.450 1363.800 1671.770 ;
        RECT 1361.300 1587.110 1361.440 1671.450 ;
        RECT 1361.240 1586.790 1361.500 1587.110 ;
        RECT 1361.240 1538.850 1361.500 1539.170 ;
        RECT 1361.300 1497.350 1361.440 1538.850 ;
        RECT 1361.240 1497.030 1361.500 1497.350 ;
        RECT 1361.240 1446.370 1361.500 1446.690 ;
        RECT 1361.300 1441.930 1361.440 1446.370 ;
        RECT 1361.240 1441.610 1361.500 1441.930 ;
        RECT 1361.700 1441.610 1361.960 1441.930 ;
        RECT 1361.760 1393.845 1361.900 1441.610 ;
        RECT 1360.770 1393.475 1361.050 1393.845 ;
        RECT 1361.690 1393.475 1361.970 1393.845 ;
        RECT 1360.840 1350.210 1360.980 1393.475 ;
        RECT 1360.840 1350.070 1361.900 1350.210 ;
        RECT 1361.760 1304.910 1361.900 1350.070 ;
        RECT 1361.700 1304.590 1361.960 1304.910 ;
        RECT 1360.780 1303.570 1361.040 1303.890 ;
        RECT 1360.840 1207.330 1360.980 1303.570 ;
        RECT 1360.780 1207.010 1361.040 1207.330 ;
        RECT 1361.700 1207.010 1361.960 1207.330 ;
        RECT 1361.760 1200.725 1361.900 1207.010 ;
        RECT 1360.770 1200.355 1361.050 1200.725 ;
        RECT 1361.690 1200.355 1361.970 1200.725 ;
        RECT 1360.840 1157.770 1360.980 1200.355 ;
        RECT 1360.840 1157.630 1361.900 1157.770 ;
        RECT 1361.760 1124.450 1361.900 1157.630 ;
        RECT 1360.840 1124.310 1361.900 1124.450 ;
        RECT 1360.840 1110.770 1360.980 1124.310 ;
        RECT 1360.780 1110.450 1361.040 1110.770 ;
        RECT 1361.240 1110.450 1361.500 1110.770 ;
        RECT 1361.300 1104.165 1361.440 1110.450 ;
        RECT 1360.310 1103.795 1360.590 1104.165 ;
        RECT 1361.230 1103.795 1361.510 1104.165 ;
        RECT 1360.380 1055.885 1360.520 1103.795 ;
        RECT 1360.310 1055.515 1360.590 1055.885 ;
        RECT 1361.230 1055.515 1361.510 1055.885 ;
        RECT 1361.300 1038.770 1361.440 1055.515 ;
        RECT 1360.380 1038.630 1361.440 1038.770 ;
        RECT 1360.380 1027.890 1360.520 1038.630 ;
        RECT 1360.380 1027.750 1360.980 1027.890 ;
        RECT 1360.840 1014.405 1360.980 1027.750 ;
        RECT 1360.770 1014.035 1361.050 1014.405 ;
        RECT 1361.690 1013.355 1361.970 1013.725 ;
        RECT 1361.760 966.010 1361.900 1013.355 ;
        RECT 1360.380 965.870 1361.900 966.010 ;
        RECT 1360.380 931.330 1360.520 965.870 ;
        RECT 1360.380 931.190 1360.980 931.330 ;
        RECT 1360.840 917.845 1360.980 931.190 ;
        RECT 1360.770 917.475 1361.050 917.845 ;
        RECT 1361.690 916.795 1361.970 917.165 ;
        RECT 1361.760 910.850 1361.900 916.795 ;
        RECT 1360.320 910.530 1360.580 910.850 ;
        RECT 1361.700 910.530 1361.960 910.850 ;
        RECT 1360.380 862.765 1360.520 910.530 ;
        RECT 1360.310 862.395 1360.590 862.765 ;
        RECT 1361.230 862.395 1361.510 862.765 ;
        RECT 1361.300 831.370 1361.440 862.395 ;
        RECT 1360.840 831.230 1361.440 831.370 ;
        RECT 1360.840 800.350 1360.980 831.230 ;
        RECT 1360.780 800.030 1361.040 800.350 ;
        RECT 1361.700 741.210 1361.960 741.530 ;
        RECT 1361.760 699.450 1361.900 741.210 ;
        RECT 1361.300 699.310 1361.900 699.450 ;
        RECT 1361.300 628.845 1361.440 699.310 ;
        RECT 1361.230 628.475 1361.510 628.845 ;
        RECT 1360.770 627.795 1361.050 628.165 ;
        RECT 1360.840 596.770 1360.980 627.795 ;
        RECT 1360.840 596.630 1361.440 596.770 ;
        RECT 1361.300 572.550 1361.440 596.630 ;
        RECT 1361.240 572.230 1361.500 572.550 ;
        RECT 1361.700 572.230 1361.960 572.550 ;
        RECT 1361.760 476.670 1361.900 572.230 ;
        RECT 1361.700 476.350 1361.960 476.670 ;
        RECT 1361.240 476.010 1361.500 476.330 ;
        RECT 1361.300 452.190 1361.440 476.010 ;
        RECT 1361.240 451.870 1361.500 452.190 ;
        RECT 1361.240 386.250 1361.500 386.570 ;
        RECT 1361.300 352.910 1361.440 386.250 ;
        RECT 1361.240 352.590 1361.500 352.910 ;
        RECT 1360.780 337.970 1361.040 338.290 ;
        RECT 1360.840 290.010 1360.980 337.970 ;
        RECT 1360.780 289.690 1361.040 290.010 ;
        RECT 1361.240 289.690 1361.500 290.010 ;
        RECT 1361.300 265.610 1361.440 289.690 ;
        RECT 1360.840 265.470 1361.440 265.610 ;
        RECT 1360.840 193.450 1360.980 265.470 ;
        RECT 1360.780 193.130 1361.040 193.450 ;
        RECT 1361.240 193.130 1361.500 193.450 ;
        RECT 1361.300 131.230 1361.440 193.130 ;
        RECT 1361.240 130.910 1361.500 131.230 ;
        RECT 530.940 54.070 531.200 54.390 ;
        RECT 531.000 15.630 531.140 54.070 ;
        RECT 525.880 15.310 526.140 15.630 ;
        RECT 530.940 15.310 531.200 15.630 ;
        RECT 525.940 2.400 526.080 15.310 ;
        RECT 525.730 -4.800 526.290 2.400 ;
      LAYER via2 ;
        RECT 1360.770 1393.520 1361.050 1393.800 ;
        RECT 1361.690 1393.520 1361.970 1393.800 ;
        RECT 1360.770 1200.400 1361.050 1200.680 ;
        RECT 1361.690 1200.400 1361.970 1200.680 ;
        RECT 1360.310 1103.840 1360.590 1104.120 ;
        RECT 1361.230 1103.840 1361.510 1104.120 ;
        RECT 1360.310 1055.560 1360.590 1055.840 ;
        RECT 1361.230 1055.560 1361.510 1055.840 ;
        RECT 1360.770 1014.080 1361.050 1014.360 ;
        RECT 1361.690 1013.400 1361.970 1013.680 ;
        RECT 1360.770 917.520 1361.050 917.800 ;
        RECT 1361.690 916.840 1361.970 917.120 ;
        RECT 1360.310 862.440 1360.590 862.720 ;
        RECT 1361.230 862.440 1361.510 862.720 ;
        RECT 1361.230 628.520 1361.510 628.800 ;
        RECT 1360.770 627.840 1361.050 628.120 ;
      LAYER met3 ;
        RECT 1360.745 1393.810 1361.075 1393.825 ;
        RECT 1361.665 1393.810 1361.995 1393.825 ;
        RECT 1360.745 1393.510 1361.995 1393.810 ;
        RECT 1360.745 1393.495 1361.075 1393.510 ;
        RECT 1361.665 1393.495 1361.995 1393.510 ;
        RECT 1360.745 1200.690 1361.075 1200.705 ;
        RECT 1361.665 1200.690 1361.995 1200.705 ;
        RECT 1360.745 1200.390 1361.995 1200.690 ;
        RECT 1360.745 1200.375 1361.075 1200.390 ;
        RECT 1361.665 1200.375 1361.995 1200.390 ;
        RECT 1360.285 1104.130 1360.615 1104.145 ;
        RECT 1361.205 1104.130 1361.535 1104.145 ;
        RECT 1360.285 1103.830 1361.535 1104.130 ;
        RECT 1360.285 1103.815 1360.615 1103.830 ;
        RECT 1361.205 1103.815 1361.535 1103.830 ;
        RECT 1360.285 1055.850 1360.615 1055.865 ;
        RECT 1361.205 1055.850 1361.535 1055.865 ;
        RECT 1360.285 1055.550 1361.535 1055.850 ;
        RECT 1360.285 1055.535 1360.615 1055.550 ;
        RECT 1361.205 1055.535 1361.535 1055.550 ;
        RECT 1360.745 1014.370 1361.075 1014.385 ;
        RECT 1360.070 1014.070 1361.075 1014.370 ;
        RECT 1360.070 1013.690 1360.370 1014.070 ;
        RECT 1360.745 1014.055 1361.075 1014.070 ;
        RECT 1361.665 1013.690 1361.995 1013.705 ;
        RECT 1360.070 1013.390 1361.995 1013.690 ;
        RECT 1361.665 1013.375 1361.995 1013.390 ;
        RECT 1360.745 917.810 1361.075 917.825 ;
        RECT 1360.070 917.510 1361.075 917.810 ;
        RECT 1360.070 917.130 1360.370 917.510 ;
        RECT 1360.745 917.495 1361.075 917.510 ;
        RECT 1361.665 917.130 1361.995 917.145 ;
        RECT 1360.070 916.830 1361.995 917.130 ;
        RECT 1361.665 916.815 1361.995 916.830 ;
        RECT 1360.285 862.730 1360.615 862.745 ;
        RECT 1361.205 862.730 1361.535 862.745 ;
        RECT 1360.285 862.430 1361.535 862.730 ;
        RECT 1360.285 862.415 1360.615 862.430 ;
        RECT 1361.205 862.415 1361.535 862.430 ;
        RECT 1361.205 628.810 1361.535 628.825 ;
        RECT 1360.990 628.495 1361.535 628.810 ;
        RECT 1360.990 628.145 1361.290 628.495 ;
        RECT 1360.745 627.830 1361.290 628.145 ;
        RECT 1360.745 627.815 1361.075 627.830 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1367.725 1587.545 1367.895 1608.795 ;
        RECT 1367.725 1352.605 1367.895 1400.715 ;
        RECT 1367.725 1256.045 1367.895 1304.155 ;
        RECT 1367.725 862.665 1367.895 910.775 ;
        RECT 1367.725 724.285 1367.895 765.935 ;
        RECT 1367.725 379.525 1367.895 400.095 ;
        RECT 1367.725 282.965 1367.895 331.075 ;
        RECT 1367.265 54.485 1367.435 89.675 ;
      LAYER mcon ;
        RECT 1367.725 1608.625 1367.895 1608.795 ;
        RECT 1367.725 1400.545 1367.895 1400.715 ;
        RECT 1367.725 1303.985 1367.895 1304.155 ;
        RECT 1367.725 910.605 1367.895 910.775 ;
        RECT 1367.725 765.765 1367.895 765.935 ;
        RECT 1367.725 399.925 1367.895 400.095 ;
        RECT 1367.725 330.905 1367.895 331.075 ;
        RECT 1367.265 89.505 1367.435 89.675 ;
      LAYER met1 ;
        RECT 1367.650 1608.780 1367.970 1608.840 ;
        RECT 1367.455 1608.640 1367.970 1608.780 ;
        RECT 1367.650 1608.580 1367.970 1608.640 ;
        RECT 1367.650 1587.700 1367.970 1587.760 ;
        RECT 1367.455 1587.560 1367.970 1587.700 ;
        RECT 1367.650 1587.500 1367.970 1587.560 ;
        RECT 1367.650 1587.020 1367.970 1587.080 ;
        RECT 1367.650 1586.880 1368.340 1587.020 ;
        RECT 1367.650 1586.820 1367.970 1586.880 ;
        RECT 1368.200 1586.740 1368.340 1586.880 ;
        RECT 1368.110 1586.480 1368.430 1586.740 ;
        RECT 1367.650 1497.060 1367.970 1497.320 ;
        RECT 1367.740 1496.640 1367.880 1497.060 ;
        RECT 1367.650 1496.380 1367.970 1496.640 ;
        RECT 1367.650 1400.700 1367.970 1400.760 ;
        RECT 1367.455 1400.560 1367.970 1400.700 ;
        RECT 1367.650 1400.500 1367.970 1400.560 ;
        RECT 1367.650 1352.760 1367.970 1352.820 ;
        RECT 1367.455 1352.620 1367.970 1352.760 ;
        RECT 1367.650 1352.560 1367.970 1352.620 ;
        RECT 1367.650 1304.140 1367.970 1304.200 ;
        RECT 1367.455 1304.000 1367.970 1304.140 ;
        RECT 1367.650 1303.940 1367.970 1304.000 ;
        RECT 1367.650 1256.200 1367.970 1256.260 ;
        RECT 1367.455 1256.060 1367.970 1256.200 ;
        RECT 1367.650 1256.000 1367.970 1256.060 ;
        RECT 1367.650 1159.300 1367.970 1159.360 ;
        RECT 1368.570 1159.300 1368.890 1159.360 ;
        RECT 1367.650 1159.160 1368.890 1159.300 ;
        RECT 1367.650 1159.100 1367.970 1159.160 ;
        RECT 1368.570 1159.100 1368.890 1159.160 ;
        RECT 1367.650 1062.740 1367.970 1062.800 ;
        RECT 1368.570 1062.740 1368.890 1062.800 ;
        RECT 1367.650 1062.600 1368.890 1062.740 ;
        RECT 1367.650 1062.540 1367.970 1062.600 ;
        RECT 1368.570 1062.540 1368.890 1062.600 ;
        RECT 1367.650 966.180 1367.970 966.240 ;
        RECT 1368.570 966.180 1368.890 966.240 ;
        RECT 1367.650 966.040 1368.890 966.180 ;
        RECT 1367.650 965.980 1367.970 966.040 ;
        RECT 1368.570 965.980 1368.890 966.040 ;
        RECT 1367.665 910.760 1367.955 910.805 ;
        RECT 1368.570 910.760 1368.890 910.820 ;
        RECT 1367.665 910.620 1368.890 910.760 ;
        RECT 1367.665 910.575 1367.955 910.620 ;
        RECT 1368.570 910.560 1368.890 910.620 ;
        RECT 1367.650 862.820 1367.970 862.880 ;
        RECT 1367.455 862.680 1367.970 862.820 ;
        RECT 1367.650 862.620 1367.970 862.680 ;
        RECT 1367.650 765.920 1367.970 765.980 ;
        RECT 1367.455 765.780 1367.970 765.920 ;
        RECT 1367.650 765.720 1367.970 765.780 ;
        RECT 1367.650 724.440 1367.970 724.500 ;
        RECT 1367.455 724.300 1367.970 724.440 ;
        RECT 1367.650 724.240 1367.970 724.300 ;
        RECT 1367.650 676.500 1367.970 676.560 ;
        RECT 1368.110 676.500 1368.430 676.560 ;
        RECT 1367.650 676.360 1368.430 676.500 ;
        RECT 1367.650 676.300 1367.970 676.360 ;
        RECT 1368.110 676.300 1368.430 676.360 ;
        RECT 1367.650 400.080 1367.970 400.140 ;
        RECT 1367.455 399.940 1367.970 400.080 ;
        RECT 1367.650 399.880 1367.970 399.940 ;
        RECT 1367.650 379.680 1367.970 379.740 ;
        RECT 1367.455 379.540 1367.970 379.680 ;
        RECT 1367.650 379.480 1367.970 379.540 ;
        RECT 1367.650 331.060 1367.970 331.120 ;
        RECT 1367.455 330.920 1367.970 331.060 ;
        RECT 1367.650 330.860 1367.970 330.920 ;
        RECT 1367.650 283.120 1367.970 283.180 ;
        RECT 1367.455 282.980 1367.970 283.120 ;
        RECT 1367.650 282.920 1367.970 282.980 ;
        RECT 1367.650 255.380 1367.970 255.640 ;
        RECT 1367.740 254.620 1367.880 255.380 ;
        RECT 1367.650 254.360 1367.970 254.620 ;
        RECT 1367.190 89.660 1367.510 89.720 ;
        RECT 1366.995 89.520 1367.510 89.660 ;
        RECT 1367.190 89.460 1367.510 89.520 ;
        RECT 544.710 54.640 545.030 54.700 ;
        RECT 1367.205 54.640 1367.495 54.685 ;
        RECT 544.710 54.500 1367.495 54.640 ;
        RECT 544.710 54.440 545.030 54.500 ;
        RECT 1367.205 54.455 1367.495 54.500 ;
      LAYER via ;
        RECT 1367.680 1608.580 1367.940 1608.840 ;
        RECT 1367.680 1587.500 1367.940 1587.760 ;
        RECT 1367.680 1586.820 1367.940 1587.080 ;
        RECT 1368.140 1586.480 1368.400 1586.740 ;
        RECT 1367.680 1497.060 1367.940 1497.320 ;
        RECT 1367.680 1496.380 1367.940 1496.640 ;
        RECT 1367.680 1400.500 1367.940 1400.760 ;
        RECT 1367.680 1352.560 1367.940 1352.820 ;
        RECT 1367.680 1303.940 1367.940 1304.200 ;
        RECT 1367.680 1256.000 1367.940 1256.260 ;
        RECT 1367.680 1159.100 1367.940 1159.360 ;
        RECT 1368.600 1159.100 1368.860 1159.360 ;
        RECT 1367.680 1062.540 1367.940 1062.800 ;
        RECT 1368.600 1062.540 1368.860 1062.800 ;
        RECT 1367.680 965.980 1367.940 966.240 ;
        RECT 1368.600 965.980 1368.860 966.240 ;
        RECT 1368.600 910.560 1368.860 910.820 ;
        RECT 1367.680 862.620 1367.940 862.880 ;
        RECT 1367.680 765.720 1367.940 765.980 ;
        RECT 1367.680 724.240 1367.940 724.500 ;
        RECT 1367.680 676.300 1367.940 676.560 ;
        RECT 1368.140 676.300 1368.400 676.560 ;
        RECT 1367.680 399.880 1367.940 400.140 ;
        RECT 1367.680 379.480 1367.940 379.740 ;
        RECT 1367.680 330.860 1367.940 331.120 ;
        RECT 1367.680 282.920 1367.940 283.180 ;
        RECT 1367.680 255.380 1367.940 255.640 ;
        RECT 1367.680 254.360 1367.940 254.620 ;
        RECT 1367.220 89.460 1367.480 89.720 ;
        RECT 544.740 54.440 545.000 54.700 ;
      LAYER met2 ;
        RECT 1372.665 1700.410 1372.945 1704.000 ;
        RECT 1371.420 1700.270 1372.945 1700.410 ;
        RECT 1371.420 1656.210 1371.560 1700.270 ;
        RECT 1372.665 1700.000 1372.945 1700.270 ;
        RECT 1367.740 1656.070 1371.560 1656.210 ;
        RECT 1367.740 1608.870 1367.880 1656.070 ;
        RECT 1367.680 1608.550 1367.940 1608.870 ;
        RECT 1367.680 1587.470 1367.940 1587.790 ;
        RECT 1367.740 1587.110 1367.880 1587.470 ;
        RECT 1367.680 1586.790 1367.940 1587.110 ;
        RECT 1368.140 1586.450 1368.400 1586.770 ;
        RECT 1368.200 1545.370 1368.340 1586.450 ;
        RECT 1367.740 1545.230 1368.340 1545.370 ;
        RECT 1367.740 1497.350 1367.880 1545.230 ;
        RECT 1367.680 1497.030 1367.940 1497.350 ;
        RECT 1367.680 1496.350 1367.940 1496.670 ;
        RECT 1367.740 1400.790 1367.880 1496.350 ;
        RECT 1367.680 1400.470 1367.940 1400.790 ;
        RECT 1367.680 1352.530 1367.940 1352.850 ;
        RECT 1367.740 1304.230 1367.880 1352.530 ;
        RECT 1367.680 1303.910 1367.940 1304.230 ;
        RECT 1367.680 1255.970 1367.940 1256.290 ;
        RECT 1367.740 1207.525 1367.880 1255.970 ;
        RECT 1367.670 1207.155 1367.950 1207.525 ;
        RECT 1368.590 1207.155 1368.870 1207.525 ;
        RECT 1368.660 1159.390 1368.800 1207.155 ;
        RECT 1367.680 1159.070 1367.940 1159.390 ;
        RECT 1368.600 1159.070 1368.860 1159.390 ;
        RECT 1367.740 1110.965 1367.880 1159.070 ;
        RECT 1367.670 1110.595 1367.950 1110.965 ;
        RECT 1368.590 1110.595 1368.870 1110.965 ;
        RECT 1368.660 1062.830 1368.800 1110.595 ;
        RECT 1367.680 1062.510 1367.940 1062.830 ;
        RECT 1368.600 1062.510 1368.860 1062.830 ;
        RECT 1367.740 1014.405 1367.880 1062.510 ;
        RECT 1367.670 1014.035 1367.950 1014.405 ;
        RECT 1368.590 1014.035 1368.870 1014.405 ;
        RECT 1368.660 966.270 1368.800 1014.035 ;
        RECT 1367.680 965.950 1367.940 966.270 ;
        RECT 1368.600 965.950 1368.860 966.270 ;
        RECT 1367.740 917.845 1367.880 965.950 ;
        RECT 1367.670 917.475 1367.950 917.845 ;
        RECT 1368.590 917.475 1368.870 917.845 ;
        RECT 1368.660 910.850 1368.800 917.475 ;
        RECT 1368.600 910.530 1368.860 910.850 ;
        RECT 1367.680 862.590 1367.940 862.910 ;
        RECT 1367.740 766.010 1367.880 862.590 ;
        RECT 1367.680 765.690 1367.940 766.010 ;
        RECT 1367.680 724.210 1367.940 724.530 ;
        RECT 1367.740 717.810 1367.880 724.210 ;
        RECT 1367.740 717.670 1368.340 717.810 ;
        RECT 1368.200 676.590 1368.340 717.670 ;
        RECT 1367.680 676.270 1367.940 676.590 ;
        RECT 1368.140 676.270 1368.400 676.590 ;
        RECT 1367.740 628.845 1367.880 676.270 ;
        RECT 1367.670 628.475 1367.950 628.845 ;
        RECT 1367.670 627.795 1367.950 628.165 ;
        RECT 1367.740 594.050 1367.880 627.795 ;
        RECT 1367.740 593.910 1368.340 594.050 ;
        RECT 1368.200 592.690 1368.340 593.910 ;
        RECT 1367.740 592.550 1368.340 592.690 ;
        RECT 1367.740 497.490 1367.880 592.550 ;
        RECT 1367.280 497.350 1367.880 497.490 ;
        RECT 1367.280 496.810 1367.420 497.350 ;
        RECT 1367.280 496.670 1367.880 496.810 ;
        RECT 1367.740 400.170 1367.880 496.670 ;
        RECT 1367.680 399.850 1367.940 400.170 ;
        RECT 1367.680 379.450 1367.940 379.770 ;
        RECT 1367.740 331.150 1367.880 379.450 ;
        RECT 1367.680 330.830 1367.940 331.150 ;
        RECT 1367.680 282.890 1367.940 283.210 ;
        RECT 1367.740 255.670 1367.880 282.890 ;
        RECT 1367.680 255.350 1367.940 255.670 ;
        RECT 1367.680 254.330 1367.940 254.650 ;
        RECT 1367.740 110.570 1367.880 254.330 ;
        RECT 1367.280 110.430 1367.880 110.570 ;
        RECT 1367.280 89.750 1367.420 110.430 ;
        RECT 1367.220 89.430 1367.480 89.750 ;
        RECT 544.740 54.410 545.000 54.730 ;
        RECT 544.800 17.410 544.940 54.410 ;
        RECT 543.880 17.270 544.940 17.410 ;
        RECT 543.880 2.400 544.020 17.270 ;
        RECT 543.670 -4.800 544.230 2.400 ;
      LAYER via2 ;
        RECT 1367.670 1207.200 1367.950 1207.480 ;
        RECT 1368.590 1207.200 1368.870 1207.480 ;
        RECT 1367.670 1110.640 1367.950 1110.920 ;
        RECT 1368.590 1110.640 1368.870 1110.920 ;
        RECT 1367.670 1014.080 1367.950 1014.360 ;
        RECT 1368.590 1014.080 1368.870 1014.360 ;
        RECT 1367.670 917.520 1367.950 917.800 ;
        RECT 1368.590 917.520 1368.870 917.800 ;
        RECT 1367.670 628.520 1367.950 628.800 ;
        RECT 1367.670 627.840 1367.950 628.120 ;
      LAYER met3 ;
        RECT 1367.645 1207.490 1367.975 1207.505 ;
        RECT 1368.565 1207.490 1368.895 1207.505 ;
        RECT 1367.645 1207.190 1368.895 1207.490 ;
        RECT 1367.645 1207.175 1367.975 1207.190 ;
        RECT 1368.565 1207.175 1368.895 1207.190 ;
        RECT 1367.645 1110.930 1367.975 1110.945 ;
        RECT 1368.565 1110.930 1368.895 1110.945 ;
        RECT 1367.645 1110.630 1368.895 1110.930 ;
        RECT 1367.645 1110.615 1367.975 1110.630 ;
        RECT 1368.565 1110.615 1368.895 1110.630 ;
        RECT 1367.645 1014.370 1367.975 1014.385 ;
        RECT 1368.565 1014.370 1368.895 1014.385 ;
        RECT 1367.645 1014.070 1368.895 1014.370 ;
        RECT 1367.645 1014.055 1367.975 1014.070 ;
        RECT 1368.565 1014.055 1368.895 1014.070 ;
        RECT 1367.645 917.810 1367.975 917.825 ;
        RECT 1368.565 917.810 1368.895 917.825 ;
        RECT 1367.645 917.510 1368.895 917.810 ;
        RECT 1367.645 917.495 1367.975 917.510 ;
        RECT 1368.565 917.495 1368.895 917.510 ;
        RECT 1367.645 628.810 1367.975 628.825 ;
        RECT 1367.430 628.495 1367.975 628.810 ;
        RECT 1367.430 628.145 1367.730 628.495 ;
        RECT 1367.430 627.830 1367.975 628.145 ;
        RECT 1367.645 627.815 1367.975 627.830 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 565.410 54.980 565.730 55.040 ;
        RECT 1380.070 54.980 1380.390 55.040 ;
        RECT 565.410 54.840 1380.390 54.980 ;
        RECT 565.410 54.780 565.730 54.840 ;
        RECT 1380.070 54.780 1380.390 54.840 ;
        RECT 561.730 14.860 562.050 14.920 ;
        RECT 565.410 14.860 565.730 14.920 ;
        RECT 561.730 14.720 565.730 14.860 ;
        RECT 561.730 14.660 562.050 14.720 ;
        RECT 565.410 14.660 565.730 14.720 ;
      LAYER via ;
        RECT 565.440 54.780 565.700 55.040 ;
        RECT 1380.100 54.780 1380.360 55.040 ;
        RECT 561.760 14.660 562.020 14.920 ;
        RECT 565.440 14.660 565.700 14.920 ;
      LAYER met2 ;
        RECT 1380.025 1700.000 1380.305 1704.000 ;
        RECT 1380.160 55.070 1380.300 1700.000 ;
        RECT 565.440 54.750 565.700 55.070 ;
        RECT 1380.100 54.750 1380.360 55.070 ;
        RECT 565.500 14.950 565.640 54.750 ;
        RECT 561.760 14.630 562.020 14.950 ;
        RECT 565.440 14.630 565.700 14.950 ;
        RECT 561.820 2.400 561.960 14.630 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 585.650 51.240 585.970 51.300 ;
        RECT 1387.890 51.240 1388.210 51.300 ;
        RECT 585.650 51.100 1388.210 51.240 ;
        RECT 585.650 51.040 585.970 51.100 ;
        RECT 1387.890 51.040 1388.210 51.100 ;
        RECT 579.670 14.860 579.990 14.920 ;
        RECT 584.730 14.860 585.050 14.920 ;
        RECT 579.670 14.720 585.050 14.860 ;
        RECT 579.670 14.660 579.990 14.720 ;
        RECT 584.730 14.660 585.050 14.720 ;
      LAYER via ;
        RECT 585.680 51.040 585.940 51.300 ;
        RECT 1387.920 51.040 1388.180 51.300 ;
        RECT 579.700 14.660 579.960 14.920 ;
        RECT 584.760 14.660 585.020 14.920 ;
      LAYER met2 ;
        RECT 1387.385 1700.410 1387.665 1704.000 ;
        RECT 1387.385 1700.270 1388.120 1700.410 ;
        RECT 1387.385 1700.000 1387.665 1700.270 ;
        RECT 1387.980 51.330 1388.120 1700.270 ;
        RECT 585.680 51.010 585.940 51.330 ;
        RECT 1387.920 51.010 1388.180 51.330 ;
        RECT 585.740 18.090 585.880 51.010 ;
        RECT 584.820 17.950 585.880 18.090 ;
        RECT 584.820 14.950 584.960 17.950 ;
        RECT 579.700 14.630 579.960 14.950 ;
        RECT 584.760 14.630 585.020 14.950 ;
        RECT 579.760 2.400 579.900 14.630 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1180.430 1678.140 1180.750 1678.200 ;
        RECT 1182.730 1678.140 1183.050 1678.200 ;
        RECT 1180.430 1678.000 1183.050 1678.140 ;
        RECT 1180.430 1677.940 1180.750 1678.000 ;
        RECT 1182.730 1677.940 1183.050 1678.000 ;
        RECT 86.090 25.740 86.410 25.800 ;
        RECT 1180.430 25.740 1180.750 25.800 ;
        RECT 86.090 25.600 1180.750 25.740 ;
        RECT 86.090 25.540 86.410 25.600 ;
        RECT 1180.430 25.540 1180.750 25.600 ;
      LAYER via ;
        RECT 1180.460 1677.940 1180.720 1678.200 ;
        RECT 1182.760 1677.940 1183.020 1678.200 ;
        RECT 86.120 25.540 86.380 25.800 ;
        RECT 1180.460 25.540 1180.720 25.800 ;
      LAYER met2 ;
        RECT 1184.065 1700.410 1184.345 1704.000 ;
        RECT 1182.820 1700.270 1184.345 1700.410 ;
        RECT 1182.820 1678.230 1182.960 1700.270 ;
        RECT 1184.065 1700.000 1184.345 1700.270 ;
        RECT 1180.460 1677.910 1180.720 1678.230 ;
        RECT 1182.760 1677.910 1183.020 1678.230 ;
        RECT 1180.520 25.830 1180.660 1677.910 ;
        RECT 86.120 25.510 86.380 25.830 ;
        RECT 1180.460 25.510 1180.720 25.830 ;
        RECT 86.180 2.400 86.320 25.510 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1394.330 1677.120 1394.650 1677.180 ;
        RECT 1394.330 1676.980 1395.020 1677.120 ;
        RECT 1394.330 1676.920 1394.650 1676.980 ;
        RECT 1394.880 1676.160 1395.020 1676.980 ;
        RECT 1394.790 1675.900 1395.110 1676.160 ;
        RECT 599.910 50.900 600.230 50.960 ;
        RECT 1394.790 50.900 1395.110 50.960 ;
        RECT 599.910 50.760 1395.110 50.900 ;
        RECT 599.910 50.700 600.230 50.760 ;
        RECT 1394.790 50.700 1395.110 50.760 ;
        RECT 597.150 14.860 597.470 14.920 ;
        RECT 599.910 14.860 600.230 14.920 ;
        RECT 597.150 14.720 600.230 14.860 ;
        RECT 597.150 14.660 597.470 14.720 ;
        RECT 599.910 14.660 600.230 14.720 ;
      LAYER via ;
        RECT 1394.360 1676.920 1394.620 1677.180 ;
        RECT 1394.820 1675.900 1395.080 1676.160 ;
        RECT 599.940 50.700 600.200 50.960 ;
        RECT 1394.820 50.700 1395.080 50.960 ;
        RECT 597.180 14.660 597.440 14.920 ;
        RECT 599.940 14.660 600.200 14.920 ;
      LAYER met2 ;
        RECT 1394.745 1700.410 1395.025 1704.000 ;
        RECT 1394.420 1700.270 1395.025 1700.410 ;
        RECT 1394.420 1677.210 1394.560 1700.270 ;
        RECT 1394.745 1700.000 1395.025 1700.270 ;
        RECT 1394.360 1676.890 1394.620 1677.210 ;
        RECT 1394.820 1675.870 1395.080 1676.190 ;
        RECT 1394.880 50.990 1395.020 1675.870 ;
        RECT 599.940 50.670 600.200 50.990 ;
        RECT 1394.820 50.670 1395.080 50.990 ;
        RECT 600.000 14.950 600.140 50.670 ;
        RECT 597.180 14.630 597.440 14.950 ;
        RECT 599.940 14.630 600.200 14.950 ;
        RECT 597.240 2.400 597.380 14.630 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 620.610 50.560 620.930 50.620 ;
        RECT 1401.690 50.560 1402.010 50.620 ;
        RECT 620.610 50.420 1402.010 50.560 ;
        RECT 620.610 50.360 620.930 50.420 ;
        RECT 1401.690 50.360 1402.010 50.420 ;
      LAYER via ;
        RECT 620.640 50.360 620.900 50.620 ;
        RECT 1401.720 50.360 1401.980 50.620 ;
      LAYER met2 ;
        RECT 1402.105 1700.410 1402.385 1704.000 ;
        RECT 1401.780 1700.270 1402.385 1700.410 ;
        RECT 1401.780 50.650 1401.920 1700.270 ;
        RECT 1402.105 1700.000 1402.385 1700.270 ;
        RECT 620.640 50.330 620.900 50.650 ;
        RECT 1401.720 50.330 1401.980 50.650 ;
        RECT 620.700 17.410 620.840 50.330 ;
        RECT 615.180 17.270 620.840 17.410 ;
        RECT 615.180 2.400 615.320 17.270 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 109.550 38.660 109.870 38.720 ;
        RECT 1194.230 38.660 1194.550 38.720 ;
        RECT 109.550 38.520 1194.550 38.660 ;
        RECT 109.550 38.460 109.870 38.520 ;
        RECT 1194.230 38.460 1194.550 38.520 ;
      LAYER via ;
        RECT 109.580 38.460 109.840 38.720 ;
        RECT 1194.260 38.460 1194.520 38.720 ;
      LAYER met2 ;
        RECT 1193.725 1700.410 1194.005 1704.000 ;
        RECT 1193.725 1700.270 1194.460 1700.410 ;
        RECT 1193.725 1700.000 1194.005 1700.270 ;
        RECT 1194.320 38.750 1194.460 1700.270 ;
        RECT 109.580 38.430 109.840 38.750 ;
        RECT 1194.260 38.430 1194.520 38.750 ;
        RECT 109.640 2.400 109.780 38.430 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 133.470 39.000 133.790 39.060 ;
        RECT 1202.050 39.000 1202.370 39.060 ;
        RECT 133.470 38.860 1202.370 39.000 ;
        RECT 133.470 38.800 133.790 38.860 ;
        RECT 1202.050 38.800 1202.370 38.860 ;
      LAYER via ;
        RECT 133.500 38.800 133.760 39.060 ;
        RECT 1202.080 38.800 1202.340 39.060 ;
      LAYER met2 ;
        RECT 1203.845 1700.410 1204.125 1704.000 ;
        RECT 1202.140 1700.270 1204.125 1700.410 ;
        RECT 1202.140 39.090 1202.280 1700.270 ;
        RECT 1203.845 1700.000 1204.125 1700.270 ;
        RECT 133.500 38.770 133.760 39.090 ;
        RECT 1202.080 38.770 1202.340 39.090 ;
        RECT 133.560 2.400 133.700 38.770 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 151.410 39.340 151.730 39.400 ;
        RECT 1208.950 39.340 1209.270 39.400 ;
        RECT 151.410 39.200 1209.270 39.340 ;
        RECT 151.410 39.140 151.730 39.200 ;
        RECT 1208.950 39.140 1209.270 39.200 ;
      LAYER via ;
        RECT 151.440 39.140 151.700 39.400 ;
        RECT 1208.980 39.140 1209.240 39.400 ;
      LAYER met2 ;
        RECT 1211.205 1700.410 1211.485 1704.000 ;
        RECT 1209.040 1700.270 1211.485 1700.410 ;
        RECT 1209.040 39.430 1209.180 1700.270 ;
        RECT 1211.205 1700.000 1211.485 1700.270 ;
        RECT 151.440 39.110 151.700 39.430 ;
        RECT 1208.980 39.110 1209.240 39.430 ;
        RECT 151.500 2.400 151.640 39.110 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1214.930 1660.460 1215.250 1660.520 ;
        RECT 1217.230 1660.460 1217.550 1660.520 ;
        RECT 1214.930 1660.320 1217.550 1660.460 ;
        RECT 1214.930 1660.260 1215.250 1660.320 ;
        RECT 1217.230 1660.260 1217.550 1660.320 ;
        RECT 169.350 39.680 169.670 39.740 ;
        RECT 1214.930 39.680 1215.250 39.740 ;
        RECT 169.350 39.540 1215.250 39.680 ;
        RECT 169.350 39.480 169.670 39.540 ;
        RECT 1214.930 39.480 1215.250 39.540 ;
      LAYER via ;
        RECT 1214.960 1660.260 1215.220 1660.520 ;
        RECT 1217.260 1660.260 1217.520 1660.520 ;
        RECT 169.380 39.480 169.640 39.740 ;
        RECT 1214.960 39.480 1215.220 39.740 ;
      LAYER met2 ;
        RECT 1218.565 1700.410 1218.845 1704.000 ;
        RECT 1217.320 1700.270 1218.845 1700.410 ;
        RECT 1217.320 1660.550 1217.460 1700.270 ;
        RECT 1218.565 1700.000 1218.845 1700.270 ;
        RECT 1214.960 1660.230 1215.220 1660.550 ;
        RECT 1217.260 1660.230 1217.520 1660.550 ;
        RECT 1215.020 39.770 1215.160 1660.230 ;
        RECT 169.380 39.450 169.640 39.770 ;
        RECT 1214.960 39.450 1215.220 39.770 ;
        RECT 169.440 2.400 169.580 39.450 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1221.905 1062.245 1222.075 1103.895 ;
        RECT 1221.905 517.565 1222.075 565.675 ;
        RECT 1221.905 282.965 1222.075 331.075 ;
        RECT 1220.985 83.045 1221.155 110.755 ;
      LAYER mcon ;
        RECT 1221.905 1103.725 1222.075 1103.895 ;
        RECT 1221.905 565.505 1222.075 565.675 ;
        RECT 1221.905 330.905 1222.075 331.075 ;
        RECT 1220.985 110.585 1221.155 110.755 ;
      LAYER met1 ;
        RECT 1221.830 1559.620 1222.150 1559.880 ;
        RECT 1221.920 1558.800 1222.060 1559.620 ;
        RECT 1222.290 1558.800 1222.610 1558.860 ;
        RECT 1221.920 1558.660 1222.610 1558.800 ;
        RECT 1222.290 1558.600 1222.610 1558.660 ;
        RECT 1222.290 1442.180 1222.610 1442.240 ;
        RECT 1222.750 1442.180 1223.070 1442.240 ;
        RECT 1222.290 1442.040 1223.070 1442.180 ;
        RECT 1222.290 1441.980 1222.610 1442.040 ;
        RECT 1222.750 1441.980 1223.070 1442.040 ;
        RECT 1221.830 1297.340 1222.150 1297.400 ;
        RECT 1222.290 1297.340 1222.610 1297.400 ;
        RECT 1221.830 1297.200 1222.610 1297.340 ;
        RECT 1221.830 1297.140 1222.150 1297.200 ;
        RECT 1222.290 1297.140 1222.610 1297.200 ;
        RECT 1221.830 1200.780 1222.150 1200.840 ;
        RECT 1222.750 1200.780 1223.070 1200.840 ;
        RECT 1221.830 1200.640 1223.070 1200.780 ;
        RECT 1221.830 1200.580 1222.150 1200.640 ;
        RECT 1222.750 1200.580 1223.070 1200.640 ;
        RECT 1222.290 1173.240 1222.610 1173.300 ;
        RECT 1221.920 1173.100 1222.610 1173.240 ;
        RECT 1221.920 1172.960 1222.060 1173.100 ;
        RECT 1222.290 1173.040 1222.610 1173.100 ;
        RECT 1221.830 1172.700 1222.150 1172.960 ;
        RECT 1221.830 1103.880 1222.150 1103.940 ;
        RECT 1221.635 1103.740 1222.150 1103.880 ;
        RECT 1221.830 1103.680 1222.150 1103.740 ;
        RECT 1221.845 1062.400 1222.135 1062.445 ;
        RECT 1222.290 1062.400 1222.610 1062.460 ;
        RECT 1221.845 1062.260 1222.610 1062.400 ;
        RECT 1221.845 1062.215 1222.135 1062.260 ;
        RECT 1222.290 1062.200 1222.610 1062.260 ;
        RECT 1221.830 1014.460 1222.150 1014.520 ;
        RECT 1222.750 1014.460 1223.070 1014.520 ;
        RECT 1221.830 1014.320 1223.070 1014.460 ;
        RECT 1221.830 1014.260 1222.150 1014.320 ;
        RECT 1222.750 1014.260 1223.070 1014.320 ;
        RECT 1221.830 966.180 1222.150 966.240 ;
        RECT 1222.290 966.180 1222.610 966.240 ;
        RECT 1221.830 966.040 1222.610 966.180 ;
        RECT 1221.830 965.980 1222.150 966.040 ;
        RECT 1222.290 965.980 1222.610 966.040 ;
        RECT 1221.830 855.140 1222.150 855.400 ;
        RECT 1221.920 855.000 1222.060 855.140 ;
        RECT 1222.750 855.000 1223.070 855.060 ;
        RECT 1221.920 854.860 1223.070 855.000 ;
        RECT 1222.750 854.800 1223.070 854.860 ;
        RECT 1221.830 690.240 1222.150 690.500 ;
        RECT 1221.920 689.820 1222.060 690.240 ;
        RECT 1221.830 689.560 1222.150 689.820 ;
        RECT 1221.370 572.800 1221.690 572.860 ;
        RECT 1222.290 572.800 1222.610 572.860 ;
        RECT 1221.370 572.660 1222.610 572.800 ;
        RECT 1221.370 572.600 1221.690 572.660 ;
        RECT 1222.290 572.600 1222.610 572.660 ;
        RECT 1221.370 565.660 1221.690 565.720 ;
        RECT 1221.845 565.660 1222.135 565.705 ;
        RECT 1221.370 565.520 1222.135 565.660 ;
        RECT 1221.370 565.460 1221.690 565.520 ;
        RECT 1221.845 565.475 1222.135 565.520 ;
        RECT 1221.830 517.720 1222.150 517.780 ;
        RECT 1221.635 517.580 1222.150 517.720 ;
        RECT 1221.830 517.520 1222.150 517.580 ;
        RECT 1221.830 517.040 1222.150 517.100 ;
        RECT 1222.750 517.040 1223.070 517.100 ;
        RECT 1221.830 516.900 1223.070 517.040 ;
        RECT 1221.830 516.840 1222.150 516.900 ;
        RECT 1222.750 516.840 1223.070 516.900 ;
        RECT 1221.830 331.060 1222.150 331.120 ;
        RECT 1221.635 330.920 1222.150 331.060 ;
        RECT 1221.830 330.860 1222.150 330.920 ;
        RECT 1221.845 283.120 1222.135 283.165 ;
        RECT 1222.290 283.120 1222.610 283.180 ;
        RECT 1221.845 282.980 1222.610 283.120 ;
        RECT 1221.845 282.935 1222.135 282.980 ;
        RECT 1222.290 282.920 1222.610 282.980 ;
        RECT 1221.830 241.640 1222.150 241.700 ;
        RECT 1222.750 241.640 1223.070 241.700 ;
        RECT 1221.830 241.500 1223.070 241.640 ;
        RECT 1221.830 241.440 1222.150 241.500 ;
        RECT 1222.750 241.440 1223.070 241.500 ;
        RECT 1221.830 193.500 1222.150 193.760 ;
        RECT 1221.920 193.360 1222.060 193.500 ;
        RECT 1222.290 193.360 1222.610 193.420 ;
        RECT 1221.920 193.220 1222.610 193.360 ;
        RECT 1222.290 193.160 1222.610 193.220 ;
        RECT 1220.925 110.740 1221.215 110.785 ;
        RECT 1222.290 110.740 1222.610 110.800 ;
        RECT 1220.925 110.600 1222.610 110.740 ;
        RECT 1220.925 110.555 1221.215 110.600 ;
        RECT 1222.290 110.540 1222.610 110.600 ;
        RECT 1220.910 83.200 1221.230 83.260 ;
        RECT 1220.715 83.060 1221.230 83.200 ;
        RECT 1220.910 83.000 1221.230 83.060 ;
        RECT 186.830 40.020 187.150 40.080 ;
        RECT 1221.370 40.020 1221.690 40.080 ;
        RECT 186.830 39.880 1221.690 40.020 ;
        RECT 186.830 39.820 187.150 39.880 ;
        RECT 1221.370 39.820 1221.690 39.880 ;
      LAYER via ;
        RECT 1221.860 1559.620 1222.120 1559.880 ;
        RECT 1222.320 1558.600 1222.580 1558.860 ;
        RECT 1222.320 1441.980 1222.580 1442.240 ;
        RECT 1222.780 1441.980 1223.040 1442.240 ;
        RECT 1221.860 1297.140 1222.120 1297.400 ;
        RECT 1222.320 1297.140 1222.580 1297.400 ;
        RECT 1221.860 1200.580 1222.120 1200.840 ;
        RECT 1222.780 1200.580 1223.040 1200.840 ;
        RECT 1222.320 1173.040 1222.580 1173.300 ;
        RECT 1221.860 1172.700 1222.120 1172.960 ;
        RECT 1221.860 1103.680 1222.120 1103.940 ;
        RECT 1222.320 1062.200 1222.580 1062.460 ;
        RECT 1221.860 1014.260 1222.120 1014.520 ;
        RECT 1222.780 1014.260 1223.040 1014.520 ;
        RECT 1221.860 965.980 1222.120 966.240 ;
        RECT 1222.320 965.980 1222.580 966.240 ;
        RECT 1221.860 855.140 1222.120 855.400 ;
        RECT 1222.780 854.800 1223.040 855.060 ;
        RECT 1221.860 690.240 1222.120 690.500 ;
        RECT 1221.860 689.560 1222.120 689.820 ;
        RECT 1221.400 572.600 1221.660 572.860 ;
        RECT 1222.320 572.600 1222.580 572.860 ;
        RECT 1221.400 565.460 1221.660 565.720 ;
        RECT 1221.860 517.520 1222.120 517.780 ;
        RECT 1221.860 516.840 1222.120 517.100 ;
        RECT 1222.780 516.840 1223.040 517.100 ;
        RECT 1221.860 330.860 1222.120 331.120 ;
        RECT 1222.320 282.920 1222.580 283.180 ;
        RECT 1221.860 241.440 1222.120 241.700 ;
        RECT 1222.780 241.440 1223.040 241.700 ;
        RECT 1221.860 193.500 1222.120 193.760 ;
        RECT 1222.320 193.160 1222.580 193.420 ;
        RECT 1222.320 110.540 1222.580 110.800 ;
        RECT 1220.940 83.000 1221.200 83.260 ;
        RECT 186.860 39.820 187.120 40.080 ;
        RECT 1221.400 39.820 1221.660 40.080 ;
      LAYER met2 ;
        RECT 1225.925 1701.090 1226.205 1704.000 ;
        RECT 1223.760 1700.950 1226.205 1701.090 ;
        RECT 1223.760 1656.210 1223.900 1700.950 ;
        RECT 1225.925 1700.000 1226.205 1700.950 ;
        RECT 1222.380 1656.070 1223.900 1656.210 ;
        RECT 1222.380 1587.530 1222.520 1656.070 ;
        RECT 1221.920 1587.390 1222.520 1587.530 ;
        RECT 1221.920 1559.910 1222.060 1587.390 ;
        RECT 1221.860 1559.590 1222.120 1559.910 ;
        RECT 1222.320 1558.570 1222.580 1558.890 ;
        RECT 1222.380 1442.270 1222.520 1558.570 ;
        RECT 1222.320 1441.950 1222.580 1442.270 ;
        RECT 1222.780 1441.950 1223.040 1442.270 ;
        RECT 1222.840 1352.760 1222.980 1441.950 ;
        RECT 1222.380 1352.620 1222.980 1352.760 ;
        RECT 1222.380 1297.430 1222.520 1352.620 ;
        RECT 1221.860 1297.110 1222.120 1297.430 ;
        RECT 1222.320 1297.110 1222.580 1297.430 ;
        RECT 1221.920 1249.005 1222.060 1297.110 ;
        RECT 1221.850 1248.635 1222.130 1249.005 ;
        RECT 1222.770 1248.635 1223.050 1249.005 ;
        RECT 1221.920 1200.870 1222.060 1201.025 ;
        RECT 1222.840 1200.870 1222.980 1248.635 ;
        RECT 1221.860 1200.610 1222.120 1200.870 ;
        RECT 1221.860 1200.550 1222.520 1200.610 ;
        RECT 1222.780 1200.550 1223.040 1200.870 ;
        RECT 1221.920 1200.470 1222.520 1200.550 ;
        RECT 1222.380 1173.330 1222.520 1200.470 ;
        RECT 1222.320 1173.010 1222.580 1173.330 ;
        RECT 1221.860 1172.670 1222.120 1172.990 ;
        RECT 1221.920 1103.970 1222.060 1172.670 ;
        RECT 1221.860 1103.650 1222.120 1103.970 ;
        RECT 1222.320 1062.170 1222.580 1062.490 ;
        RECT 1222.380 1055.770 1222.520 1062.170 ;
        RECT 1222.380 1055.630 1222.980 1055.770 ;
        RECT 1222.840 1014.550 1222.980 1055.630 ;
        RECT 1221.860 1014.230 1222.120 1014.550 ;
        RECT 1222.780 1014.230 1223.040 1014.550 ;
        RECT 1221.920 966.270 1222.060 1014.230 ;
        RECT 1221.860 965.950 1222.120 966.270 ;
        RECT 1222.320 965.950 1222.580 966.270 ;
        RECT 1222.380 927.930 1222.520 965.950 ;
        RECT 1222.380 927.790 1222.980 927.930 ;
        RECT 1222.840 910.250 1222.980 927.790 ;
        RECT 1221.920 910.110 1222.980 910.250 ;
        RECT 1221.920 855.430 1222.060 910.110 ;
        RECT 1221.860 855.110 1222.120 855.430 ;
        RECT 1222.780 854.770 1223.040 855.090 ;
        RECT 1222.840 724.725 1222.980 854.770 ;
        RECT 1221.850 724.355 1222.130 724.725 ;
        RECT 1222.770 724.355 1223.050 724.725 ;
        RECT 1221.920 690.530 1222.060 724.355 ;
        RECT 1221.860 690.210 1222.120 690.530 ;
        RECT 1221.860 689.530 1222.120 689.850 ;
        RECT 1221.920 651.850 1222.060 689.530 ;
        RECT 1221.920 651.710 1222.520 651.850 ;
        RECT 1222.380 572.890 1222.520 651.710 ;
        RECT 1221.400 572.570 1221.660 572.890 ;
        RECT 1222.320 572.570 1222.580 572.890 ;
        RECT 1221.460 565.750 1221.600 572.570 ;
        RECT 1221.400 565.430 1221.660 565.750 ;
        RECT 1221.860 517.490 1222.120 517.810 ;
        RECT 1221.920 517.130 1222.060 517.490 ;
        RECT 1221.860 516.810 1222.120 517.130 ;
        RECT 1222.780 516.810 1223.040 517.130 ;
        RECT 1222.840 482.530 1222.980 516.810 ;
        RECT 1222.380 482.390 1222.980 482.530 ;
        RECT 1222.380 356.050 1222.520 482.390 ;
        RECT 1222.380 355.910 1222.980 356.050 ;
        RECT 1222.840 332.365 1222.980 355.910 ;
        RECT 1222.770 331.995 1223.050 332.365 ;
        RECT 1221.850 331.315 1222.130 331.685 ;
        RECT 1221.920 331.150 1222.060 331.315 ;
        RECT 1221.860 330.830 1222.120 331.150 ;
        RECT 1222.320 282.890 1222.580 283.210 ;
        RECT 1222.380 266.290 1222.520 282.890 ;
        RECT 1222.380 266.150 1222.980 266.290 ;
        RECT 1222.840 241.730 1222.980 266.150 ;
        RECT 1221.860 241.410 1222.120 241.730 ;
        RECT 1222.780 241.410 1223.040 241.730 ;
        RECT 1221.920 193.790 1222.060 241.410 ;
        RECT 1221.860 193.470 1222.120 193.790 ;
        RECT 1222.320 193.130 1222.580 193.450 ;
        RECT 1222.380 110.830 1222.520 193.130 ;
        RECT 1222.320 110.510 1222.580 110.830 ;
        RECT 1220.940 82.970 1221.200 83.290 ;
        RECT 1221.000 55.490 1221.140 82.970 ;
        RECT 1221.000 55.350 1221.600 55.490 ;
        RECT 1221.460 40.110 1221.600 55.350 ;
        RECT 186.860 39.790 187.120 40.110 ;
        RECT 1221.400 39.790 1221.660 40.110 ;
        RECT 186.920 2.400 187.060 39.790 ;
        RECT 186.710 -4.800 187.270 2.400 ;
      LAYER via2 ;
        RECT 1221.850 1248.680 1222.130 1248.960 ;
        RECT 1222.770 1248.680 1223.050 1248.960 ;
        RECT 1221.850 724.400 1222.130 724.680 ;
        RECT 1222.770 724.400 1223.050 724.680 ;
        RECT 1222.770 332.040 1223.050 332.320 ;
        RECT 1221.850 331.360 1222.130 331.640 ;
      LAYER met3 ;
        RECT 1221.825 1248.970 1222.155 1248.985 ;
        RECT 1222.745 1248.970 1223.075 1248.985 ;
        RECT 1221.825 1248.670 1223.075 1248.970 ;
        RECT 1221.825 1248.655 1222.155 1248.670 ;
        RECT 1222.745 1248.655 1223.075 1248.670 ;
        RECT 1221.825 724.690 1222.155 724.705 ;
        RECT 1222.745 724.690 1223.075 724.705 ;
        RECT 1221.825 724.390 1223.075 724.690 ;
        RECT 1221.825 724.375 1222.155 724.390 ;
        RECT 1222.745 724.375 1223.075 724.390 ;
        RECT 1222.745 332.330 1223.075 332.345 ;
        RECT 1221.150 332.030 1223.075 332.330 ;
        RECT 1221.150 331.650 1221.450 332.030 ;
        RECT 1222.745 332.015 1223.075 332.030 ;
        RECT 1221.825 331.650 1222.155 331.665 ;
        RECT 1221.150 331.350 1222.155 331.650 ;
        RECT 1221.825 331.335 1222.155 331.350 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1229.265 945.285 1229.435 959.395 ;
        RECT 1229.265 689.605 1229.435 717.655 ;
        RECT 1229.725 572.645 1229.895 579.955 ;
        RECT 1229.725 483.225 1229.895 531.335 ;
        RECT 1229.265 83.045 1229.435 131.155 ;
      LAYER mcon ;
        RECT 1229.265 959.225 1229.435 959.395 ;
        RECT 1229.265 717.485 1229.435 717.655 ;
        RECT 1229.725 579.785 1229.895 579.955 ;
        RECT 1229.725 531.165 1229.895 531.335 ;
        RECT 1229.265 130.985 1229.435 131.155 ;
      LAYER met1 ;
        RECT 1229.190 1559.620 1229.510 1559.880 ;
        RECT 1229.280 1558.800 1229.420 1559.620 ;
        RECT 1229.650 1558.800 1229.970 1558.860 ;
        RECT 1229.280 1558.660 1229.970 1558.800 ;
        RECT 1229.650 1558.600 1229.970 1558.660 ;
        RECT 1229.650 1345.620 1229.970 1345.680 ;
        RECT 1230.570 1345.620 1230.890 1345.680 ;
        RECT 1229.650 1345.480 1230.890 1345.620 ;
        RECT 1229.650 1345.420 1229.970 1345.480 ;
        RECT 1230.570 1345.420 1230.890 1345.480 ;
        RECT 1229.190 1249.060 1229.510 1249.120 ;
        RECT 1230.110 1249.060 1230.430 1249.120 ;
        RECT 1229.190 1248.920 1230.430 1249.060 ;
        RECT 1229.190 1248.860 1229.510 1248.920 ;
        RECT 1230.110 1248.860 1230.430 1248.920 ;
        RECT 1229.650 1200.780 1229.970 1200.840 ;
        RECT 1230.570 1200.780 1230.890 1200.840 ;
        RECT 1229.650 1200.640 1230.890 1200.780 ;
        RECT 1229.650 1200.580 1229.970 1200.640 ;
        RECT 1230.570 1200.580 1230.890 1200.640 ;
        RECT 1229.190 1104.220 1229.510 1104.280 ;
        RECT 1230.110 1104.220 1230.430 1104.280 ;
        RECT 1229.190 1104.080 1230.430 1104.220 ;
        RECT 1229.190 1104.020 1229.510 1104.080 ;
        RECT 1230.110 1104.020 1230.430 1104.080 ;
        RECT 1229.190 1062.740 1229.510 1062.800 ;
        RECT 1229.650 1062.740 1229.970 1062.800 ;
        RECT 1229.190 1062.600 1229.970 1062.740 ;
        RECT 1229.190 1062.540 1229.510 1062.600 ;
        RECT 1229.650 1062.540 1229.970 1062.600 ;
        RECT 1229.190 1014.460 1229.510 1014.520 ;
        RECT 1229.650 1014.460 1229.970 1014.520 ;
        RECT 1229.190 1014.320 1229.970 1014.460 ;
        RECT 1229.190 1014.260 1229.510 1014.320 ;
        RECT 1229.650 1014.260 1229.970 1014.320 ;
        RECT 1229.190 959.380 1229.510 959.440 ;
        RECT 1228.995 959.240 1229.510 959.380 ;
        RECT 1229.190 959.180 1229.510 959.240 ;
        RECT 1226.890 945.440 1227.210 945.500 ;
        RECT 1229.205 945.440 1229.495 945.485 ;
        RECT 1226.890 945.300 1229.495 945.440 ;
        RECT 1226.890 945.240 1227.210 945.300 ;
        RECT 1229.205 945.255 1229.495 945.300 ;
        RECT 1226.890 903.280 1227.210 903.340 ;
        RECT 1229.190 903.280 1229.510 903.340 ;
        RECT 1226.890 903.140 1229.510 903.280 ;
        RECT 1226.890 903.080 1227.210 903.140 ;
        RECT 1229.190 903.080 1229.510 903.140 ;
        RECT 1229.190 782.920 1229.510 782.980 ;
        RECT 1230.110 782.920 1230.430 782.980 ;
        RECT 1229.190 782.780 1230.430 782.920 ;
        RECT 1229.190 782.720 1229.510 782.780 ;
        RECT 1230.110 782.720 1230.430 782.780 ;
        RECT 1229.190 717.640 1229.510 717.700 ;
        RECT 1228.995 717.500 1229.510 717.640 ;
        RECT 1229.190 717.440 1229.510 717.500 ;
        RECT 1229.190 689.760 1229.510 689.820 ;
        RECT 1228.995 689.620 1229.510 689.760 ;
        RECT 1229.190 689.560 1229.510 689.620 ;
        RECT 1229.650 579.940 1229.970 580.000 ;
        RECT 1229.455 579.800 1229.970 579.940 ;
        RECT 1229.650 579.740 1229.970 579.800 ;
        RECT 1229.650 572.800 1229.970 572.860 ;
        RECT 1229.455 572.660 1229.970 572.800 ;
        RECT 1229.650 572.600 1229.970 572.660 ;
        RECT 1229.650 531.320 1229.970 531.380 ;
        RECT 1229.455 531.180 1229.970 531.320 ;
        RECT 1229.650 531.120 1229.970 531.180 ;
        RECT 1229.650 483.380 1229.970 483.440 ;
        RECT 1229.455 483.240 1229.970 483.380 ;
        RECT 1229.650 483.180 1229.970 483.240 ;
        RECT 1229.650 338.340 1229.970 338.600 ;
        RECT 1229.740 337.580 1229.880 338.340 ;
        RECT 1229.650 337.320 1229.970 337.580 ;
        RECT 1229.650 331.060 1229.970 331.120 ;
        RECT 1229.650 330.920 1230.340 331.060 ;
        RECT 1229.650 330.860 1229.970 330.920 ;
        RECT 1230.200 330.780 1230.340 330.920 ;
        RECT 1230.110 330.520 1230.430 330.780 ;
        RECT 1227.810 201.860 1228.130 201.920 ;
        RECT 1229.650 201.860 1229.970 201.920 ;
        RECT 1227.810 201.720 1229.970 201.860 ;
        RECT 1227.810 201.660 1228.130 201.720 ;
        RECT 1229.650 201.660 1229.970 201.720 ;
        RECT 1229.205 131.140 1229.495 131.185 ;
        RECT 1229.650 131.140 1229.970 131.200 ;
        RECT 1229.205 131.000 1229.970 131.140 ;
        RECT 1229.205 130.955 1229.495 131.000 ;
        RECT 1229.650 130.940 1229.970 131.000 ;
        RECT 1229.190 83.200 1229.510 83.260 ;
        RECT 1228.995 83.060 1229.510 83.200 ;
        RECT 1229.190 83.000 1229.510 83.060 ;
        RECT 204.770 40.360 205.090 40.420 ;
        RECT 1229.650 40.360 1229.970 40.420 ;
        RECT 204.770 40.220 1229.970 40.360 ;
        RECT 204.770 40.160 205.090 40.220 ;
        RECT 1229.650 40.160 1229.970 40.220 ;
      LAYER via ;
        RECT 1229.220 1559.620 1229.480 1559.880 ;
        RECT 1229.680 1558.600 1229.940 1558.860 ;
        RECT 1229.680 1345.420 1229.940 1345.680 ;
        RECT 1230.600 1345.420 1230.860 1345.680 ;
        RECT 1229.220 1248.860 1229.480 1249.120 ;
        RECT 1230.140 1248.860 1230.400 1249.120 ;
        RECT 1229.680 1200.580 1229.940 1200.840 ;
        RECT 1230.600 1200.580 1230.860 1200.840 ;
        RECT 1229.220 1104.020 1229.480 1104.280 ;
        RECT 1230.140 1104.020 1230.400 1104.280 ;
        RECT 1229.220 1062.540 1229.480 1062.800 ;
        RECT 1229.680 1062.540 1229.940 1062.800 ;
        RECT 1229.220 1014.260 1229.480 1014.520 ;
        RECT 1229.680 1014.260 1229.940 1014.520 ;
        RECT 1229.220 959.180 1229.480 959.440 ;
        RECT 1226.920 945.240 1227.180 945.500 ;
        RECT 1226.920 903.080 1227.180 903.340 ;
        RECT 1229.220 903.080 1229.480 903.340 ;
        RECT 1229.220 782.720 1229.480 782.980 ;
        RECT 1230.140 782.720 1230.400 782.980 ;
        RECT 1229.220 717.440 1229.480 717.700 ;
        RECT 1229.220 689.560 1229.480 689.820 ;
        RECT 1229.680 579.740 1229.940 580.000 ;
        RECT 1229.680 572.600 1229.940 572.860 ;
        RECT 1229.680 531.120 1229.940 531.380 ;
        RECT 1229.680 483.180 1229.940 483.440 ;
        RECT 1229.680 338.340 1229.940 338.600 ;
        RECT 1229.680 337.320 1229.940 337.580 ;
        RECT 1229.680 330.860 1229.940 331.120 ;
        RECT 1230.140 330.520 1230.400 330.780 ;
        RECT 1227.840 201.660 1228.100 201.920 ;
        RECT 1229.680 201.660 1229.940 201.920 ;
        RECT 1229.680 130.940 1229.940 131.200 ;
        RECT 1229.220 83.000 1229.480 83.260 ;
        RECT 204.800 40.160 205.060 40.420 ;
        RECT 1229.680 40.160 1229.940 40.420 ;
      LAYER met2 ;
        RECT 1233.285 1701.090 1233.565 1704.000 ;
        RECT 1231.120 1700.950 1233.565 1701.090 ;
        RECT 1231.120 1673.210 1231.260 1700.950 ;
        RECT 1233.285 1700.000 1233.565 1700.950 ;
        RECT 1229.740 1673.070 1231.260 1673.210 ;
        RECT 1229.740 1587.530 1229.880 1673.070 ;
        RECT 1229.280 1587.390 1229.880 1587.530 ;
        RECT 1229.280 1559.910 1229.420 1587.390 ;
        RECT 1229.220 1559.590 1229.480 1559.910 ;
        RECT 1229.680 1558.570 1229.940 1558.890 ;
        RECT 1229.740 1393.845 1229.880 1558.570 ;
        RECT 1229.670 1393.475 1229.950 1393.845 ;
        RECT 1230.590 1393.475 1230.870 1393.845 ;
        RECT 1230.660 1345.710 1230.800 1393.475 ;
        RECT 1229.680 1345.390 1229.940 1345.710 ;
        RECT 1230.600 1345.390 1230.860 1345.710 ;
        RECT 1229.740 1328.450 1229.880 1345.390 ;
        RECT 1229.740 1328.310 1230.340 1328.450 ;
        RECT 1230.200 1317.570 1230.340 1328.310 ;
        RECT 1229.280 1317.430 1230.340 1317.570 ;
        RECT 1229.280 1297.285 1229.420 1317.430 ;
        RECT 1229.210 1296.915 1229.490 1297.285 ;
        RECT 1230.130 1296.915 1230.410 1297.285 ;
        RECT 1230.200 1249.150 1230.340 1296.915 ;
        RECT 1229.220 1249.005 1229.480 1249.150 ;
        RECT 1229.210 1248.635 1229.490 1249.005 ;
        RECT 1230.140 1248.830 1230.400 1249.150 ;
        RECT 1230.590 1248.635 1230.870 1249.005 ;
        RECT 1230.660 1200.870 1230.800 1248.635 ;
        RECT 1229.680 1200.550 1229.940 1200.870 ;
        RECT 1230.600 1200.550 1230.860 1200.870 ;
        RECT 1229.740 1136.690 1229.880 1200.550 ;
        RECT 1229.740 1136.550 1230.340 1136.690 ;
        RECT 1230.200 1104.310 1230.340 1136.550 ;
        RECT 1229.220 1103.990 1229.480 1104.310 ;
        RECT 1230.140 1103.990 1230.400 1104.310 ;
        RECT 1229.280 1062.830 1229.420 1103.990 ;
        RECT 1229.220 1062.510 1229.480 1062.830 ;
        RECT 1229.680 1062.510 1229.940 1062.830 ;
        RECT 1229.740 1014.550 1229.880 1062.510 ;
        RECT 1229.220 1014.230 1229.480 1014.550 ;
        RECT 1229.680 1014.230 1229.940 1014.550 ;
        RECT 1229.280 959.470 1229.420 1014.230 ;
        RECT 1229.220 959.150 1229.480 959.470 ;
        RECT 1226.920 945.210 1227.180 945.530 ;
        RECT 1226.980 903.370 1227.120 945.210 ;
        RECT 1226.920 903.050 1227.180 903.370 ;
        RECT 1229.220 903.050 1229.480 903.370 ;
        RECT 1229.280 783.010 1229.420 903.050 ;
        RECT 1229.220 782.690 1229.480 783.010 ;
        RECT 1230.140 782.690 1230.400 783.010 ;
        RECT 1230.200 717.925 1230.340 782.690 ;
        RECT 1229.210 717.555 1229.490 717.925 ;
        RECT 1230.130 717.555 1230.410 717.925 ;
        RECT 1229.220 717.410 1229.480 717.555 ;
        RECT 1229.220 689.530 1229.480 689.850 ;
        RECT 1229.280 651.850 1229.420 689.530 ;
        RECT 1229.280 651.710 1229.880 651.850 ;
        RECT 1229.740 580.030 1229.880 651.710 ;
        RECT 1229.680 579.710 1229.940 580.030 ;
        RECT 1229.680 572.570 1229.940 572.890 ;
        RECT 1229.740 531.410 1229.880 572.570 ;
        RECT 1229.680 531.090 1229.940 531.410 ;
        RECT 1229.680 483.150 1229.940 483.470 ;
        RECT 1229.740 338.630 1229.880 483.150 ;
        RECT 1229.680 338.310 1229.940 338.630 ;
        RECT 1229.680 337.290 1229.940 337.610 ;
        RECT 1229.740 331.150 1229.880 337.290 ;
        RECT 1229.680 330.830 1229.940 331.150 ;
        RECT 1230.140 330.490 1230.400 330.810 ;
        RECT 1230.200 303.010 1230.340 330.490 ;
        RECT 1229.740 302.870 1230.340 303.010 ;
        RECT 1229.740 241.925 1229.880 302.870 ;
        RECT 1229.670 241.555 1229.950 241.925 ;
        RECT 1227.830 240.875 1228.110 241.245 ;
        RECT 1227.900 201.950 1228.040 240.875 ;
        RECT 1227.840 201.630 1228.100 201.950 ;
        RECT 1229.680 201.630 1229.940 201.950 ;
        RECT 1229.740 131.230 1229.880 201.630 ;
        RECT 1229.680 130.910 1229.940 131.230 ;
        RECT 1229.220 82.970 1229.480 83.290 ;
        RECT 1229.280 65.690 1229.420 82.970 ;
        RECT 1229.280 65.550 1229.880 65.690 ;
        RECT 1229.740 40.450 1229.880 65.550 ;
        RECT 204.800 40.130 205.060 40.450 ;
        RECT 1229.680 40.130 1229.940 40.450 ;
        RECT 204.860 2.400 205.000 40.130 ;
        RECT 204.650 -4.800 205.210 2.400 ;
      LAYER via2 ;
        RECT 1229.670 1393.520 1229.950 1393.800 ;
        RECT 1230.590 1393.520 1230.870 1393.800 ;
        RECT 1229.210 1296.960 1229.490 1297.240 ;
        RECT 1230.130 1296.960 1230.410 1297.240 ;
        RECT 1229.210 1248.680 1229.490 1248.960 ;
        RECT 1230.590 1248.680 1230.870 1248.960 ;
        RECT 1229.210 717.600 1229.490 717.880 ;
        RECT 1230.130 717.600 1230.410 717.880 ;
        RECT 1229.670 241.600 1229.950 241.880 ;
        RECT 1227.830 240.920 1228.110 241.200 ;
      LAYER met3 ;
        RECT 1229.645 1393.810 1229.975 1393.825 ;
        RECT 1230.565 1393.810 1230.895 1393.825 ;
        RECT 1229.645 1393.510 1230.895 1393.810 ;
        RECT 1229.645 1393.495 1229.975 1393.510 ;
        RECT 1230.565 1393.495 1230.895 1393.510 ;
        RECT 1229.185 1297.250 1229.515 1297.265 ;
        RECT 1230.105 1297.250 1230.435 1297.265 ;
        RECT 1229.185 1296.950 1230.435 1297.250 ;
        RECT 1229.185 1296.935 1229.515 1296.950 ;
        RECT 1230.105 1296.935 1230.435 1296.950 ;
        RECT 1229.185 1248.970 1229.515 1248.985 ;
        RECT 1230.565 1248.970 1230.895 1248.985 ;
        RECT 1229.185 1248.670 1230.895 1248.970 ;
        RECT 1229.185 1248.655 1229.515 1248.670 ;
        RECT 1230.565 1248.655 1230.895 1248.670 ;
        RECT 1229.185 717.890 1229.515 717.905 ;
        RECT 1230.105 717.890 1230.435 717.905 ;
        RECT 1229.185 717.590 1230.435 717.890 ;
        RECT 1229.185 717.575 1229.515 717.590 ;
        RECT 1230.105 717.575 1230.435 717.590 ;
        RECT 1229.645 241.890 1229.975 241.905 ;
        RECT 1228.510 241.590 1229.975 241.890 ;
        RECT 1227.805 241.210 1228.135 241.225 ;
        RECT 1228.510 241.210 1228.810 241.590 ;
        RECT 1229.645 241.575 1229.975 241.590 ;
        RECT 1227.805 240.910 1228.810 241.210 ;
        RECT 1227.805 240.895 1228.135 240.910 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1236.165 1297.865 1236.335 1304.495 ;
        RECT 1236.165 1248.565 1236.335 1290.215 ;
        RECT 1235.705 807.245 1235.875 855.355 ;
        RECT 1236.625 572.645 1236.795 620.755 ;
        RECT 1235.705 469.285 1235.875 517.395 ;
        RECT 1235.705 365.925 1235.875 400.435 ;
        RECT 1236.165 227.885 1236.335 275.995 ;
        RECT 1236.165 131.665 1236.335 179.435 ;
        RECT 1235.705 45.645 1235.875 131.155 ;
      LAYER mcon ;
        RECT 1236.165 1304.325 1236.335 1304.495 ;
        RECT 1236.165 1290.045 1236.335 1290.215 ;
        RECT 1235.705 855.185 1235.875 855.355 ;
        RECT 1236.625 620.585 1236.795 620.755 ;
        RECT 1235.705 517.225 1235.875 517.395 ;
        RECT 1235.705 400.265 1235.875 400.435 ;
        RECT 1236.165 275.825 1236.335 275.995 ;
        RECT 1236.165 179.265 1236.335 179.435 ;
        RECT 1235.705 130.985 1235.875 131.155 ;
      LAYER met1 ;
        RECT 1235.170 1490.800 1235.490 1490.860 ;
        RECT 1236.550 1490.800 1236.870 1490.860 ;
        RECT 1235.170 1490.660 1236.870 1490.800 ;
        RECT 1235.170 1490.600 1235.490 1490.660 ;
        RECT 1236.550 1490.600 1236.870 1490.660 ;
        RECT 1235.170 1449.320 1235.490 1449.380 ;
        RECT 1236.090 1449.320 1236.410 1449.380 ;
        RECT 1235.170 1449.180 1236.410 1449.320 ;
        RECT 1235.170 1449.120 1235.490 1449.180 ;
        RECT 1236.090 1449.120 1236.410 1449.180 ;
        RECT 1235.170 1352.760 1235.490 1352.820 ;
        RECT 1236.090 1352.760 1236.410 1352.820 ;
        RECT 1235.170 1352.620 1236.410 1352.760 ;
        RECT 1235.170 1352.560 1235.490 1352.620 ;
        RECT 1236.090 1352.560 1236.410 1352.620 ;
        RECT 1235.630 1304.480 1235.950 1304.540 ;
        RECT 1236.105 1304.480 1236.395 1304.525 ;
        RECT 1235.630 1304.340 1236.395 1304.480 ;
        RECT 1235.630 1304.280 1235.950 1304.340 ;
        RECT 1236.105 1304.295 1236.395 1304.340 ;
        RECT 1236.090 1298.020 1236.410 1298.080 ;
        RECT 1235.895 1297.880 1236.410 1298.020 ;
        RECT 1236.090 1297.820 1236.410 1297.880 ;
        RECT 1236.090 1290.200 1236.410 1290.260 ;
        RECT 1235.895 1290.060 1236.410 1290.200 ;
        RECT 1236.090 1290.000 1236.410 1290.060 ;
        RECT 1236.090 1248.720 1236.410 1248.780 ;
        RECT 1235.895 1248.580 1236.410 1248.720 ;
        RECT 1236.090 1248.520 1236.410 1248.580 ;
        RECT 1234.710 1055.600 1235.030 1055.660 ;
        RECT 1236.090 1055.600 1236.410 1055.660 ;
        RECT 1234.710 1055.460 1236.410 1055.600 ;
        RECT 1234.710 1055.400 1235.030 1055.460 ;
        RECT 1236.090 1055.400 1236.410 1055.460 ;
        RECT 1235.630 966.180 1235.950 966.240 ;
        RECT 1236.090 966.180 1236.410 966.240 ;
        RECT 1235.630 966.040 1236.410 966.180 ;
        RECT 1235.630 965.980 1235.950 966.040 ;
        RECT 1236.090 965.980 1236.410 966.040 ;
        RECT 1235.630 883.700 1235.950 883.960 ;
        RECT 1235.720 883.560 1235.860 883.700 ;
        RECT 1236.090 883.560 1236.410 883.620 ;
        RECT 1235.720 883.420 1236.410 883.560 ;
        RECT 1236.090 883.360 1236.410 883.420 ;
        RECT 1235.645 855.340 1235.935 855.385 ;
        RECT 1236.090 855.340 1236.410 855.400 ;
        RECT 1235.645 855.200 1236.410 855.340 ;
        RECT 1235.645 855.155 1235.935 855.200 ;
        RECT 1236.090 855.140 1236.410 855.200 ;
        RECT 1235.630 807.400 1235.950 807.460 ;
        RECT 1235.435 807.260 1235.950 807.400 ;
        RECT 1235.630 807.200 1235.950 807.260 ;
        RECT 1235.630 766.260 1235.950 766.320 ;
        RECT 1235.260 766.120 1235.950 766.260 ;
        RECT 1235.260 765.980 1235.400 766.120 ;
        RECT 1235.630 766.060 1235.950 766.120 ;
        RECT 1235.170 765.720 1235.490 765.980 ;
        RECT 1236.550 620.740 1236.870 620.800 ;
        RECT 1236.355 620.600 1236.870 620.740 ;
        RECT 1236.550 620.540 1236.870 620.600 ;
        RECT 1235.630 572.800 1235.950 572.860 ;
        RECT 1236.565 572.800 1236.855 572.845 ;
        RECT 1235.630 572.660 1236.855 572.800 ;
        RECT 1235.630 572.600 1235.950 572.660 ;
        RECT 1236.565 572.615 1236.855 572.660 ;
        RECT 1235.630 531.460 1235.950 531.720 ;
        RECT 1235.720 531.040 1235.860 531.460 ;
        RECT 1235.630 530.780 1235.950 531.040 ;
        RECT 1235.630 517.380 1235.950 517.440 ;
        RECT 1235.435 517.240 1235.950 517.380 ;
        RECT 1235.630 517.180 1235.950 517.240 ;
        RECT 1235.645 469.440 1235.935 469.485 ;
        RECT 1236.090 469.440 1236.410 469.500 ;
        RECT 1235.645 469.300 1236.410 469.440 ;
        RECT 1235.645 469.255 1235.935 469.300 ;
        RECT 1236.090 469.240 1236.410 469.300 ;
        RECT 1235.645 400.420 1235.935 400.465 ;
        RECT 1236.090 400.420 1236.410 400.480 ;
        RECT 1235.645 400.280 1236.410 400.420 ;
        RECT 1235.645 400.235 1235.935 400.280 ;
        RECT 1236.090 400.220 1236.410 400.280 ;
        RECT 1235.630 366.080 1235.950 366.140 ;
        RECT 1235.435 365.940 1235.950 366.080 ;
        RECT 1235.630 365.880 1235.950 365.940 ;
        RECT 1236.090 275.980 1236.410 276.040 ;
        RECT 1235.895 275.840 1236.410 275.980 ;
        RECT 1236.090 275.780 1236.410 275.840 ;
        RECT 1236.090 228.040 1236.410 228.100 ;
        RECT 1235.895 227.900 1236.410 228.040 ;
        RECT 1236.090 227.840 1236.410 227.900 ;
        RECT 1236.090 179.420 1236.410 179.480 ;
        RECT 1235.895 179.280 1236.410 179.420 ;
        RECT 1236.090 179.220 1236.410 179.280 ;
        RECT 1236.090 131.820 1236.410 131.880 ;
        RECT 1235.895 131.680 1236.410 131.820 ;
        RECT 1236.090 131.620 1236.410 131.680 ;
        RECT 1235.645 131.140 1235.935 131.185 ;
        RECT 1236.090 131.140 1236.410 131.200 ;
        RECT 1235.645 131.000 1236.410 131.140 ;
        RECT 1235.645 130.955 1235.935 131.000 ;
        RECT 1236.090 130.940 1236.410 131.000 ;
        RECT 222.710 45.800 223.030 45.860 ;
        RECT 1235.645 45.800 1235.935 45.845 ;
        RECT 222.710 45.660 1235.935 45.800 ;
        RECT 222.710 45.600 223.030 45.660 ;
        RECT 1235.645 45.615 1235.935 45.660 ;
      LAYER via ;
        RECT 1235.200 1490.600 1235.460 1490.860 ;
        RECT 1236.580 1490.600 1236.840 1490.860 ;
        RECT 1235.200 1449.120 1235.460 1449.380 ;
        RECT 1236.120 1449.120 1236.380 1449.380 ;
        RECT 1235.200 1352.560 1235.460 1352.820 ;
        RECT 1236.120 1352.560 1236.380 1352.820 ;
        RECT 1235.660 1304.280 1235.920 1304.540 ;
        RECT 1236.120 1297.820 1236.380 1298.080 ;
        RECT 1236.120 1290.000 1236.380 1290.260 ;
        RECT 1236.120 1248.520 1236.380 1248.780 ;
        RECT 1234.740 1055.400 1235.000 1055.660 ;
        RECT 1236.120 1055.400 1236.380 1055.660 ;
        RECT 1235.660 965.980 1235.920 966.240 ;
        RECT 1236.120 965.980 1236.380 966.240 ;
        RECT 1235.660 883.700 1235.920 883.960 ;
        RECT 1236.120 883.360 1236.380 883.620 ;
        RECT 1236.120 855.140 1236.380 855.400 ;
        RECT 1235.660 807.200 1235.920 807.460 ;
        RECT 1235.660 766.060 1235.920 766.320 ;
        RECT 1235.200 765.720 1235.460 765.980 ;
        RECT 1236.580 620.540 1236.840 620.800 ;
        RECT 1235.660 572.600 1235.920 572.860 ;
        RECT 1235.660 531.460 1235.920 531.720 ;
        RECT 1235.660 530.780 1235.920 531.040 ;
        RECT 1235.660 517.180 1235.920 517.440 ;
        RECT 1236.120 469.240 1236.380 469.500 ;
        RECT 1236.120 400.220 1236.380 400.480 ;
        RECT 1235.660 365.880 1235.920 366.140 ;
        RECT 1236.120 275.780 1236.380 276.040 ;
        RECT 1236.120 227.840 1236.380 228.100 ;
        RECT 1236.120 179.220 1236.380 179.480 ;
        RECT 1236.120 131.620 1236.380 131.880 ;
        RECT 1236.120 130.940 1236.380 131.200 ;
        RECT 222.740 45.600 223.000 45.860 ;
      LAYER met2 ;
        RECT 1240.645 1700.410 1240.925 1704.000 ;
        RECT 1238.940 1700.270 1240.925 1700.410 ;
        RECT 1238.940 1687.490 1239.080 1700.270 ;
        RECT 1240.645 1700.000 1240.925 1700.270 ;
        RECT 1235.720 1687.350 1239.080 1687.490 ;
        RECT 1235.720 1655.530 1235.860 1687.350 ;
        RECT 1235.720 1655.390 1236.320 1655.530 ;
        RECT 1236.180 1579.370 1236.320 1655.390 ;
        RECT 1236.180 1579.230 1236.780 1579.370 ;
        RECT 1236.640 1490.890 1236.780 1579.230 ;
        RECT 1235.200 1490.570 1235.460 1490.890 ;
        RECT 1236.580 1490.570 1236.840 1490.890 ;
        RECT 1235.260 1449.410 1235.400 1490.570 ;
        RECT 1235.200 1449.090 1235.460 1449.410 ;
        RECT 1236.120 1449.090 1236.380 1449.410 ;
        RECT 1236.180 1414.810 1236.320 1449.090 ;
        RECT 1236.180 1414.670 1236.780 1414.810 ;
        RECT 1236.640 1414.130 1236.780 1414.670 ;
        RECT 1235.720 1413.990 1236.780 1414.130 ;
        RECT 1235.720 1400.530 1235.860 1413.990 ;
        RECT 1235.260 1400.390 1235.860 1400.530 ;
        RECT 1235.260 1352.850 1235.400 1400.390 ;
        RECT 1235.200 1352.530 1235.460 1352.850 ;
        RECT 1236.120 1352.530 1236.380 1352.850 ;
        RECT 1236.180 1345.450 1236.320 1352.530 ;
        RECT 1235.720 1345.310 1236.320 1345.450 ;
        RECT 1235.720 1304.570 1235.860 1345.310 ;
        RECT 1235.660 1304.250 1235.920 1304.570 ;
        RECT 1236.120 1297.790 1236.380 1298.110 ;
        RECT 1236.180 1290.290 1236.320 1297.790 ;
        RECT 1236.120 1289.970 1236.380 1290.290 ;
        RECT 1236.120 1248.490 1236.380 1248.810 ;
        RECT 1236.180 1199.930 1236.320 1248.490 ;
        RECT 1236.180 1199.790 1236.780 1199.930 ;
        RECT 1236.640 1104.165 1236.780 1199.790 ;
        RECT 1236.570 1103.795 1236.850 1104.165 ;
        RECT 1234.740 1055.370 1235.000 1055.690 ;
        RECT 1236.110 1055.515 1236.390 1055.885 ;
        RECT 1236.120 1055.370 1236.380 1055.515 ;
        RECT 1234.800 1007.605 1234.940 1055.370 ;
        RECT 1234.730 1007.235 1235.010 1007.605 ;
        RECT 1235.650 1007.235 1235.930 1007.605 ;
        RECT 1235.720 966.270 1235.860 1007.235 ;
        RECT 1235.660 965.950 1235.920 966.270 ;
        RECT 1236.120 965.950 1236.380 966.270 ;
        RECT 1236.180 910.930 1236.320 965.950 ;
        RECT 1235.720 910.790 1236.320 910.930 ;
        RECT 1235.720 883.990 1235.860 910.790 ;
        RECT 1235.660 883.670 1235.920 883.990 ;
        RECT 1236.120 883.330 1236.380 883.650 ;
        RECT 1236.180 855.430 1236.320 883.330 ;
        RECT 1236.120 855.110 1236.380 855.430 ;
        RECT 1235.660 807.170 1235.920 807.490 ;
        RECT 1235.720 766.350 1235.860 807.170 ;
        RECT 1235.660 766.030 1235.920 766.350 ;
        RECT 1235.200 765.690 1235.460 766.010 ;
        RECT 1235.260 669.645 1235.400 765.690 ;
        RECT 1235.190 669.275 1235.470 669.645 ;
        RECT 1236.570 668.595 1236.850 668.965 ;
        RECT 1236.640 620.830 1236.780 668.595 ;
        RECT 1236.580 620.510 1236.840 620.830 ;
        RECT 1235.660 572.570 1235.920 572.890 ;
        RECT 1235.720 531.750 1235.860 572.570 ;
        RECT 1235.660 531.430 1235.920 531.750 ;
        RECT 1235.660 530.750 1235.920 531.070 ;
        RECT 1235.720 517.470 1235.860 530.750 ;
        RECT 1235.660 517.150 1235.920 517.470 ;
        RECT 1236.120 469.210 1236.380 469.530 ;
        RECT 1236.180 400.510 1236.320 469.210 ;
        RECT 1236.120 400.190 1236.380 400.510 ;
        RECT 1235.660 365.850 1235.920 366.170 ;
        RECT 1235.720 347.890 1235.860 365.850 ;
        RECT 1235.720 347.750 1236.320 347.890 ;
        RECT 1236.180 276.070 1236.320 347.750 ;
        RECT 1236.120 275.750 1236.380 276.070 ;
        RECT 1236.120 227.810 1236.380 228.130 ;
        RECT 1236.180 179.510 1236.320 227.810 ;
        RECT 1236.120 179.190 1236.380 179.510 ;
        RECT 1236.120 131.590 1236.380 131.910 ;
        RECT 1236.180 131.230 1236.320 131.590 ;
        RECT 1236.120 130.910 1236.380 131.230 ;
        RECT 222.740 45.570 223.000 45.890 ;
        RECT 222.800 2.400 222.940 45.570 ;
        RECT 222.590 -4.800 223.150 2.400 ;
      LAYER via2 ;
        RECT 1236.570 1103.840 1236.850 1104.120 ;
        RECT 1236.110 1055.560 1236.390 1055.840 ;
        RECT 1234.730 1007.280 1235.010 1007.560 ;
        RECT 1235.650 1007.280 1235.930 1007.560 ;
        RECT 1235.190 669.320 1235.470 669.600 ;
        RECT 1236.570 668.640 1236.850 668.920 ;
      LAYER met3 ;
        RECT 1235.830 1104.130 1236.210 1104.140 ;
        RECT 1236.545 1104.130 1236.875 1104.145 ;
        RECT 1235.830 1103.830 1236.875 1104.130 ;
        RECT 1235.830 1103.820 1236.210 1103.830 ;
        RECT 1236.545 1103.815 1236.875 1103.830 ;
        RECT 1236.085 1055.860 1236.415 1055.865 ;
        RECT 1235.830 1055.850 1236.415 1055.860 ;
        RECT 1235.830 1055.550 1236.640 1055.850 ;
        RECT 1235.830 1055.540 1236.415 1055.550 ;
        RECT 1236.085 1055.535 1236.415 1055.540 ;
        RECT 1234.705 1007.570 1235.035 1007.585 ;
        RECT 1235.625 1007.570 1235.955 1007.585 ;
        RECT 1234.705 1007.270 1235.955 1007.570 ;
        RECT 1234.705 1007.255 1235.035 1007.270 ;
        RECT 1235.625 1007.255 1235.955 1007.270 ;
        RECT 1235.165 669.610 1235.495 669.625 ;
        RECT 1235.165 669.310 1236.170 669.610 ;
        RECT 1235.165 669.295 1235.495 669.310 ;
        RECT 1235.870 668.930 1236.170 669.310 ;
        RECT 1236.545 668.930 1236.875 668.945 ;
        RECT 1235.870 668.630 1236.875 668.930 ;
        RECT 1236.545 668.615 1236.875 668.630 ;
      LAYER via3 ;
        RECT 1235.860 1103.820 1236.180 1104.140 ;
        RECT 1235.860 1055.540 1236.180 1055.860 ;
      LAYER met4 ;
        RECT 1235.855 1103.815 1236.185 1104.145 ;
        RECT 1235.870 1055.865 1236.170 1103.815 ;
        RECT 1235.855 1055.535 1236.185 1055.865 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1154.285 1545.725 1154.455 1593.835 ;
        RECT 1154.285 669.545 1154.455 717.655 ;
        RECT 1153.825 241.485 1153.995 303.195 ;
        RECT 1153.825 186.405 1153.995 193.715 ;
        RECT 1153.825 89.845 1153.995 137.955 ;
        RECT 1153.365 55.845 1153.535 62.475 ;
      LAYER mcon ;
        RECT 1154.285 1593.665 1154.455 1593.835 ;
        RECT 1154.285 717.485 1154.455 717.655 ;
        RECT 1153.825 303.025 1153.995 303.195 ;
        RECT 1153.825 193.545 1153.995 193.715 ;
        RECT 1153.825 137.785 1153.995 137.955 ;
        RECT 1153.365 62.305 1153.535 62.475 ;
      LAYER met1 ;
        RECT 1153.750 1607.760 1154.070 1607.820 ;
        RECT 1154.670 1607.760 1154.990 1607.820 ;
        RECT 1153.750 1607.620 1154.990 1607.760 ;
        RECT 1153.750 1607.560 1154.070 1607.620 ;
        RECT 1154.670 1607.560 1154.990 1607.620 ;
        RECT 1154.225 1593.820 1154.515 1593.865 ;
        RECT 1154.670 1593.820 1154.990 1593.880 ;
        RECT 1154.225 1593.680 1154.990 1593.820 ;
        RECT 1154.225 1593.635 1154.515 1593.680 ;
        RECT 1154.670 1593.620 1154.990 1593.680 ;
        RECT 1154.210 1545.880 1154.530 1545.940 ;
        RECT 1154.015 1545.740 1154.530 1545.880 ;
        RECT 1154.210 1545.680 1154.530 1545.740 ;
        RECT 1154.210 966.180 1154.530 966.240 ;
        RECT 1155.130 966.180 1155.450 966.240 ;
        RECT 1154.210 966.040 1155.450 966.180 ;
        RECT 1154.210 965.980 1154.530 966.040 ;
        RECT 1155.130 965.980 1155.450 966.040 ;
        RECT 1154.210 869.620 1154.530 869.680 ;
        RECT 1155.130 869.620 1155.450 869.680 ;
        RECT 1154.210 869.480 1155.450 869.620 ;
        RECT 1154.210 869.420 1154.530 869.480 ;
        RECT 1155.130 869.420 1155.450 869.480 ;
        RECT 1153.290 814.200 1153.610 814.260 ;
        RECT 1153.750 814.200 1154.070 814.260 ;
        RECT 1153.290 814.060 1154.070 814.200 ;
        RECT 1153.290 814.000 1153.610 814.060 ;
        RECT 1153.750 814.000 1154.070 814.060 ;
        RECT 1154.210 717.640 1154.530 717.700 ;
        RECT 1154.015 717.500 1154.530 717.640 ;
        RECT 1154.210 717.440 1154.530 717.500 ;
        RECT 1154.210 669.700 1154.530 669.760 ;
        RECT 1154.015 669.560 1154.530 669.700 ;
        RECT 1154.210 669.500 1154.530 669.560 ;
        RECT 1153.765 303.180 1154.055 303.225 ;
        RECT 1154.210 303.180 1154.530 303.240 ;
        RECT 1153.765 303.040 1154.530 303.180 ;
        RECT 1153.765 302.995 1154.055 303.040 ;
        RECT 1154.210 302.980 1154.530 303.040 ;
        RECT 1153.750 241.640 1154.070 241.700 ;
        RECT 1153.555 241.500 1154.070 241.640 ;
        RECT 1153.750 241.440 1154.070 241.500 ;
        RECT 1153.750 193.700 1154.070 193.760 ;
        RECT 1153.555 193.560 1154.070 193.700 ;
        RECT 1153.750 193.500 1154.070 193.560 ;
        RECT 1153.750 186.560 1154.070 186.620 ;
        RECT 1153.555 186.420 1154.070 186.560 ;
        RECT 1153.750 186.360 1154.070 186.420 ;
        RECT 1153.750 137.940 1154.070 138.000 ;
        RECT 1153.555 137.800 1154.070 137.940 ;
        RECT 1153.750 137.740 1154.070 137.800 ;
        RECT 1153.750 90.000 1154.070 90.060 ;
        RECT 1153.555 89.860 1154.070 90.000 ;
        RECT 1153.750 89.800 1154.070 89.860 ;
        RECT 1153.305 62.460 1153.595 62.505 ;
        RECT 1153.750 62.460 1154.070 62.520 ;
        RECT 1153.305 62.320 1154.070 62.460 ;
        RECT 1153.305 62.275 1153.595 62.320 ;
        RECT 1153.750 62.260 1154.070 62.320 ;
        RECT 1153.290 56.000 1153.610 56.060 ;
        RECT 1153.095 55.860 1153.610 56.000 ;
        RECT 1153.290 55.800 1153.610 55.860 ;
        RECT 1153.290 38.320 1153.610 38.380 ;
        RECT 1138.200 38.180 1153.610 38.320 ;
        RECT 20.310 37.980 20.630 38.040 ;
        RECT 1138.200 37.980 1138.340 38.180 ;
        RECT 1153.290 38.120 1153.610 38.180 ;
        RECT 20.310 37.840 1138.340 37.980 ;
        RECT 20.310 37.780 20.630 37.840 ;
      LAYER via ;
        RECT 1153.780 1607.560 1154.040 1607.820 ;
        RECT 1154.700 1607.560 1154.960 1607.820 ;
        RECT 1154.700 1593.620 1154.960 1593.880 ;
        RECT 1154.240 1545.680 1154.500 1545.940 ;
        RECT 1154.240 965.980 1154.500 966.240 ;
        RECT 1155.160 965.980 1155.420 966.240 ;
        RECT 1154.240 869.420 1154.500 869.680 ;
        RECT 1155.160 869.420 1155.420 869.680 ;
        RECT 1153.320 814.000 1153.580 814.260 ;
        RECT 1153.780 814.000 1154.040 814.260 ;
        RECT 1154.240 717.440 1154.500 717.700 ;
        RECT 1154.240 669.500 1154.500 669.760 ;
        RECT 1154.240 302.980 1154.500 303.240 ;
        RECT 1153.780 241.440 1154.040 241.700 ;
        RECT 1153.780 193.500 1154.040 193.760 ;
        RECT 1153.780 186.360 1154.040 186.620 ;
        RECT 1153.780 137.740 1154.040 138.000 ;
        RECT 1153.780 89.800 1154.040 90.060 ;
        RECT 1153.780 62.260 1154.040 62.520 ;
        RECT 1153.320 55.800 1153.580 56.060 ;
        RECT 20.340 37.780 20.600 38.040 ;
        RECT 1153.320 38.120 1153.580 38.380 ;
      LAYER met2 ;
        RECT 1156.925 1701.090 1157.205 1704.000 ;
        RECT 1155.220 1700.950 1157.205 1701.090 ;
        RECT 1155.220 1688.850 1155.360 1700.950 ;
        RECT 1156.925 1700.000 1157.205 1700.950 ;
        RECT 1153.840 1688.710 1155.360 1688.850 ;
        RECT 1153.840 1607.850 1153.980 1688.710 ;
        RECT 1153.780 1607.530 1154.040 1607.850 ;
        RECT 1154.700 1607.530 1154.960 1607.850 ;
        RECT 1154.760 1593.910 1154.900 1607.530 ;
        RECT 1154.700 1593.590 1154.960 1593.910 ;
        RECT 1154.240 1545.650 1154.500 1545.970 ;
        RECT 1154.300 1027.890 1154.440 1545.650 ;
        RECT 1153.840 1027.750 1154.440 1027.890 ;
        RECT 1153.840 1014.405 1153.980 1027.750 ;
        RECT 1153.770 1014.035 1154.050 1014.405 ;
        RECT 1155.150 1014.035 1155.430 1014.405 ;
        RECT 1155.220 966.270 1155.360 1014.035 ;
        RECT 1154.240 965.950 1154.500 966.270 ;
        RECT 1155.160 965.950 1155.420 966.270 ;
        RECT 1154.300 931.330 1154.440 965.950 ;
        RECT 1153.840 931.190 1154.440 931.330 ;
        RECT 1153.840 917.845 1153.980 931.190 ;
        RECT 1153.770 917.475 1154.050 917.845 ;
        RECT 1155.150 917.475 1155.430 917.845 ;
        RECT 1155.220 869.710 1155.360 917.475 ;
        RECT 1154.240 869.390 1154.500 869.710 ;
        RECT 1155.160 869.390 1155.420 869.710 ;
        RECT 1154.300 834.770 1154.440 869.390 ;
        RECT 1153.840 834.630 1154.440 834.770 ;
        RECT 1153.840 814.290 1153.980 834.630 ;
        RECT 1153.320 813.970 1153.580 814.290 ;
        RECT 1153.780 813.970 1154.040 814.290 ;
        RECT 1153.380 766.205 1153.520 813.970 ;
        RECT 1153.310 765.835 1153.590 766.205 ;
        RECT 1154.230 765.835 1154.510 766.205 ;
        RECT 1154.300 717.730 1154.440 765.835 ;
        RECT 1154.240 717.410 1154.500 717.730 ;
        RECT 1154.240 669.470 1154.500 669.790 ;
        RECT 1154.300 303.270 1154.440 669.470 ;
        RECT 1154.240 302.950 1154.500 303.270 ;
        RECT 1153.780 241.410 1154.040 241.730 ;
        RECT 1153.840 193.790 1153.980 241.410 ;
        RECT 1153.780 193.470 1154.040 193.790 ;
        RECT 1153.780 186.330 1154.040 186.650 ;
        RECT 1153.840 138.030 1153.980 186.330 ;
        RECT 1153.780 137.710 1154.040 138.030 ;
        RECT 1153.780 89.770 1154.040 90.090 ;
        RECT 1153.840 62.550 1153.980 89.770 ;
        RECT 1153.780 62.230 1154.040 62.550 ;
        RECT 1153.320 55.770 1153.580 56.090 ;
        RECT 1153.380 38.410 1153.520 55.770 ;
        RECT 1153.320 38.090 1153.580 38.410 ;
        RECT 20.340 37.750 20.600 38.070 ;
        RECT 20.400 2.400 20.540 37.750 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 1153.770 1014.080 1154.050 1014.360 ;
        RECT 1155.150 1014.080 1155.430 1014.360 ;
        RECT 1153.770 917.520 1154.050 917.800 ;
        RECT 1155.150 917.520 1155.430 917.800 ;
        RECT 1153.310 765.880 1153.590 766.160 ;
        RECT 1154.230 765.880 1154.510 766.160 ;
      LAYER met3 ;
        RECT 1153.745 1014.370 1154.075 1014.385 ;
        RECT 1155.125 1014.370 1155.455 1014.385 ;
        RECT 1153.745 1014.070 1155.455 1014.370 ;
        RECT 1153.745 1014.055 1154.075 1014.070 ;
        RECT 1155.125 1014.055 1155.455 1014.070 ;
        RECT 1153.745 917.810 1154.075 917.825 ;
        RECT 1155.125 917.810 1155.455 917.825 ;
        RECT 1153.745 917.510 1155.455 917.810 ;
        RECT 1153.745 917.495 1154.075 917.510 ;
        RECT 1155.125 917.495 1155.455 917.510 ;
        RECT 1153.285 766.170 1153.615 766.185 ;
        RECT 1154.205 766.170 1154.535 766.185 ;
        RECT 1153.285 765.870 1154.535 766.170 ;
        RECT 1153.285 765.855 1153.615 765.870 ;
        RECT 1154.205 765.855 1154.535 765.870 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1137.725 34.765 1137.895 38.335 ;
      LAYER mcon ;
        RECT 1137.725 38.165 1137.895 38.335 ;
      LAYER met1 ;
        RECT 44.230 38.320 44.550 38.380 ;
        RECT 1137.665 38.320 1137.955 38.365 ;
        RECT 44.230 38.180 1137.955 38.320 ;
        RECT 44.230 38.120 44.550 38.180 ;
        RECT 1137.665 38.135 1137.955 38.180 ;
        RECT 1137.665 34.920 1137.955 34.965 ;
        RECT 1167.090 34.920 1167.410 34.980 ;
        RECT 1137.665 34.780 1167.410 34.920 ;
        RECT 1137.665 34.735 1137.955 34.780 ;
        RECT 1167.090 34.720 1167.410 34.780 ;
      LAYER via ;
        RECT 44.260 38.120 44.520 38.380 ;
        RECT 1167.120 34.720 1167.380 34.980 ;
      LAYER met2 ;
        RECT 1167.045 1700.000 1167.325 1704.000 ;
        RECT 44.260 38.090 44.520 38.410 ;
        RECT 44.320 2.400 44.460 38.090 ;
        RECT 1167.180 35.010 1167.320 1700.000 ;
        RECT 1167.120 34.690 1167.380 35.010 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 246.630 46.140 246.950 46.200 ;
        RECT 1249.430 46.140 1249.750 46.200 ;
        RECT 246.630 46.000 1249.750 46.140 ;
        RECT 246.630 45.940 246.950 46.000 ;
        RECT 1249.430 45.940 1249.750 46.000 ;
      LAYER via ;
        RECT 246.660 45.940 246.920 46.200 ;
        RECT 1249.460 45.940 1249.720 46.200 ;
      LAYER met2 ;
        RECT 1250.305 1700.410 1250.585 1704.000 ;
        RECT 1249.520 1700.270 1250.585 1700.410 ;
        RECT 1249.520 46.230 1249.660 1700.270 ;
        RECT 1250.305 1700.000 1250.585 1700.270 ;
        RECT 246.660 45.910 246.920 46.230 ;
        RECT 1249.460 45.910 1249.720 46.230 ;
        RECT 246.720 2.400 246.860 45.910 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1256.330 821.480 1256.650 821.740 ;
        RECT 1256.420 821.060 1256.560 821.480 ;
        RECT 1256.330 820.800 1256.650 821.060 ;
        RECT 268.710 51.580 269.030 51.640 ;
        RECT 1256.330 51.580 1256.650 51.640 ;
        RECT 268.710 51.440 1256.650 51.580 ;
        RECT 268.710 51.380 269.030 51.440 ;
        RECT 1256.330 51.380 1256.650 51.440 ;
        RECT 264.110 15.880 264.430 15.940 ;
        RECT 268.710 15.880 269.030 15.940 ;
        RECT 264.110 15.740 269.030 15.880 ;
        RECT 264.110 15.680 264.430 15.740 ;
        RECT 268.710 15.680 269.030 15.740 ;
      LAYER via ;
        RECT 1256.360 821.480 1256.620 821.740 ;
        RECT 1256.360 820.800 1256.620 821.060 ;
        RECT 268.740 51.380 269.000 51.640 ;
        RECT 1256.360 51.380 1256.620 51.640 ;
        RECT 264.140 15.680 264.400 15.940 ;
        RECT 268.740 15.680 269.000 15.940 ;
      LAYER met2 ;
        RECT 1257.665 1700.410 1257.945 1704.000 ;
        RECT 1256.420 1700.270 1257.945 1700.410 ;
        RECT 1256.420 821.770 1256.560 1700.270 ;
        RECT 1257.665 1700.000 1257.945 1700.270 ;
        RECT 1256.360 821.450 1256.620 821.770 ;
        RECT 1256.360 820.770 1256.620 821.090 ;
        RECT 1256.420 51.670 1256.560 820.770 ;
        RECT 268.740 51.350 269.000 51.670 ;
        RECT 1256.360 51.350 1256.620 51.670 ;
        RECT 268.800 15.970 268.940 51.350 ;
        RECT 264.140 15.650 264.400 15.970 ;
        RECT 268.740 15.650 269.000 15.970 ;
        RECT 264.200 2.400 264.340 15.650 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.510 51.920 282.830 51.980 ;
        RECT 1263.230 51.920 1263.550 51.980 ;
        RECT 282.510 51.780 1263.550 51.920 ;
        RECT 282.510 51.720 282.830 51.780 ;
        RECT 1263.230 51.720 1263.550 51.780 ;
      LAYER via ;
        RECT 282.540 51.720 282.800 51.980 ;
        RECT 1263.260 51.720 1263.520 51.980 ;
      LAYER met2 ;
        RECT 1265.025 1700.410 1265.305 1704.000 ;
        RECT 1263.320 1700.270 1265.305 1700.410 ;
        RECT 1263.320 52.010 1263.460 1700.270 ;
        RECT 1265.025 1700.000 1265.305 1700.270 ;
        RECT 282.540 51.690 282.800 52.010 ;
        RECT 1263.260 51.690 1263.520 52.010 ;
        RECT 282.600 17.410 282.740 51.690 ;
        RECT 282.140 17.270 282.740 17.410 ;
        RECT 282.140 2.400 282.280 17.270 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 303.210 52.260 303.530 52.320 ;
        RECT 1270.130 52.260 1270.450 52.320 ;
        RECT 303.210 52.120 1270.450 52.260 ;
        RECT 303.210 52.060 303.530 52.120 ;
        RECT 1270.130 52.060 1270.450 52.120 ;
        RECT 299.990 16.900 300.310 16.960 ;
        RECT 303.210 16.900 303.530 16.960 ;
        RECT 299.990 16.760 303.530 16.900 ;
        RECT 299.990 16.700 300.310 16.760 ;
        RECT 303.210 16.700 303.530 16.760 ;
      LAYER via ;
        RECT 303.240 52.060 303.500 52.320 ;
        RECT 1270.160 52.060 1270.420 52.320 ;
        RECT 300.020 16.700 300.280 16.960 ;
        RECT 303.240 16.700 303.500 16.960 ;
      LAYER met2 ;
        RECT 1272.385 1700.410 1272.665 1704.000 ;
        RECT 1270.220 1700.270 1272.665 1700.410 ;
        RECT 1270.220 52.350 1270.360 1700.270 ;
        RECT 1272.385 1700.000 1272.665 1700.270 ;
        RECT 303.240 52.030 303.500 52.350 ;
        RECT 1270.160 52.030 1270.420 52.350 ;
        RECT 303.300 16.990 303.440 52.030 ;
        RECT 300.020 16.670 300.280 16.990 ;
        RECT 303.240 16.670 303.500 16.990 ;
        RECT 300.080 2.400 300.220 16.670 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 323.910 52.600 324.230 52.660 ;
        RECT 1277.950 52.600 1278.270 52.660 ;
        RECT 323.910 52.460 1278.270 52.600 ;
        RECT 323.910 52.400 324.230 52.460 ;
        RECT 1277.950 52.400 1278.270 52.460 ;
        RECT 317.930 16.220 318.250 16.280 ;
        RECT 323.910 16.220 324.230 16.280 ;
        RECT 317.930 16.080 324.230 16.220 ;
        RECT 317.930 16.020 318.250 16.080 ;
        RECT 323.910 16.020 324.230 16.080 ;
      LAYER via ;
        RECT 323.940 52.400 324.200 52.660 ;
        RECT 1277.980 52.400 1278.240 52.660 ;
        RECT 317.960 16.020 318.220 16.280 ;
        RECT 323.940 16.020 324.200 16.280 ;
      LAYER met2 ;
        RECT 1279.745 1700.410 1280.025 1704.000 ;
        RECT 1278.040 1700.270 1280.025 1700.410 ;
        RECT 1278.040 52.690 1278.180 1700.270 ;
        RECT 1279.745 1700.000 1280.025 1700.270 ;
        RECT 323.940 52.370 324.200 52.690 ;
        RECT 1277.980 52.370 1278.240 52.690 ;
        RECT 324.000 16.310 324.140 52.370 ;
        RECT 317.960 15.990 318.220 16.310 ;
        RECT 323.940 15.990 324.200 16.310 ;
        RECT 318.020 2.400 318.160 15.990 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 335.870 26.420 336.190 26.480 ;
        RECT 1284.850 26.420 1285.170 26.480 ;
        RECT 335.870 26.280 1285.170 26.420 ;
        RECT 335.870 26.220 336.190 26.280 ;
        RECT 1284.850 26.220 1285.170 26.280 ;
      LAYER via ;
        RECT 335.900 26.220 336.160 26.480 ;
        RECT 1284.880 26.220 1285.140 26.480 ;
      LAYER met2 ;
        RECT 1287.105 1700.410 1287.385 1704.000 ;
        RECT 1284.940 1700.270 1287.385 1700.410 ;
        RECT 1284.940 26.510 1285.080 1700.270 ;
        RECT 1287.105 1700.000 1287.385 1700.270 ;
        RECT 335.900 26.190 336.160 26.510 ;
        RECT 1284.880 26.190 1285.140 26.510 ;
        RECT 335.960 2.400 336.100 26.190 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1290.830 1673.040 1291.150 1673.100 ;
        RECT 1292.670 1673.040 1292.990 1673.100 ;
        RECT 1290.830 1672.900 1292.990 1673.040 ;
        RECT 1290.830 1672.840 1291.150 1672.900 ;
        RECT 1292.670 1672.840 1292.990 1672.900 ;
        RECT 358.410 65.860 358.730 65.920 ;
        RECT 1290.830 65.860 1291.150 65.920 ;
        RECT 358.410 65.720 1291.150 65.860 ;
        RECT 358.410 65.660 358.730 65.720 ;
        RECT 1290.830 65.660 1291.150 65.720 ;
        RECT 353.350 16.560 353.670 16.620 ;
        RECT 358.410 16.560 358.730 16.620 ;
        RECT 353.350 16.420 358.730 16.560 ;
        RECT 353.350 16.360 353.670 16.420 ;
        RECT 358.410 16.360 358.730 16.420 ;
      LAYER via ;
        RECT 1290.860 1672.840 1291.120 1673.100 ;
        RECT 1292.700 1672.840 1292.960 1673.100 ;
        RECT 358.440 65.660 358.700 65.920 ;
        RECT 1290.860 65.660 1291.120 65.920 ;
        RECT 353.380 16.360 353.640 16.620 ;
        RECT 358.440 16.360 358.700 16.620 ;
      LAYER met2 ;
        RECT 1294.465 1700.410 1294.745 1704.000 ;
        RECT 1292.760 1700.270 1294.745 1700.410 ;
        RECT 1292.760 1673.130 1292.900 1700.270 ;
        RECT 1294.465 1700.000 1294.745 1700.270 ;
        RECT 1290.860 1672.810 1291.120 1673.130 ;
        RECT 1292.700 1672.810 1292.960 1673.130 ;
        RECT 1290.920 65.950 1291.060 1672.810 ;
        RECT 358.440 65.630 358.700 65.950 ;
        RECT 1290.860 65.630 1291.120 65.950 ;
        RECT 358.500 16.650 358.640 65.630 ;
        RECT 353.380 16.330 353.640 16.650 ;
        RECT 358.440 16.330 358.700 16.650 ;
        RECT 353.440 2.400 353.580 16.330 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1299.185 1594.005 1299.355 1642.115 ;
        RECT 1298.265 1483.505 1298.435 1511.555 ;
        RECT 1298.265 1207.765 1298.435 1273.215 ;
        RECT 1298.725 737.885 1298.895 772.735 ;
        RECT 1298.265 614.125 1298.435 662.235 ;
        RECT 1298.725 386.325 1298.895 475.915 ;
        RECT 1299.645 228.225 1299.815 282.795 ;
        RECT 1297.805 131.665 1297.975 179.435 ;
        RECT 1297.805 89.505 1297.975 131.155 ;
      LAYER mcon ;
        RECT 1299.185 1641.945 1299.355 1642.115 ;
        RECT 1298.265 1511.385 1298.435 1511.555 ;
        RECT 1298.265 1273.045 1298.435 1273.215 ;
        RECT 1298.725 772.565 1298.895 772.735 ;
        RECT 1298.265 662.065 1298.435 662.235 ;
        RECT 1298.725 475.745 1298.895 475.915 ;
        RECT 1299.645 282.625 1299.815 282.795 ;
        RECT 1297.805 179.265 1297.975 179.435 ;
        RECT 1297.805 130.985 1297.975 131.155 ;
      LAYER met1 ;
        RECT 1298.190 1689.020 1298.510 1689.080 ;
        RECT 1300.490 1689.020 1300.810 1689.080 ;
        RECT 1298.190 1688.880 1300.810 1689.020 ;
        RECT 1298.190 1688.820 1298.510 1688.880 ;
        RECT 1300.490 1688.820 1300.810 1688.880 ;
        RECT 1298.190 1656.040 1298.510 1656.100 ;
        RECT 1299.110 1656.040 1299.430 1656.100 ;
        RECT 1298.190 1655.900 1299.430 1656.040 ;
        RECT 1298.190 1655.840 1298.510 1655.900 ;
        RECT 1299.110 1655.840 1299.430 1655.900 ;
        RECT 1299.110 1642.100 1299.430 1642.160 ;
        RECT 1298.915 1641.960 1299.430 1642.100 ;
        RECT 1299.110 1641.900 1299.430 1641.960 ;
        RECT 1299.125 1594.160 1299.415 1594.205 ;
        RECT 1299.570 1594.160 1299.890 1594.220 ;
        RECT 1299.125 1594.020 1299.890 1594.160 ;
        RECT 1299.125 1593.975 1299.415 1594.020 ;
        RECT 1299.570 1593.960 1299.890 1594.020 ;
        RECT 1298.650 1559.480 1298.970 1559.540 ;
        RECT 1299.570 1559.480 1299.890 1559.540 ;
        RECT 1298.650 1559.340 1299.890 1559.480 ;
        RECT 1298.650 1559.280 1298.970 1559.340 ;
        RECT 1299.570 1559.280 1299.890 1559.340 ;
        RECT 1298.205 1511.540 1298.495 1511.585 ;
        RECT 1298.650 1511.540 1298.970 1511.600 ;
        RECT 1298.205 1511.400 1298.970 1511.540 ;
        RECT 1298.205 1511.355 1298.495 1511.400 ;
        RECT 1298.650 1511.340 1298.970 1511.400 ;
        RECT 1298.190 1483.660 1298.510 1483.720 ;
        RECT 1297.995 1483.520 1298.510 1483.660 ;
        RECT 1298.190 1483.460 1298.510 1483.520 ;
        RECT 1298.190 1345.620 1298.510 1345.680 ;
        RECT 1298.650 1345.620 1298.970 1345.680 ;
        RECT 1298.190 1345.480 1298.970 1345.620 ;
        RECT 1298.190 1345.420 1298.510 1345.480 ;
        RECT 1298.650 1345.420 1298.970 1345.480 ;
        RECT 1298.205 1273.200 1298.495 1273.245 ;
        RECT 1298.650 1273.200 1298.970 1273.260 ;
        RECT 1298.205 1273.060 1298.970 1273.200 ;
        RECT 1298.205 1273.015 1298.495 1273.060 ;
        RECT 1298.650 1273.000 1298.970 1273.060 ;
        RECT 1298.190 1207.920 1298.510 1207.980 ;
        RECT 1297.995 1207.780 1298.510 1207.920 ;
        RECT 1298.190 1207.720 1298.510 1207.780 ;
        RECT 1297.730 1152.500 1298.050 1152.560 ;
        RECT 1298.190 1152.500 1298.510 1152.560 ;
        RECT 1297.730 1152.360 1298.510 1152.500 ;
        RECT 1297.730 1152.300 1298.050 1152.360 ;
        RECT 1298.190 1152.300 1298.510 1152.360 ;
        RECT 1298.650 966.180 1298.970 966.240 ;
        RECT 1299.570 966.180 1299.890 966.240 ;
        RECT 1298.650 966.040 1299.890 966.180 ;
        RECT 1298.650 965.980 1298.970 966.040 ;
        RECT 1299.570 965.980 1299.890 966.040 ;
        RECT 1298.650 869.620 1298.970 869.680 ;
        RECT 1299.570 869.620 1299.890 869.680 ;
        RECT 1298.650 869.480 1299.890 869.620 ;
        RECT 1298.650 869.420 1298.970 869.480 ;
        RECT 1299.570 869.420 1299.890 869.480 ;
        RECT 1298.650 772.720 1298.970 772.780 ;
        RECT 1298.455 772.580 1298.970 772.720 ;
        RECT 1298.650 772.520 1298.970 772.580 ;
        RECT 1298.650 738.040 1298.970 738.100 ;
        RECT 1298.455 737.900 1298.970 738.040 ;
        RECT 1298.650 737.840 1298.970 737.900 ;
        RECT 1298.190 690.100 1298.510 690.160 ;
        RECT 1299.110 690.100 1299.430 690.160 ;
        RECT 1298.190 689.960 1299.430 690.100 ;
        RECT 1298.190 689.900 1298.510 689.960 ;
        RECT 1299.110 689.900 1299.430 689.960 ;
        RECT 1298.205 662.220 1298.495 662.265 ;
        RECT 1298.650 662.220 1298.970 662.280 ;
        RECT 1298.205 662.080 1298.970 662.220 ;
        RECT 1298.205 662.035 1298.495 662.080 ;
        RECT 1298.650 662.020 1298.970 662.080 ;
        RECT 1298.190 614.280 1298.510 614.340 ;
        RECT 1297.995 614.140 1298.510 614.280 ;
        RECT 1298.190 614.080 1298.510 614.140 ;
        RECT 1298.650 566.000 1298.970 566.060 ;
        RECT 1299.570 566.000 1299.890 566.060 ;
        RECT 1298.650 565.860 1299.890 566.000 ;
        RECT 1298.650 565.800 1298.970 565.860 ;
        RECT 1299.570 565.800 1299.890 565.860 ;
        RECT 1298.190 475.900 1298.510 475.960 ;
        RECT 1298.665 475.900 1298.955 475.945 ;
        RECT 1298.190 475.760 1298.955 475.900 ;
        RECT 1298.190 475.700 1298.510 475.760 ;
        RECT 1298.665 475.715 1298.955 475.760 ;
        RECT 1298.650 386.480 1298.970 386.540 ;
        RECT 1298.455 386.340 1298.970 386.480 ;
        RECT 1298.650 386.280 1298.970 386.340 ;
        RECT 1298.650 313.180 1298.970 313.440 ;
        RECT 1298.740 313.040 1298.880 313.180 ;
        RECT 1299.570 313.040 1299.890 313.100 ;
        RECT 1298.740 312.900 1299.890 313.040 ;
        RECT 1299.570 312.840 1299.890 312.900 ;
        RECT 1299.570 282.780 1299.890 282.840 ;
        RECT 1299.570 282.640 1300.085 282.780 ;
        RECT 1299.570 282.580 1299.890 282.640 ;
        RECT 1299.585 228.380 1299.875 228.425 ;
        RECT 1298.740 228.240 1299.875 228.380 ;
        RECT 1298.740 228.100 1298.880 228.240 ;
        RECT 1299.585 228.195 1299.875 228.240 ;
        RECT 1298.650 227.840 1298.970 228.100 ;
        RECT 1298.190 185.880 1298.510 185.940 ;
        RECT 1298.650 185.880 1298.970 185.940 ;
        RECT 1298.190 185.740 1298.970 185.880 ;
        RECT 1298.190 185.680 1298.510 185.740 ;
        RECT 1298.650 185.680 1298.970 185.740 ;
        RECT 1297.745 179.420 1298.035 179.465 ;
        RECT 1298.190 179.420 1298.510 179.480 ;
        RECT 1297.745 179.280 1298.510 179.420 ;
        RECT 1297.745 179.235 1298.035 179.280 ;
        RECT 1298.190 179.220 1298.510 179.280 ;
        RECT 1297.730 131.820 1298.050 131.880 ;
        RECT 1297.535 131.680 1298.050 131.820 ;
        RECT 1297.730 131.620 1298.050 131.680 ;
        RECT 1297.730 131.140 1298.050 131.200 ;
        RECT 1297.535 131.000 1298.050 131.140 ;
        RECT 1297.730 130.940 1298.050 131.000 ;
        RECT 1297.730 89.660 1298.050 89.720 ;
        RECT 1297.535 89.520 1298.050 89.660 ;
        RECT 1297.730 89.460 1298.050 89.520 ;
        RECT 372.210 72.320 372.530 72.380 ;
        RECT 1297.730 72.320 1298.050 72.380 ;
        RECT 372.210 72.180 1298.050 72.320 ;
        RECT 372.210 72.120 372.530 72.180 ;
        RECT 1297.730 72.120 1298.050 72.180 ;
      LAYER via ;
        RECT 1298.220 1688.820 1298.480 1689.080 ;
        RECT 1300.520 1688.820 1300.780 1689.080 ;
        RECT 1298.220 1655.840 1298.480 1656.100 ;
        RECT 1299.140 1655.840 1299.400 1656.100 ;
        RECT 1299.140 1641.900 1299.400 1642.160 ;
        RECT 1299.600 1593.960 1299.860 1594.220 ;
        RECT 1298.680 1559.280 1298.940 1559.540 ;
        RECT 1299.600 1559.280 1299.860 1559.540 ;
        RECT 1298.680 1511.340 1298.940 1511.600 ;
        RECT 1298.220 1483.460 1298.480 1483.720 ;
        RECT 1298.220 1345.420 1298.480 1345.680 ;
        RECT 1298.680 1345.420 1298.940 1345.680 ;
        RECT 1298.680 1273.000 1298.940 1273.260 ;
        RECT 1298.220 1207.720 1298.480 1207.980 ;
        RECT 1297.760 1152.300 1298.020 1152.560 ;
        RECT 1298.220 1152.300 1298.480 1152.560 ;
        RECT 1298.680 965.980 1298.940 966.240 ;
        RECT 1299.600 965.980 1299.860 966.240 ;
        RECT 1298.680 869.420 1298.940 869.680 ;
        RECT 1299.600 869.420 1299.860 869.680 ;
        RECT 1298.680 772.520 1298.940 772.780 ;
        RECT 1298.680 737.840 1298.940 738.100 ;
        RECT 1298.220 689.900 1298.480 690.160 ;
        RECT 1299.140 689.900 1299.400 690.160 ;
        RECT 1298.680 662.020 1298.940 662.280 ;
        RECT 1298.220 614.080 1298.480 614.340 ;
        RECT 1298.680 565.800 1298.940 566.060 ;
        RECT 1299.600 565.800 1299.860 566.060 ;
        RECT 1298.220 475.700 1298.480 475.960 ;
        RECT 1298.680 386.280 1298.940 386.540 ;
        RECT 1298.680 313.180 1298.940 313.440 ;
        RECT 1299.600 312.840 1299.860 313.100 ;
        RECT 1299.600 282.580 1299.860 282.840 ;
        RECT 1298.680 227.840 1298.940 228.100 ;
        RECT 1298.220 185.680 1298.480 185.940 ;
        RECT 1298.680 185.680 1298.940 185.940 ;
        RECT 1298.220 179.220 1298.480 179.480 ;
        RECT 1297.760 131.620 1298.020 131.880 ;
        RECT 1297.760 130.940 1298.020 131.200 ;
        RECT 1297.760 89.460 1298.020 89.720 ;
        RECT 372.240 72.120 372.500 72.380 ;
        RECT 1297.760 72.120 1298.020 72.380 ;
      LAYER met2 ;
        RECT 1301.825 1700.410 1302.105 1704.000 ;
        RECT 1300.580 1700.270 1302.105 1700.410 ;
        RECT 1300.580 1689.110 1300.720 1700.270 ;
        RECT 1301.825 1700.000 1302.105 1700.270 ;
        RECT 1298.220 1688.790 1298.480 1689.110 ;
        RECT 1300.520 1688.790 1300.780 1689.110 ;
        RECT 1298.280 1656.130 1298.420 1688.790 ;
        RECT 1298.220 1655.810 1298.480 1656.130 ;
        RECT 1299.140 1655.810 1299.400 1656.130 ;
        RECT 1299.200 1642.190 1299.340 1655.810 ;
        RECT 1299.140 1641.870 1299.400 1642.190 ;
        RECT 1299.600 1593.930 1299.860 1594.250 ;
        RECT 1299.660 1559.570 1299.800 1593.930 ;
        RECT 1298.680 1559.250 1298.940 1559.570 ;
        RECT 1299.600 1559.250 1299.860 1559.570 ;
        RECT 1298.740 1511.630 1298.880 1559.250 ;
        RECT 1298.680 1511.310 1298.940 1511.630 ;
        RECT 1298.220 1483.430 1298.480 1483.750 ;
        RECT 1298.280 1345.710 1298.420 1483.430 ;
        RECT 1298.220 1345.390 1298.480 1345.710 ;
        RECT 1298.680 1345.390 1298.940 1345.710 ;
        RECT 1298.740 1328.450 1298.880 1345.390 ;
        RECT 1297.820 1328.310 1298.880 1328.450 ;
        RECT 1297.820 1317.570 1297.960 1328.310 ;
        RECT 1297.820 1317.430 1298.420 1317.570 ;
        RECT 1298.280 1303.970 1298.420 1317.430 ;
        RECT 1298.280 1303.830 1298.880 1303.970 ;
        RECT 1298.740 1273.290 1298.880 1303.830 ;
        RECT 1298.680 1272.970 1298.940 1273.290 ;
        RECT 1298.220 1207.690 1298.480 1208.010 ;
        RECT 1298.280 1152.590 1298.420 1207.690 ;
        RECT 1297.760 1152.270 1298.020 1152.590 ;
        RECT 1298.220 1152.270 1298.480 1152.590 ;
        RECT 1297.820 1135.330 1297.960 1152.270 ;
        RECT 1297.820 1135.190 1298.420 1135.330 ;
        RECT 1298.280 1110.965 1298.420 1135.190 ;
        RECT 1298.210 1110.595 1298.490 1110.965 ;
        RECT 1298.670 1109.235 1298.950 1109.605 ;
        RECT 1298.740 1027.890 1298.880 1109.235 ;
        RECT 1298.280 1027.750 1298.880 1027.890 ;
        RECT 1298.280 1014.405 1298.420 1027.750 ;
        RECT 1298.210 1014.035 1298.490 1014.405 ;
        RECT 1299.590 1014.035 1299.870 1014.405 ;
        RECT 1299.660 966.270 1299.800 1014.035 ;
        RECT 1298.680 965.950 1298.940 966.270 ;
        RECT 1299.600 965.950 1299.860 966.270 ;
        RECT 1298.740 931.330 1298.880 965.950 ;
        RECT 1298.280 931.190 1298.880 931.330 ;
        RECT 1298.280 917.845 1298.420 931.190 ;
        RECT 1298.210 917.475 1298.490 917.845 ;
        RECT 1299.590 917.475 1299.870 917.845 ;
        RECT 1299.660 869.710 1299.800 917.475 ;
        RECT 1298.680 869.390 1298.940 869.710 ;
        RECT 1299.600 869.390 1299.860 869.710 ;
        RECT 1298.740 787.170 1298.880 869.390 ;
        RECT 1298.280 787.030 1298.880 787.170 ;
        RECT 1298.280 786.490 1298.420 787.030 ;
        RECT 1298.280 786.350 1298.880 786.490 ;
        RECT 1298.740 772.810 1298.880 786.350 ;
        RECT 1298.680 772.490 1298.940 772.810 ;
        RECT 1298.680 737.810 1298.940 738.130 ;
        RECT 1298.740 724.610 1298.880 737.810 ;
        RECT 1298.740 724.470 1299.340 724.610 ;
        RECT 1298.280 690.190 1298.420 690.345 ;
        RECT 1299.200 690.190 1299.340 724.470 ;
        RECT 1298.220 689.930 1298.480 690.190 ;
        RECT 1298.220 689.870 1298.880 689.930 ;
        RECT 1299.140 689.870 1299.400 690.190 ;
        RECT 1298.280 689.790 1298.880 689.870 ;
        RECT 1298.740 662.310 1298.880 689.790 ;
        RECT 1298.680 661.990 1298.940 662.310 ;
        RECT 1298.220 614.050 1298.480 614.370 ;
        RECT 1298.280 613.770 1298.420 614.050 ;
        RECT 1298.670 613.770 1298.950 613.885 ;
        RECT 1298.280 613.630 1298.950 613.770 ;
        RECT 1298.670 613.515 1298.950 613.630 ;
        RECT 1299.590 613.515 1299.870 613.885 ;
        RECT 1299.660 566.090 1299.800 613.515 ;
        RECT 1298.680 565.770 1298.940 566.090 ;
        RECT 1299.600 565.770 1299.860 566.090 ;
        RECT 1298.740 524.010 1298.880 565.770 ;
        RECT 1298.280 523.870 1298.880 524.010 ;
        RECT 1298.280 475.990 1298.420 523.870 ;
        RECT 1298.220 475.670 1298.480 475.990 ;
        RECT 1298.680 386.250 1298.940 386.570 ;
        RECT 1298.740 313.470 1298.880 386.250 ;
        RECT 1298.680 313.150 1298.940 313.470 ;
        RECT 1299.600 312.810 1299.860 313.130 ;
        RECT 1299.660 282.870 1299.800 312.810 ;
        RECT 1299.600 282.550 1299.860 282.870 ;
        RECT 1298.680 227.810 1298.940 228.130 ;
        RECT 1298.740 185.970 1298.880 227.810 ;
        RECT 1298.220 185.650 1298.480 185.970 ;
        RECT 1298.680 185.650 1298.940 185.970 ;
        RECT 1298.280 179.510 1298.420 185.650 ;
        RECT 1298.220 179.190 1298.480 179.510 ;
        RECT 1297.760 131.590 1298.020 131.910 ;
        RECT 1297.820 131.230 1297.960 131.590 ;
        RECT 1297.760 130.910 1298.020 131.230 ;
        RECT 1297.760 89.430 1298.020 89.750 ;
        RECT 1297.820 72.410 1297.960 89.430 ;
        RECT 372.240 72.090 372.500 72.410 ;
        RECT 1297.760 72.090 1298.020 72.410 ;
        RECT 372.300 16.900 372.440 72.090 ;
        RECT 371.380 16.760 372.440 16.900 ;
        RECT 371.380 2.400 371.520 16.760 ;
        RECT 371.170 -4.800 371.730 2.400 ;
      LAYER via2 ;
        RECT 1298.210 1110.640 1298.490 1110.920 ;
        RECT 1298.670 1109.280 1298.950 1109.560 ;
        RECT 1298.210 1014.080 1298.490 1014.360 ;
        RECT 1299.590 1014.080 1299.870 1014.360 ;
        RECT 1298.210 917.520 1298.490 917.800 ;
        RECT 1299.590 917.520 1299.870 917.800 ;
        RECT 1298.670 613.560 1298.950 613.840 ;
        RECT 1299.590 613.560 1299.870 613.840 ;
      LAYER met3 ;
        RECT 1298.185 1110.930 1298.515 1110.945 ;
        RECT 1297.510 1110.630 1298.515 1110.930 ;
        RECT 1297.510 1109.570 1297.810 1110.630 ;
        RECT 1298.185 1110.615 1298.515 1110.630 ;
        RECT 1298.645 1109.570 1298.975 1109.585 ;
        RECT 1297.510 1109.270 1298.975 1109.570 ;
        RECT 1298.645 1109.255 1298.975 1109.270 ;
        RECT 1298.185 1014.370 1298.515 1014.385 ;
        RECT 1299.565 1014.370 1299.895 1014.385 ;
        RECT 1298.185 1014.070 1299.895 1014.370 ;
        RECT 1298.185 1014.055 1298.515 1014.070 ;
        RECT 1299.565 1014.055 1299.895 1014.070 ;
        RECT 1298.185 917.810 1298.515 917.825 ;
        RECT 1299.565 917.810 1299.895 917.825 ;
        RECT 1298.185 917.510 1299.895 917.810 ;
        RECT 1298.185 917.495 1298.515 917.510 ;
        RECT 1299.565 917.495 1299.895 917.510 ;
        RECT 1298.645 613.850 1298.975 613.865 ;
        RECT 1299.565 613.850 1299.895 613.865 ;
        RECT 1298.645 613.550 1299.895 613.850 ;
        RECT 1298.645 613.535 1298.975 613.550 ;
        RECT 1299.565 613.535 1299.895 613.550 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1304.630 1678.140 1304.950 1678.200 ;
        RECT 1307.390 1678.140 1307.710 1678.200 ;
        RECT 1304.630 1678.000 1307.710 1678.140 ;
        RECT 1304.630 1677.940 1304.950 1678.000 ;
        RECT 1307.390 1677.940 1307.710 1678.000 ;
        RECT 392.910 72.660 393.230 72.720 ;
        RECT 1304.630 72.660 1304.950 72.720 ;
        RECT 392.910 72.520 1304.950 72.660 ;
        RECT 392.910 72.460 393.230 72.520 ;
        RECT 1304.630 72.460 1304.950 72.520 ;
        RECT 389.230 16.220 389.550 16.280 ;
        RECT 392.910 16.220 393.230 16.280 ;
        RECT 389.230 16.080 393.230 16.220 ;
        RECT 389.230 16.020 389.550 16.080 ;
        RECT 392.910 16.020 393.230 16.080 ;
      LAYER via ;
        RECT 1304.660 1677.940 1304.920 1678.200 ;
        RECT 1307.420 1677.940 1307.680 1678.200 ;
        RECT 392.940 72.460 393.200 72.720 ;
        RECT 1304.660 72.460 1304.920 72.720 ;
        RECT 389.260 16.020 389.520 16.280 ;
        RECT 392.940 16.020 393.200 16.280 ;
      LAYER met2 ;
        RECT 1309.185 1700.410 1309.465 1704.000 ;
        RECT 1307.480 1700.270 1309.465 1700.410 ;
        RECT 1307.480 1678.230 1307.620 1700.270 ;
        RECT 1309.185 1700.000 1309.465 1700.270 ;
        RECT 1304.660 1677.910 1304.920 1678.230 ;
        RECT 1307.420 1677.910 1307.680 1678.230 ;
        RECT 1304.720 72.750 1304.860 1677.910 ;
        RECT 392.940 72.430 393.200 72.750 ;
        RECT 1304.660 72.430 1304.920 72.750 ;
        RECT 393.000 16.310 393.140 72.430 ;
        RECT 389.260 15.990 389.520 16.310 ;
        RECT 392.940 15.990 393.200 16.310 ;
        RECT 389.320 2.400 389.460 15.990 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1312.985 1483.505 1313.155 1498.295 ;
        RECT 1312.985 614.125 1313.155 662.235 ;
        RECT 1312.525 524.365 1312.695 548.675 ;
        RECT 1312.985 421.345 1313.155 469.115 ;
      LAYER mcon ;
        RECT 1312.985 1498.125 1313.155 1498.295 ;
        RECT 1312.985 662.065 1313.155 662.235 ;
        RECT 1312.525 548.505 1312.695 548.675 ;
        RECT 1312.985 468.945 1313.155 469.115 ;
      LAYER met1 ;
        RECT 1312.910 1678.140 1313.230 1678.200 ;
        RECT 1315.210 1678.140 1315.530 1678.200 ;
        RECT 1312.910 1678.000 1315.530 1678.140 ;
        RECT 1312.910 1677.940 1313.230 1678.000 ;
        RECT 1315.210 1677.940 1315.530 1678.000 ;
        RECT 1312.910 1656.040 1313.230 1656.100 ;
        RECT 1313.830 1656.040 1314.150 1656.100 ;
        RECT 1312.910 1655.900 1314.150 1656.040 ;
        RECT 1312.910 1655.840 1313.230 1655.900 ;
        RECT 1313.830 1655.840 1314.150 1655.900 ;
        RECT 1313.830 1607.900 1314.150 1608.160 ;
        RECT 1313.920 1607.420 1314.060 1607.900 ;
        RECT 1314.290 1607.420 1314.610 1607.480 ;
        RECT 1313.920 1607.280 1314.610 1607.420 ;
        RECT 1314.290 1607.220 1314.610 1607.280 ;
        RECT 1312.925 1498.280 1313.215 1498.325 ;
        RECT 1313.370 1498.280 1313.690 1498.340 ;
        RECT 1312.925 1498.140 1313.690 1498.280 ;
        RECT 1312.925 1498.095 1313.215 1498.140 ;
        RECT 1313.370 1498.080 1313.690 1498.140 ;
        RECT 1312.910 1483.660 1313.230 1483.720 ;
        RECT 1312.715 1483.520 1313.230 1483.660 ;
        RECT 1312.910 1483.460 1313.230 1483.520 ;
        RECT 1311.530 1290.200 1311.850 1290.260 ;
        RECT 1312.910 1290.200 1313.230 1290.260 ;
        RECT 1311.530 1290.060 1313.230 1290.200 ;
        RECT 1311.530 1290.000 1311.850 1290.060 ;
        RECT 1312.910 1290.000 1313.230 1290.060 ;
        RECT 1312.450 1200.780 1312.770 1200.840 ;
        RECT 1312.910 1200.780 1313.230 1200.840 ;
        RECT 1312.450 1200.640 1313.230 1200.780 ;
        RECT 1312.450 1200.580 1312.770 1200.640 ;
        RECT 1312.910 1200.580 1313.230 1200.640 ;
        RECT 1312.450 1060.700 1312.770 1060.760 ;
        RECT 1313.370 1060.700 1313.690 1060.760 ;
        RECT 1312.450 1060.560 1313.690 1060.700 ;
        RECT 1312.450 1060.500 1312.770 1060.560 ;
        RECT 1313.370 1060.500 1313.690 1060.560 ;
        RECT 1312.450 1014.460 1312.770 1014.520 ;
        RECT 1312.910 1014.460 1313.230 1014.520 ;
        RECT 1312.450 1014.320 1313.230 1014.460 ;
        RECT 1312.450 1014.260 1312.770 1014.320 ;
        RECT 1312.910 1014.260 1313.230 1014.320 ;
        RECT 1312.925 662.220 1313.215 662.265 ;
        RECT 1313.370 662.220 1313.690 662.280 ;
        RECT 1312.925 662.080 1313.690 662.220 ;
        RECT 1312.925 662.035 1313.215 662.080 ;
        RECT 1313.370 662.020 1313.690 662.080 ;
        RECT 1312.910 614.280 1313.230 614.340 ;
        RECT 1312.715 614.140 1313.230 614.280 ;
        RECT 1312.910 614.080 1313.230 614.140 ;
        RECT 1312.465 548.660 1312.755 548.705 ;
        RECT 1312.910 548.660 1313.230 548.720 ;
        RECT 1312.465 548.520 1313.230 548.660 ;
        RECT 1312.465 548.475 1312.755 548.520 ;
        RECT 1312.910 548.460 1313.230 548.520 ;
        RECT 1312.450 524.520 1312.770 524.580 ;
        RECT 1312.255 524.380 1312.770 524.520 ;
        RECT 1312.450 524.320 1312.770 524.380 ;
        RECT 1312.450 476.240 1312.770 476.300 ;
        RECT 1312.910 476.240 1313.230 476.300 ;
        RECT 1312.450 476.100 1313.230 476.240 ;
        RECT 1312.450 476.040 1312.770 476.100 ;
        RECT 1312.910 476.040 1313.230 476.100 ;
        RECT 1312.910 469.100 1313.230 469.160 ;
        RECT 1312.715 468.960 1313.230 469.100 ;
        RECT 1312.910 468.900 1313.230 468.960 ;
        RECT 1312.925 421.500 1313.215 421.545 ;
        RECT 1312.925 421.360 1313.600 421.500 ;
        RECT 1312.925 421.315 1313.215 421.360 ;
        RECT 1313.460 421.220 1313.600 421.360 ;
        RECT 1313.370 420.960 1313.690 421.220 ;
        RECT 1313.830 307.260 1314.150 307.320 ;
        RECT 1314.750 307.260 1315.070 307.320 ;
        RECT 1313.830 307.120 1315.070 307.260 ;
        RECT 1313.830 307.060 1314.150 307.120 ;
        RECT 1314.750 307.060 1315.070 307.120 ;
        RECT 1313.370 145.080 1313.690 145.140 ;
        RECT 1313.830 145.080 1314.150 145.140 ;
        RECT 1313.370 144.940 1314.150 145.080 ;
        RECT 1313.370 144.880 1313.690 144.940 ;
        RECT 1313.830 144.880 1314.150 144.940 ;
        RECT 413.610 73.000 413.930 73.060 ;
        RECT 1312.910 73.000 1313.230 73.060 ;
        RECT 413.610 72.860 1313.230 73.000 ;
        RECT 413.610 72.800 413.930 72.860 ;
        RECT 1312.910 72.800 1313.230 72.860 ;
        RECT 407.170 16.220 407.490 16.280 ;
        RECT 413.610 16.220 413.930 16.280 ;
        RECT 407.170 16.080 413.930 16.220 ;
        RECT 407.170 16.020 407.490 16.080 ;
        RECT 413.610 16.020 413.930 16.080 ;
      LAYER via ;
        RECT 1312.940 1677.940 1313.200 1678.200 ;
        RECT 1315.240 1677.940 1315.500 1678.200 ;
        RECT 1312.940 1655.840 1313.200 1656.100 ;
        RECT 1313.860 1655.840 1314.120 1656.100 ;
        RECT 1313.860 1607.900 1314.120 1608.160 ;
        RECT 1314.320 1607.220 1314.580 1607.480 ;
        RECT 1313.400 1498.080 1313.660 1498.340 ;
        RECT 1312.940 1483.460 1313.200 1483.720 ;
        RECT 1311.560 1290.000 1311.820 1290.260 ;
        RECT 1312.940 1290.000 1313.200 1290.260 ;
        RECT 1312.480 1200.580 1312.740 1200.840 ;
        RECT 1312.940 1200.580 1313.200 1200.840 ;
        RECT 1312.480 1060.500 1312.740 1060.760 ;
        RECT 1313.400 1060.500 1313.660 1060.760 ;
        RECT 1312.480 1014.260 1312.740 1014.520 ;
        RECT 1312.940 1014.260 1313.200 1014.520 ;
        RECT 1313.400 662.020 1313.660 662.280 ;
        RECT 1312.940 614.080 1313.200 614.340 ;
        RECT 1312.940 548.460 1313.200 548.720 ;
        RECT 1312.480 524.320 1312.740 524.580 ;
        RECT 1312.480 476.040 1312.740 476.300 ;
        RECT 1312.940 476.040 1313.200 476.300 ;
        RECT 1312.940 468.900 1313.200 469.160 ;
        RECT 1313.400 420.960 1313.660 421.220 ;
        RECT 1313.860 307.060 1314.120 307.320 ;
        RECT 1314.780 307.060 1315.040 307.320 ;
        RECT 1313.400 144.880 1313.660 145.140 ;
        RECT 1313.860 144.880 1314.120 145.140 ;
        RECT 413.640 72.800 413.900 73.060 ;
        RECT 1312.940 72.800 1313.200 73.060 ;
        RECT 407.200 16.020 407.460 16.280 ;
        RECT 413.640 16.020 413.900 16.280 ;
      LAYER met2 ;
        RECT 1316.545 1700.410 1316.825 1704.000 ;
        RECT 1315.300 1700.270 1316.825 1700.410 ;
        RECT 1315.300 1678.230 1315.440 1700.270 ;
        RECT 1316.545 1700.000 1316.825 1700.270 ;
        RECT 1312.940 1677.910 1313.200 1678.230 ;
        RECT 1315.240 1677.910 1315.500 1678.230 ;
        RECT 1313.000 1656.130 1313.140 1677.910 ;
        RECT 1312.940 1655.810 1313.200 1656.130 ;
        RECT 1313.860 1655.810 1314.120 1656.130 ;
        RECT 1313.920 1608.190 1314.060 1655.810 ;
        RECT 1313.860 1607.870 1314.120 1608.190 ;
        RECT 1314.320 1607.190 1314.580 1607.510 ;
        RECT 1314.380 1546.050 1314.520 1607.190 ;
        RECT 1313.460 1545.910 1314.520 1546.050 ;
        RECT 1313.460 1498.370 1313.600 1545.910 ;
        RECT 1313.400 1498.050 1313.660 1498.370 ;
        RECT 1312.940 1483.430 1313.200 1483.750 ;
        RECT 1313.000 1345.565 1313.140 1483.430 ;
        RECT 1312.930 1345.195 1313.210 1345.565 ;
        RECT 1313.390 1344.515 1313.670 1344.885 ;
        RECT 1313.460 1317.570 1313.600 1344.515 ;
        RECT 1313.000 1317.430 1313.600 1317.570 ;
        RECT 1313.000 1290.290 1313.140 1317.430 ;
        RECT 1311.560 1289.970 1311.820 1290.290 ;
        RECT 1312.940 1289.970 1313.200 1290.290 ;
        RECT 1311.620 1242.205 1311.760 1289.970 ;
        RECT 1311.550 1241.835 1311.830 1242.205 ;
        RECT 1312.470 1241.835 1312.750 1242.205 ;
        RECT 1312.540 1200.870 1312.680 1241.835 ;
        RECT 1313.000 1200.870 1313.140 1201.025 ;
        RECT 1312.480 1200.550 1312.740 1200.870 ;
        RECT 1312.940 1200.610 1313.200 1200.870 ;
        RECT 1312.940 1200.550 1313.600 1200.610 ;
        RECT 1313.000 1200.470 1313.600 1200.550 ;
        RECT 1313.460 1060.790 1313.600 1200.470 ;
        RECT 1312.480 1060.470 1312.740 1060.790 ;
        RECT 1313.400 1060.470 1313.660 1060.790 ;
        RECT 1312.540 1014.550 1312.680 1060.470 ;
        RECT 1312.480 1014.230 1312.740 1014.550 ;
        RECT 1312.940 1014.405 1313.200 1014.550 ;
        RECT 1312.930 1014.035 1313.210 1014.405 ;
        RECT 1313.390 1013.355 1313.670 1013.725 ;
        RECT 1313.460 931.330 1313.600 1013.355 ;
        RECT 1313.000 931.190 1313.600 931.330 ;
        RECT 1313.000 917.845 1313.140 931.190 ;
        RECT 1312.930 917.475 1313.210 917.845 ;
        RECT 1313.390 916.795 1313.670 917.165 ;
        RECT 1313.460 787.170 1313.600 916.795 ;
        RECT 1313.000 787.030 1313.600 787.170 ;
        RECT 1313.000 786.490 1313.140 787.030 ;
        RECT 1313.000 786.350 1313.600 786.490 ;
        RECT 1313.460 748.410 1313.600 786.350 ;
        RECT 1313.460 748.270 1314.520 748.410 ;
        RECT 1314.380 738.210 1314.520 748.270 ;
        RECT 1313.920 738.070 1314.520 738.210 ;
        RECT 1313.920 724.440 1314.060 738.070 ;
        RECT 1313.920 724.300 1314.520 724.440 ;
        RECT 1314.380 676.445 1314.520 724.300 ;
        RECT 1313.390 676.075 1313.670 676.445 ;
        RECT 1314.310 676.075 1314.590 676.445 ;
        RECT 1313.460 662.310 1313.600 676.075 ;
        RECT 1313.400 661.990 1313.660 662.310 ;
        RECT 1312.940 614.050 1313.200 614.370 ;
        RECT 1313.000 548.750 1313.140 614.050 ;
        RECT 1312.940 548.430 1313.200 548.750 ;
        RECT 1312.480 524.290 1312.740 524.610 ;
        RECT 1312.540 476.330 1312.680 524.290 ;
        RECT 1312.480 476.010 1312.740 476.330 ;
        RECT 1312.940 476.010 1313.200 476.330 ;
        RECT 1313.000 469.190 1313.140 476.010 ;
        RECT 1312.940 468.870 1313.200 469.190 ;
        RECT 1313.400 420.930 1313.660 421.250 ;
        RECT 1313.460 331.005 1313.600 420.930 ;
        RECT 1313.390 330.635 1313.670 331.005 ;
        RECT 1314.770 330.635 1315.050 331.005 ;
        RECT 1314.840 307.350 1314.980 330.635 ;
        RECT 1313.860 307.030 1314.120 307.350 ;
        RECT 1314.780 307.030 1315.040 307.350 ;
        RECT 1313.920 145.170 1314.060 307.030 ;
        RECT 1313.400 144.850 1313.660 145.170 ;
        RECT 1313.860 144.850 1314.120 145.170 ;
        RECT 1313.460 110.570 1313.600 144.850 ;
        RECT 1313.000 110.430 1313.600 110.570 ;
        RECT 1313.000 73.090 1313.140 110.430 ;
        RECT 413.640 72.770 413.900 73.090 ;
        RECT 1312.940 72.770 1313.200 73.090 ;
        RECT 413.700 16.310 413.840 72.770 ;
        RECT 407.200 15.990 407.460 16.310 ;
        RECT 413.640 15.990 413.900 16.310 ;
        RECT 407.260 2.400 407.400 15.990 ;
        RECT 407.050 -4.800 407.610 2.400 ;
      LAYER via2 ;
        RECT 1312.930 1345.240 1313.210 1345.520 ;
        RECT 1313.390 1344.560 1313.670 1344.840 ;
        RECT 1311.550 1241.880 1311.830 1242.160 ;
        RECT 1312.470 1241.880 1312.750 1242.160 ;
        RECT 1312.930 1014.080 1313.210 1014.360 ;
        RECT 1313.390 1013.400 1313.670 1013.680 ;
        RECT 1312.930 917.520 1313.210 917.800 ;
        RECT 1313.390 916.840 1313.670 917.120 ;
        RECT 1313.390 676.120 1313.670 676.400 ;
        RECT 1314.310 676.120 1314.590 676.400 ;
        RECT 1313.390 330.680 1313.670 330.960 ;
        RECT 1314.770 330.680 1315.050 330.960 ;
      LAYER met3 ;
        RECT 1312.905 1345.530 1313.235 1345.545 ;
        RECT 1312.905 1345.215 1313.450 1345.530 ;
        RECT 1313.150 1344.865 1313.450 1345.215 ;
        RECT 1313.150 1344.550 1313.695 1344.865 ;
        RECT 1313.365 1344.535 1313.695 1344.550 ;
        RECT 1311.525 1242.170 1311.855 1242.185 ;
        RECT 1312.445 1242.170 1312.775 1242.185 ;
        RECT 1311.525 1241.870 1312.775 1242.170 ;
        RECT 1311.525 1241.855 1311.855 1241.870 ;
        RECT 1312.445 1241.855 1312.775 1241.870 ;
        RECT 1312.905 1014.370 1313.235 1014.385 ;
        RECT 1312.905 1014.055 1313.450 1014.370 ;
        RECT 1313.150 1013.705 1313.450 1014.055 ;
        RECT 1313.150 1013.390 1313.695 1013.705 ;
        RECT 1313.365 1013.375 1313.695 1013.390 ;
        RECT 1312.905 917.810 1313.235 917.825 ;
        RECT 1312.905 917.495 1313.450 917.810 ;
        RECT 1313.150 917.145 1313.450 917.495 ;
        RECT 1313.150 916.830 1313.695 917.145 ;
        RECT 1313.365 916.815 1313.695 916.830 ;
        RECT 1313.365 676.410 1313.695 676.425 ;
        RECT 1314.285 676.410 1314.615 676.425 ;
        RECT 1313.365 676.110 1314.615 676.410 ;
        RECT 1313.365 676.095 1313.695 676.110 ;
        RECT 1314.285 676.095 1314.615 676.110 ;
        RECT 1313.365 330.970 1313.695 330.985 ;
        RECT 1314.745 330.970 1315.075 330.985 ;
        RECT 1313.365 330.670 1315.075 330.970 ;
        RECT 1313.365 330.655 1313.695 330.670 ;
        RECT 1314.745 330.655 1315.075 330.670 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 68.150 44.780 68.470 44.840 ;
        RECT 1173.990 44.780 1174.310 44.840 ;
        RECT 68.150 44.640 1174.310 44.780 ;
        RECT 68.150 44.580 68.470 44.640 ;
        RECT 1173.990 44.580 1174.310 44.640 ;
      LAYER via ;
        RECT 68.180 44.580 68.440 44.840 ;
        RECT 1174.020 44.580 1174.280 44.840 ;
      LAYER met2 ;
        RECT 1176.705 1700.410 1176.985 1704.000 ;
        RECT 1175.460 1700.270 1176.985 1700.410 ;
        RECT 1175.460 1678.650 1175.600 1700.270 ;
        RECT 1176.705 1700.000 1176.985 1700.270 ;
        RECT 1174.080 1678.510 1175.600 1678.650 ;
        RECT 1174.080 44.870 1174.220 1678.510 ;
        RECT 68.180 44.550 68.440 44.870 ;
        RECT 1174.020 44.550 1174.280 44.870 ;
        RECT 68.240 2.400 68.380 44.550 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1318.430 1678.140 1318.750 1678.200 ;
        RECT 1322.110 1678.140 1322.430 1678.200 ;
        RECT 1318.430 1678.000 1322.430 1678.140 ;
        RECT 1318.430 1677.940 1318.750 1678.000 ;
        RECT 1322.110 1677.940 1322.430 1678.000 ;
        RECT 427.410 73.340 427.730 73.400 ;
        RECT 1318.430 73.340 1318.750 73.400 ;
        RECT 427.410 73.200 1318.750 73.340 ;
        RECT 427.410 73.140 427.730 73.200 ;
        RECT 1318.430 73.140 1318.750 73.200 ;
        RECT 424.650 16.220 424.970 16.280 ;
        RECT 427.410 16.220 427.730 16.280 ;
        RECT 424.650 16.080 427.730 16.220 ;
        RECT 424.650 16.020 424.970 16.080 ;
        RECT 427.410 16.020 427.730 16.080 ;
      LAYER via ;
        RECT 1318.460 1677.940 1318.720 1678.200 ;
        RECT 1322.140 1677.940 1322.400 1678.200 ;
        RECT 427.440 73.140 427.700 73.400 ;
        RECT 1318.460 73.140 1318.720 73.400 ;
        RECT 424.680 16.020 424.940 16.280 ;
        RECT 427.440 16.020 427.700 16.280 ;
      LAYER met2 ;
        RECT 1323.905 1700.410 1324.185 1704.000 ;
        RECT 1322.200 1700.270 1324.185 1700.410 ;
        RECT 1322.200 1678.230 1322.340 1700.270 ;
        RECT 1323.905 1700.000 1324.185 1700.270 ;
        RECT 1318.460 1677.910 1318.720 1678.230 ;
        RECT 1322.140 1677.910 1322.400 1678.230 ;
        RECT 1318.520 73.430 1318.660 1677.910 ;
        RECT 427.440 73.110 427.700 73.430 ;
        RECT 1318.460 73.110 1318.720 73.430 ;
        RECT 427.500 16.310 427.640 73.110 ;
        RECT 424.680 15.990 424.940 16.310 ;
        RECT 427.440 15.990 427.700 16.310 ;
        RECT 424.740 2.400 424.880 15.990 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1325.330 1678.140 1325.650 1678.200 ;
        RECT 1329.470 1678.140 1329.790 1678.200 ;
        RECT 1325.330 1678.000 1329.790 1678.140 ;
        RECT 1325.330 1677.940 1325.650 1678.000 ;
        RECT 1329.470 1677.940 1329.790 1678.000 ;
        RECT 448.110 73.680 448.430 73.740 ;
        RECT 1325.330 73.680 1325.650 73.740 ;
        RECT 448.110 73.540 1325.650 73.680 ;
        RECT 448.110 73.480 448.430 73.540 ;
        RECT 1325.330 73.480 1325.650 73.540 ;
        RECT 442.590 16.220 442.910 16.280 ;
        RECT 448.110 16.220 448.430 16.280 ;
        RECT 442.590 16.080 448.430 16.220 ;
        RECT 442.590 16.020 442.910 16.080 ;
        RECT 448.110 16.020 448.430 16.080 ;
      LAYER via ;
        RECT 1325.360 1677.940 1325.620 1678.200 ;
        RECT 1329.500 1677.940 1329.760 1678.200 ;
        RECT 448.140 73.480 448.400 73.740 ;
        RECT 1325.360 73.480 1325.620 73.740 ;
        RECT 442.620 16.020 442.880 16.280 ;
        RECT 448.140 16.020 448.400 16.280 ;
      LAYER met2 ;
        RECT 1331.265 1700.410 1331.545 1704.000 ;
        RECT 1329.560 1700.270 1331.545 1700.410 ;
        RECT 1329.560 1678.230 1329.700 1700.270 ;
        RECT 1331.265 1700.000 1331.545 1700.270 ;
        RECT 1325.360 1677.910 1325.620 1678.230 ;
        RECT 1329.500 1677.910 1329.760 1678.230 ;
        RECT 1325.420 73.770 1325.560 1677.910 ;
        RECT 448.140 73.450 448.400 73.770 ;
        RECT 1325.360 73.450 1325.620 73.770 ;
        RECT 448.200 16.310 448.340 73.450 ;
        RECT 442.620 15.990 442.880 16.310 ;
        RECT 448.140 15.990 448.400 16.310 ;
        RECT 442.680 2.400 442.820 15.990 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1332.230 1678.140 1332.550 1678.200 ;
        RECT 1336.830 1678.140 1337.150 1678.200 ;
        RECT 1332.230 1678.000 1337.150 1678.140 ;
        RECT 1332.230 1677.940 1332.550 1678.000 ;
        RECT 1336.830 1677.940 1337.150 1678.000 ;
        RECT 461.910 74.020 462.230 74.080 ;
        RECT 1332.230 74.020 1332.550 74.080 ;
        RECT 461.910 73.880 1332.550 74.020 ;
        RECT 461.910 73.820 462.230 73.880 ;
        RECT 1332.230 73.820 1332.550 73.880 ;
      LAYER via ;
        RECT 1332.260 1677.940 1332.520 1678.200 ;
        RECT 1336.860 1677.940 1337.120 1678.200 ;
        RECT 461.940 73.820 462.200 74.080 ;
        RECT 1332.260 73.820 1332.520 74.080 ;
      LAYER met2 ;
        RECT 1338.165 1700.410 1338.445 1704.000 ;
        RECT 1336.920 1700.270 1338.445 1700.410 ;
        RECT 1336.920 1678.230 1337.060 1700.270 ;
        RECT 1338.165 1700.000 1338.445 1700.270 ;
        RECT 1332.260 1677.910 1332.520 1678.230 ;
        RECT 1336.860 1677.910 1337.120 1678.230 ;
        RECT 1332.320 74.110 1332.460 1677.910 ;
        RECT 461.940 73.790 462.200 74.110 ;
        RECT 1332.260 73.790 1332.520 74.110 ;
        RECT 462.000 16.730 462.140 73.790 ;
        RECT 460.620 16.590 462.140 16.730 ;
        RECT 460.620 2.400 460.760 16.590 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 482.610 74.360 482.930 74.420 ;
        RECT 1346.030 74.360 1346.350 74.420 ;
        RECT 482.610 74.220 1346.350 74.360 ;
        RECT 482.610 74.160 482.930 74.220 ;
        RECT 1346.030 74.160 1346.350 74.220 ;
        RECT 478.470 15.540 478.790 15.600 ;
        RECT 482.610 15.540 482.930 15.600 ;
        RECT 478.470 15.400 482.930 15.540 ;
        RECT 478.470 15.340 478.790 15.400 ;
        RECT 482.610 15.340 482.930 15.400 ;
      LAYER via ;
        RECT 482.640 74.160 482.900 74.420 ;
        RECT 1346.060 74.160 1346.320 74.420 ;
        RECT 478.500 15.340 478.760 15.600 ;
        RECT 482.640 15.340 482.900 15.600 ;
      LAYER met2 ;
        RECT 1345.525 1700.410 1345.805 1704.000 ;
        RECT 1345.525 1700.270 1346.260 1700.410 ;
        RECT 1345.525 1700.000 1345.805 1700.270 ;
        RECT 1346.120 74.450 1346.260 1700.270 ;
        RECT 482.640 74.130 482.900 74.450 ;
        RECT 1346.060 74.130 1346.320 74.450 ;
        RECT 482.700 15.630 482.840 74.130 ;
        RECT 478.500 15.310 478.760 15.630 ;
        RECT 482.640 15.310 482.900 15.630 ;
        RECT 478.560 2.400 478.700 15.310 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 496.410 74.700 496.730 74.760 ;
        RECT 1352.930 74.700 1353.250 74.760 ;
        RECT 496.410 74.560 1353.250 74.700 ;
        RECT 496.410 74.500 496.730 74.560 ;
        RECT 1352.930 74.500 1353.250 74.560 ;
      LAYER via ;
        RECT 496.440 74.500 496.700 74.760 ;
        RECT 1352.960 74.500 1353.220 74.760 ;
      LAYER met2 ;
        RECT 1352.885 1700.000 1353.165 1704.000 ;
        RECT 1353.020 74.790 1353.160 1700.000 ;
        RECT 496.440 74.470 496.700 74.790 ;
        RECT 1352.960 74.470 1353.220 74.790 ;
        RECT 496.500 2.400 496.640 74.470 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 517.110 75.040 517.430 75.100 ;
        RECT 1359.830 75.040 1360.150 75.100 ;
        RECT 517.110 74.900 1360.150 75.040 ;
        RECT 517.110 74.840 517.430 74.900 ;
        RECT 1359.830 74.840 1360.150 74.900 ;
        RECT 513.890 15.540 514.210 15.600 ;
        RECT 517.110 15.540 517.430 15.600 ;
        RECT 513.890 15.400 517.430 15.540 ;
        RECT 513.890 15.340 514.210 15.400 ;
        RECT 517.110 15.340 517.430 15.400 ;
      LAYER via ;
        RECT 517.140 74.840 517.400 75.100 ;
        RECT 1359.860 74.840 1360.120 75.100 ;
        RECT 513.920 15.340 514.180 15.600 ;
        RECT 517.140 15.340 517.400 15.600 ;
      LAYER met2 ;
        RECT 1360.245 1700.410 1360.525 1704.000 ;
        RECT 1359.920 1700.270 1360.525 1700.410 ;
        RECT 1359.920 75.130 1360.060 1700.270 ;
        RECT 1360.245 1700.000 1360.525 1700.270 ;
        RECT 517.140 74.810 517.400 75.130 ;
        RECT 1359.860 74.810 1360.120 75.130 ;
        RECT 517.200 15.630 517.340 74.810 ;
        RECT 513.920 15.310 514.180 15.630 ;
        RECT 517.140 15.310 517.400 15.630 ;
        RECT 513.980 2.400 514.120 15.310 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 537.350 75.380 537.670 75.440 ;
        RECT 1366.730 75.380 1367.050 75.440 ;
        RECT 537.350 75.240 1367.050 75.380 ;
        RECT 537.350 75.180 537.670 75.240 ;
        RECT 1366.730 75.180 1367.050 75.240 ;
        RECT 531.830 15.540 532.150 15.600 ;
        RECT 537.350 15.540 537.670 15.600 ;
        RECT 531.830 15.400 537.670 15.540 ;
        RECT 531.830 15.340 532.150 15.400 ;
        RECT 537.350 15.340 537.670 15.400 ;
      LAYER via ;
        RECT 537.380 75.180 537.640 75.440 ;
        RECT 1366.760 75.180 1367.020 75.440 ;
        RECT 531.860 15.340 532.120 15.600 ;
        RECT 537.380 15.340 537.640 15.600 ;
      LAYER met2 ;
        RECT 1367.605 1700.410 1367.885 1704.000 ;
        RECT 1366.820 1700.270 1367.885 1700.410 ;
        RECT 1366.820 75.470 1366.960 1700.270 ;
        RECT 1367.605 1700.000 1367.885 1700.270 ;
        RECT 537.380 75.150 537.640 75.470 ;
        RECT 1366.760 75.150 1367.020 75.470 ;
        RECT 537.440 15.630 537.580 75.150 ;
        RECT 531.860 15.310 532.120 15.630 ;
        RECT 537.380 15.310 537.640 15.630 ;
        RECT 531.920 2.400 532.060 15.310 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 75.720 551.930 75.780 ;
        RECT 1373.630 75.720 1373.950 75.780 ;
        RECT 551.610 75.580 1373.950 75.720 ;
        RECT 551.610 75.520 551.930 75.580 ;
        RECT 1373.630 75.520 1373.950 75.580 ;
      LAYER via ;
        RECT 551.640 75.520 551.900 75.780 ;
        RECT 1373.660 75.520 1373.920 75.780 ;
      LAYER met2 ;
        RECT 1374.965 1700.410 1375.245 1704.000 ;
        RECT 1373.720 1700.270 1375.245 1700.410 ;
        RECT 1373.720 75.810 1373.860 1700.270 ;
        RECT 1374.965 1700.000 1375.245 1700.270 ;
        RECT 551.640 75.490 551.900 75.810 ;
        RECT 1373.660 75.490 1373.920 75.810 ;
        RECT 551.700 17.410 551.840 75.490 ;
        RECT 549.860 17.270 551.840 17.410 ;
        RECT 549.860 2.400 550.000 17.270 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 572.310 71.980 572.630 72.040 ;
        RECT 1380.530 71.980 1380.850 72.040 ;
        RECT 572.310 71.840 1380.850 71.980 ;
        RECT 572.310 71.780 572.630 71.840 ;
        RECT 1380.530 71.780 1380.850 71.840 ;
        RECT 567.710 14.860 568.030 14.920 ;
        RECT 572.310 14.860 572.630 14.920 ;
        RECT 567.710 14.720 572.630 14.860 ;
        RECT 567.710 14.660 568.030 14.720 ;
        RECT 572.310 14.660 572.630 14.720 ;
      LAYER via ;
        RECT 572.340 71.780 572.600 72.040 ;
        RECT 1380.560 71.780 1380.820 72.040 ;
        RECT 567.740 14.660 568.000 14.920 ;
        RECT 572.340 14.660 572.600 14.920 ;
      LAYER met2 ;
        RECT 1382.325 1700.410 1382.605 1704.000 ;
        RECT 1380.620 1700.270 1382.605 1700.410 ;
        RECT 1380.620 72.070 1380.760 1700.270 ;
        RECT 1382.325 1700.000 1382.605 1700.270 ;
        RECT 572.340 71.750 572.600 72.070 ;
        RECT 1380.560 71.750 1380.820 72.070 ;
        RECT 572.400 14.950 572.540 71.750 ;
        RECT 567.740 14.630 568.000 14.950 ;
        RECT 572.340 14.630 572.600 14.950 ;
        RECT 567.800 2.400 567.940 14.630 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 586.110 71.640 586.430 71.700 ;
        RECT 1388.350 71.640 1388.670 71.700 ;
        RECT 586.110 71.500 1388.670 71.640 ;
        RECT 586.110 71.440 586.430 71.500 ;
        RECT 1388.350 71.440 1388.670 71.500 ;
      LAYER via ;
        RECT 586.140 71.440 586.400 71.700 ;
        RECT 1388.380 71.440 1388.640 71.700 ;
      LAYER met2 ;
        RECT 1389.685 1700.410 1389.965 1704.000 ;
        RECT 1388.440 1700.270 1389.965 1700.410 ;
        RECT 1388.440 71.730 1388.580 1700.270 ;
        RECT 1389.685 1700.000 1389.965 1700.270 ;
        RECT 586.140 71.410 586.400 71.730 ;
        RECT 1388.380 71.410 1388.640 71.730 ;
        RECT 586.200 17.410 586.340 71.410 ;
        RECT 585.740 17.270 586.340 17.410 ;
        RECT 585.740 2.400 585.880 17.270 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1180.890 1678.480 1181.210 1678.540 ;
        RECT 1185.030 1678.480 1185.350 1678.540 ;
        RECT 1180.890 1678.340 1185.350 1678.480 ;
        RECT 1180.890 1678.280 1181.210 1678.340 ;
        RECT 1185.030 1678.280 1185.350 1678.340 ;
        RECT 91.610 45.120 91.930 45.180 ;
        RECT 1180.890 45.120 1181.210 45.180 ;
        RECT 91.610 44.980 1181.210 45.120 ;
        RECT 91.610 44.920 91.930 44.980 ;
        RECT 1180.890 44.920 1181.210 44.980 ;
      LAYER via ;
        RECT 1180.920 1678.280 1181.180 1678.540 ;
        RECT 1185.060 1678.280 1185.320 1678.540 ;
        RECT 91.640 44.920 91.900 45.180 ;
        RECT 1180.920 44.920 1181.180 45.180 ;
      LAYER met2 ;
        RECT 1186.365 1700.410 1186.645 1704.000 ;
        RECT 1185.120 1700.270 1186.645 1700.410 ;
        RECT 1185.120 1678.570 1185.260 1700.270 ;
        RECT 1186.365 1700.000 1186.645 1700.270 ;
        RECT 1180.920 1678.250 1181.180 1678.570 ;
        RECT 1185.060 1678.250 1185.320 1678.570 ;
        RECT 1180.980 45.210 1181.120 1678.250 ;
        RECT 91.640 44.890 91.900 45.210 ;
        RECT 1180.920 44.890 1181.180 45.210 ;
        RECT 91.700 2.400 91.840 44.890 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1394.405 241.485 1394.575 255.935 ;
      LAYER mcon ;
        RECT 1394.405 255.765 1394.575 255.935 ;
      LAYER met1 ;
        RECT 1394.330 1666.580 1394.650 1666.640 ;
        RECT 1395.250 1666.580 1395.570 1666.640 ;
        RECT 1394.330 1666.440 1395.570 1666.580 ;
        RECT 1394.330 1666.380 1394.650 1666.440 ;
        RECT 1395.250 1666.380 1395.570 1666.440 ;
        RECT 1394.330 835.280 1394.650 835.340 ;
        RECT 1393.960 835.140 1394.650 835.280 ;
        RECT 1393.960 834.660 1394.100 835.140 ;
        RECT 1394.330 835.080 1394.650 835.140 ;
        RECT 1393.870 834.400 1394.190 834.660 ;
        RECT 1394.330 593.680 1394.650 593.940 ;
        RECT 1394.420 593.260 1394.560 593.680 ;
        RECT 1394.330 593.000 1394.650 593.260 ;
        RECT 1394.330 400.560 1394.650 400.820 ;
        RECT 1394.420 400.140 1394.560 400.560 ;
        RECT 1394.330 399.880 1394.650 400.140 ;
        RECT 1394.330 255.920 1394.650 255.980 ;
        RECT 1394.135 255.780 1394.650 255.920 ;
        RECT 1394.330 255.720 1394.650 255.780 ;
        RECT 1394.330 241.640 1394.650 241.700 ;
        RECT 1394.135 241.500 1394.650 241.640 ;
        RECT 1394.330 241.440 1394.650 241.500 ;
        RECT 606.810 71.300 607.130 71.360 ;
        RECT 1393.870 71.300 1394.190 71.360 ;
        RECT 606.810 71.160 1394.190 71.300 ;
        RECT 606.810 71.100 607.130 71.160 ;
        RECT 1393.870 71.100 1394.190 71.160 ;
        RECT 603.130 14.860 603.450 14.920 ;
        RECT 606.810 14.860 607.130 14.920 ;
        RECT 603.130 14.720 607.130 14.860 ;
        RECT 603.130 14.660 603.450 14.720 ;
        RECT 606.810 14.660 607.130 14.720 ;
      LAYER via ;
        RECT 1394.360 1666.380 1394.620 1666.640 ;
        RECT 1395.280 1666.380 1395.540 1666.640 ;
        RECT 1394.360 835.080 1394.620 835.340 ;
        RECT 1393.900 834.400 1394.160 834.660 ;
        RECT 1394.360 593.680 1394.620 593.940 ;
        RECT 1394.360 593.000 1394.620 593.260 ;
        RECT 1394.360 400.560 1394.620 400.820 ;
        RECT 1394.360 399.880 1394.620 400.140 ;
        RECT 1394.360 255.720 1394.620 255.980 ;
        RECT 1394.360 241.440 1394.620 241.700 ;
        RECT 606.840 71.100 607.100 71.360 ;
        RECT 1393.900 71.100 1394.160 71.360 ;
        RECT 603.160 14.660 603.420 14.920 ;
        RECT 606.840 14.660 607.100 14.920 ;
      LAYER met2 ;
        RECT 1397.045 1700.410 1397.325 1704.000 ;
        RECT 1395.340 1700.270 1397.325 1700.410 ;
        RECT 1395.340 1666.670 1395.480 1700.270 ;
        RECT 1397.045 1700.000 1397.325 1700.270 ;
        RECT 1394.360 1666.350 1394.620 1666.670 ;
        RECT 1395.280 1666.350 1395.540 1666.670 ;
        RECT 1394.420 1511.370 1394.560 1666.350 ;
        RECT 1393.960 1511.230 1394.560 1511.370 ;
        RECT 1393.960 1510.690 1394.100 1511.230 ;
        RECT 1393.960 1510.550 1394.560 1510.690 ;
        RECT 1394.420 1414.810 1394.560 1510.550 ;
        RECT 1393.960 1414.670 1394.560 1414.810 ;
        RECT 1393.960 1414.130 1394.100 1414.670 ;
        RECT 1393.960 1413.990 1394.560 1414.130 ;
        RECT 1394.420 1318.250 1394.560 1413.990 ;
        RECT 1393.960 1318.110 1394.560 1318.250 ;
        RECT 1393.960 1317.570 1394.100 1318.110 ;
        RECT 1393.960 1317.430 1394.560 1317.570 ;
        RECT 1394.420 1221.690 1394.560 1317.430 ;
        RECT 1393.960 1221.550 1394.560 1221.690 ;
        RECT 1393.960 1221.010 1394.100 1221.550 ;
        RECT 1393.960 1220.870 1394.560 1221.010 ;
        RECT 1394.420 1125.130 1394.560 1220.870 ;
        RECT 1393.960 1124.990 1394.560 1125.130 ;
        RECT 1393.960 1124.450 1394.100 1124.990 ;
        RECT 1393.960 1124.310 1394.560 1124.450 ;
        RECT 1394.420 1028.570 1394.560 1124.310 ;
        RECT 1393.960 1028.430 1394.560 1028.570 ;
        RECT 1393.960 1027.890 1394.100 1028.430 ;
        RECT 1393.960 1027.750 1394.560 1027.890 ;
        RECT 1394.420 932.010 1394.560 1027.750 ;
        RECT 1393.960 931.870 1394.560 932.010 ;
        RECT 1393.960 931.330 1394.100 931.870 ;
        RECT 1393.960 931.190 1394.560 931.330 ;
        RECT 1394.420 835.370 1394.560 931.190 ;
        RECT 1394.360 835.050 1394.620 835.370 ;
        RECT 1393.900 834.370 1394.160 834.690 ;
        RECT 1393.960 700.130 1394.100 834.370 ;
        RECT 1393.960 699.990 1394.560 700.130 ;
        RECT 1394.420 593.970 1394.560 699.990 ;
        RECT 1394.360 593.650 1394.620 593.970 ;
        RECT 1394.360 592.970 1394.620 593.290 ;
        RECT 1394.420 400.850 1394.560 592.970 ;
        RECT 1394.360 400.530 1394.620 400.850 ;
        RECT 1394.360 399.850 1394.620 400.170 ;
        RECT 1394.420 256.010 1394.560 399.850 ;
        RECT 1394.360 255.690 1394.620 256.010 ;
        RECT 1394.360 241.410 1394.620 241.730 ;
        RECT 1394.420 158.850 1394.560 241.410 ;
        RECT 1393.960 158.710 1394.560 158.850 ;
        RECT 1393.960 71.390 1394.100 158.710 ;
        RECT 606.840 71.070 607.100 71.390 ;
        RECT 1393.900 71.070 1394.160 71.390 ;
        RECT 606.900 14.950 607.040 71.070 ;
        RECT 603.160 14.630 603.420 14.950 ;
        RECT 606.840 14.630 607.100 14.950 ;
        RECT 603.220 2.400 603.360 14.630 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1401.230 1678.140 1401.550 1678.200 ;
        RECT 1403.070 1678.140 1403.390 1678.200 ;
        RECT 1401.230 1678.000 1403.390 1678.140 ;
        RECT 1401.230 1677.940 1401.550 1678.000 ;
        RECT 1403.070 1677.940 1403.390 1678.000 ;
        RECT 627.050 70.960 627.370 71.020 ;
        RECT 1401.230 70.960 1401.550 71.020 ;
        RECT 627.050 70.820 1401.550 70.960 ;
        RECT 627.050 70.760 627.370 70.820 ;
        RECT 1401.230 70.760 1401.550 70.820 ;
        RECT 621.070 20.980 621.390 21.040 ;
        RECT 627.050 20.980 627.370 21.040 ;
        RECT 621.070 20.840 627.370 20.980 ;
        RECT 621.070 20.780 621.390 20.840 ;
        RECT 627.050 20.780 627.370 20.840 ;
      LAYER via ;
        RECT 1401.260 1677.940 1401.520 1678.200 ;
        RECT 1403.100 1677.940 1403.360 1678.200 ;
        RECT 627.080 70.760 627.340 71.020 ;
        RECT 1401.260 70.760 1401.520 71.020 ;
        RECT 621.100 20.780 621.360 21.040 ;
        RECT 627.080 20.780 627.340 21.040 ;
      LAYER met2 ;
        RECT 1404.405 1700.410 1404.685 1704.000 ;
        RECT 1403.160 1700.270 1404.685 1700.410 ;
        RECT 1403.160 1678.230 1403.300 1700.270 ;
        RECT 1404.405 1700.000 1404.685 1700.270 ;
        RECT 1401.260 1677.910 1401.520 1678.230 ;
        RECT 1403.100 1677.910 1403.360 1678.230 ;
        RECT 1401.320 71.050 1401.460 1677.910 ;
        RECT 627.080 70.730 627.340 71.050 ;
        RECT 1401.260 70.730 1401.520 71.050 ;
        RECT 627.140 21.070 627.280 70.730 ;
        RECT 621.100 20.750 621.360 21.070 ;
        RECT 627.080 20.750 627.340 21.070 ;
        RECT 621.160 2.400 621.300 20.750 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 116.910 58.720 117.230 58.780 ;
        RECT 1194.690 58.720 1195.010 58.780 ;
        RECT 116.910 58.580 1195.010 58.720 ;
        RECT 116.910 58.520 117.230 58.580 ;
        RECT 1194.690 58.520 1195.010 58.580 ;
        RECT 115.530 2.960 115.850 3.020 ;
        RECT 116.910 2.960 117.230 3.020 ;
        RECT 115.530 2.820 117.230 2.960 ;
        RECT 115.530 2.760 115.850 2.820 ;
        RECT 116.910 2.760 117.230 2.820 ;
      LAYER via ;
        RECT 116.940 58.520 117.200 58.780 ;
        RECT 1194.720 58.520 1194.980 58.780 ;
        RECT 115.560 2.760 115.820 3.020 ;
        RECT 116.940 2.760 117.200 3.020 ;
      LAYER met2 ;
        RECT 1196.485 1700.410 1196.765 1704.000 ;
        RECT 1194.780 1700.270 1196.765 1700.410 ;
        RECT 1194.780 58.810 1194.920 1700.270 ;
        RECT 1196.485 1700.000 1196.765 1700.270 ;
        RECT 116.940 58.490 117.200 58.810 ;
        RECT 1194.720 58.490 1194.980 58.810 ;
        RECT 117.000 3.050 117.140 58.490 ;
        RECT 115.560 2.730 115.820 3.050 ;
        RECT 116.940 2.730 117.200 3.050 ;
        RECT 115.620 2.400 115.760 2.730 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1169.390 1686.980 1169.710 1687.040 ;
        RECT 1206.190 1686.980 1206.510 1687.040 ;
        RECT 1169.390 1686.840 1206.510 1686.980 ;
        RECT 1169.390 1686.780 1169.710 1686.840 ;
        RECT 1206.190 1686.780 1206.510 1686.840 ;
        RECT 139.450 45.460 139.770 45.520 ;
        RECT 1169.390 45.460 1169.710 45.520 ;
        RECT 139.450 45.320 1169.710 45.460 ;
        RECT 139.450 45.260 139.770 45.320 ;
        RECT 1169.390 45.260 1169.710 45.320 ;
      LAYER via ;
        RECT 1169.420 1686.780 1169.680 1687.040 ;
        RECT 1206.220 1686.780 1206.480 1687.040 ;
        RECT 139.480 45.260 139.740 45.520 ;
        RECT 1169.420 45.260 1169.680 45.520 ;
      LAYER met2 ;
        RECT 1206.145 1700.000 1206.425 1704.000 ;
        RECT 1206.280 1687.070 1206.420 1700.000 ;
        RECT 1169.420 1686.750 1169.680 1687.070 ;
        RECT 1206.220 1686.750 1206.480 1687.070 ;
        RECT 1169.480 45.550 1169.620 1686.750 ;
        RECT 139.480 45.230 139.740 45.550 ;
        RECT 1169.420 45.230 1169.680 45.550 ;
        RECT 139.540 2.400 139.680 45.230 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1208.030 1678.140 1208.350 1678.200 ;
        RECT 1211.710 1678.140 1212.030 1678.200 ;
        RECT 1208.030 1678.000 1212.030 1678.140 ;
        RECT 1208.030 1677.940 1208.350 1678.000 ;
        RECT 1211.710 1677.940 1212.030 1678.000 ;
        RECT 158.310 65.520 158.630 65.580 ;
        RECT 1208.030 65.520 1208.350 65.580 ;
        RECT 158.310 65.380 1208.350 65.520 ;
        RECT 158.310 65.320 158.630 65.380 ;
        RECT 1208.030 65.320 1208.350 65.380 ;
      LAYER via ;
        RECT 1208.060 1677.940 1208.320 1678.200 ;
        RECT 1211.740 1677.940 1212.000 1678.200 ;
        RECT 158.340 65.320 158.600 65.580 ;
        RECT 1208.060 65.320 1208.320 65.580 ;
      LAYER met2 ;
        RECT 1213.505 1700.410 1213.785 1704.000 ;
        RECT 1211.800 1700.270 1213.785 1700.410 ;
        RECT 1211.800 1678.230 1211.940 1700.270 ;
        RECT 1213.505 1700.000 1213.785 1700.270 ;
        RECT 1208.060 1677.910 1208.320 1678.230 ;
        RECT 1211.740 1677.910 1212.000 1678.230 ;
        RECT 1208.120 65.610 1208.260 1677.910 ;
        RECT 158.340 65.290 158.600 65.610 ;
        RECT 1208.060 65.290 1208.320 65.610 ;
        RECT 158.400 3.130 158.540 65.290 ;
        RECT 157.480 2.990 158.540 3.130 ;
        RECT 157.480 2.400 157.620 2.990 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 286.190 1689.020 286.510 1689.080 ;
        RECT 1220.910 1689.020 1221.230 1689.080 ;
        RECT 286.190 1688.880 1221.230 1689.020 ;
        RECT 286.190 1688.820 286.510 1688.880 ;
        RECT 1220.910 1688.820 1221.230 1688.880 ;
        RECT 174.870 16.900 175.190 16.960 ;
        RECT 286.190 16.900 286.510 16.960 ;
        RECT 174.870 16.760 286.510 16.900 ;
        RECT 174.870 16.700 175.190 16.760 ;
        RECT 286.190 16.700 286.510 16.760 ;
      LAYER via ;
        RECT 286.220 1688.820 286.480 1689.080 ;
        RECT 1220.940 1688.820 1221.200 1689.080 ;
        RECT 174.900 16.700 175.160 16.960 ;
        RECT 286.220 16.700 286.480 16.960 ;
      LAYER met2 ;
        RECT 1220.865 1700.000 1221.145 1704.000 ;
        RECT 1221.000 1689.110 1221.140 1700.000 ;
        RECT 286.220 1688.790 286.480 1689.110 ;
        RECT 1220.940 1688.790 1221.200 1689.110 ;
        RECT 286.280 16.990 286.420 1688.790 ;
        RECT 174.900 16.670 175.160 16.990 ;
        RECT 286.220 16.670 286.480 16.990 ;
        RECT 174.960 2.400 175.100 16.670 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1228.270 904.100 1228.590 904.360 ;
        RECT 1228.360 903.680 1228.500 904.100 ;
        RECT 1228.270 903.420 1228.590 903.680 ;
        RECT 192.810 18.940 193.130 19.000 ;
        RECT 1228.270 18.940 1228.590 19.000 ;
        RECT 192.810 18.800 1228.590 18.940 ;
        RECT 192.810 18.740 193.130 18.800 ;
        RECT 1228.270 18.740 1228.590 18.800 ;
      LAYER via ;
        RECT 1228.300 904.100 1228.560 904.360 ;
        RECT 1228.300 903.420 1228.560 903.680 ;
        RECT 192.840 18.740 193.100 19.000 ;
        RECT 1228.300 18.740 1228.560 19.000 ;
      LAYER met2 ;
        RECT 1228.225 1700.000 1228.505 1704.000 ;
        RECT 1228.360 904.390 1228.500 1700.000 ;
        RECT 1228.300 904.070 1228.560 904.390 ;
        RECT 1228.300 903.390 1228.560 903.710 ;
        RECT 1228.360 19.030 1228.500 903.390 ;
        RECT 192.840 18.710 193.100 19.030 ;
        RECT 1228.300 18.710 1228.560 19.030 ;
        RECT 192.900 2.400 193.040 18.710 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 334.490 1689.700 334.810 1689.760 ;
        RECT 1235.630 1689.700 1235.950 1689.760 ;
        RECT 334.490 1689.560 1235.950 1689.700 ;
        RECT 334.490 1689.500 334.810 1689.560 ;
        RECT 1235.630 1689.500 1235.950 1689.560 ;
        RECT 210.750 16.560 211.070 16.620 ;
        RECT 334.490 16.560 334.810 16.620 ;
        RECT 210.750 16.420 334.810 16.560 ;
        RECT 210.750 16.360 211.070 16.420 ;
        RECT 334.490 16.360 334.810 16.420 ;
      LAYER via ;
        RECT 334.520 1689.500 334.780 1689.760 ;
        RECT 1235.660 1689.500 1235.920 1689.760 ;
        RECT 210.780 16.360 211.040 16.620 ;
        RECT 334.520 16.360 334.780 16.620 ;
      LAYER met2 ;
        RECT 1235.585 1700.000 1235.865 1704.000 ;
        RECT 1235.720 1689.790 1235.860 1700.000 ;
        RECT 334.520 1689.470 334.780 1689.790 ;
        RECT 1235.660 1689.470 1235.920 1689.790 ;
        RECT 334.580 16.650 334.720 1689.470 ;
        RECT 210.780 16.330 211.040 16.650 ;
        RECT 334.520 16.330 334.780 16.650 ;
        RECT 210.840 2.400 210.980 16.330 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1238.390 1686.980 1238.710 1687.040 ;
        RECT 1242.990 1686.980 1243.310 1687.040 ;
        RECT 1238.390 1686.840 1243.310 1686.980 ;
        RECT 1238.390 1686.780 1238.710 1686.840 ;
        RECT 1242.990 1686.780 1243.310 1686.840 ;
        RECT 228.690 19.620 229.010 19.680 ;
        RECT 1238.390 19.620 1238.710 19.680 ;
        RECT 228.690 19.480 1238.710 19.620 ;
        RECT 228.690 19.420 229.010 19.480 ;
        RECT 1238.390 19.420 1238.710 19.480 ;
      LAYER via ;
        RECT 1238.420 1686.780 1238.680 1687.040 ;
        RECT 1243.020 1686.780 1243.280 1687.040 ;
        RECT 228.720 19.420 228.980 19.680 ;
        RECT 1238.420 19.420 1238.680 19.680 ;
      LAYER met2 ;
        RECT 1242.945 1700.000 1243.225 1704.000 ;
        RECT 1243.080 1687.070 1243.220 1700.000 ;
        RECT 1238.420 1686.750 1238.680 1687.070 ;
        RECT 1243.020 1686.750 1243.280 1687.070 ;
        RECT 1238.480 19.710 1238.620 1686.750 ;
        RECT 228.720 19.390 228.980 19.710 ;
        RECT 1238.420 19.390 1238.680 19.710 ;
        RECT 228.780 2.400 228.920 19.390 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 65.390 1686.980 65.710 1687.040 ;
        RECT 1167.550 1686.980 1167.870 1687.040 ;
        RECT 65.390 1686.840 1167.870 1686.980 ;
        RECT 65.390 1686.780 65.710 1686.840 ;
        RECT 1167.550 1686.780 1167.870 1686.840 ;
        RECT 50.210 16.560 50.530 16.620 ;
        RECT 65.390 16.560 65.710 16.620 ;
        RECT 50.210 16.420 65.710 16.560 ;
        RECT 50.210 16.360 50.530 16.420 ;
        RECT 65.390 16.360 65.710 16.420 ;
      LAYER via ;
        RECT 65.420 1686.780 65.680 1687.040 ;
        RECT 1167.580 1686.780 1167.840 1687.040 ;
        RECT 50.240 16.360 50.500 16.620 ;
        RECT 65.420 16.360 65.680 16.620 ;
      LAYER met2 ;
        RECT 1169.345 1700.410 1169.625 1704.000 ;
        RECT 1167.640 1700.270 1169.625 1700.410 ;
        RECT 1167.640 1687.070 1167.780 1700.270 ;
        RECT 1169.345 1700.000 1169.625 1700.270 ;
        RECT 65.420 1686.750 65.680 1687.070 ;
        RECT 1167.580 1686.750 1167.840 1687.070 ;
        RECT 65.480 16.650 65.620 1686.750 ;
        RECT 50.240 16.330 50.500 16.650 ;
        RECT 65.420 16.330 65.680 16.650 ;
        RECT 50.300 2.400 50.440 16.330 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1245.290 1686.980 1245.610 1687.040 ;
        RECT 1252.650 1686.980 1252.970 1687.040 ;
        RECT 1245.290 1686.840 1252.970 1686.980 ;
        RECT 1245.290 1686.780 1245.610 1686.840 ;
        RECT 1252.650 1686.780 1252.970 1686.840 ;
        RECT 252.610 20.300 252.930 20.360 ;
        RECT 1245.290 20.300 1245.610 20.360 ;
        RECT 252.610 20.160 1245.610 20.300 ;
        RECT 252.610 20.100 252.930 20.160 ;
        RECT 1245.290 20.100 1245.610 20.160 ;
      LAYER via ;
        RECT 1245.320 1686.780 1245.580 1687.040 ;
        RECT 1252.680 1686.780 1252.940 1687.040 ;
        RECT 252.640 20.100 252.900 20.360 ;
        RECT 1245.320 20.100 1245.580 20.360 ;
      LAYER met2 ;
        RECT 1252.605 1700.000 1252.885 1704.000 ;
        RECT 1252.740 1687.070 1252.880 1700.000 ;
        RECT 1245.320 1686.750 1245.580 1687.070 ;
        RECT 1252.680 1686.750 1252.940 1687.070 ;
        RECT 1245.380 20.390 1245.520 1686.750 ;
        RECT 252.640 20.070 252.900 20.390 ;
        RECT 1245.320 20.070 1245.580 20.390 ;
        RECT 252.700 2.400 252.840 20.070 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 355.190 1690.040 355.510 1690.100 ;
        RECT 1260.010 1690.040 1260.330 1690.100 ;
        RECT 355.190 1689.900 1260.330 1690.040 ;
        RECT 355.190 1689.840 355.510 1689.900 ;
        RECT 1260.010 1689.840 1260.330 1689.900 ;
        RECT 270.090 15.880 270.410 15.940 ;
        RECT 355.190 15.880 355.510 15.940 ;
        RECT 270.090 15.740 355.510 15.880 ;
        RECT 270.090 15.680 270.410 15.740 ;
        RECT 355.190 15.680 355.510 15.740 ;
      LAYER via ;
        RECT 355.220 1689.840 355.480 1690.100 ;
        RECT 1260.040 1689.840 1260.300 1690.100 ;
        RECT 270.120 15.680 270.380 15.940 ;
        RECT 355.220 15.680 355.480 15.940 ;
      LAYER met2 ;
        RECT 1259.965 1700.000 1260.245 1704.000 ;
        RECT 1260.100 1690.130 1260.240 1700.000 ;
        RECT 355.220 1689.810 355.480 1690.130 ;
        RECT 1260.040 1689.810 1260.300 1690.130 ;
        RECT 355.280 15.970 355.420 1689.810 ;
        RECT 270.120 15.650 270.380 15.970 ;
        RECT 355.220 15.650 355.480 15.970 ;
        RECT 270.180 2.400 270.320 15.650 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1253.570 1686.980 1253.890 1687.040 ;
        RECT 1267.370 1686.980 1267.690 1687.040 ;
        RECT 1253.570 1686.840 1267.690 1686.980 ;
        RECT 1253.570 1686.780 1253.890 1686.840 ;
        RECT 1267.370 1686.780 1267.690 1686.840 ;
        RECT 288.030 20.640 288.350 20.700 ;
        RECT 1252.190 20.640 1252.510 20.700 ;
        RECT 288.030 20.500 1252.510 20.640 ;
        RECT 288.030 20.440 288.350 20.500 ;
        RECT 1252.190 20.440 1252.510 20.500 ;
      LAYER via ;
        RECT 1253.600 1686.780 1253.860 1687.040 ;
        RECT 1267.400 1686.780 1267.660 1687.040 ;
        RECT 288.060 20.440 288.320 20.700 ;
        RECT 1252.220 20.440 1252.480 20.700 ;
      LAYER met2 ;
        RECT 1267.325 1700.000 1267.605 1704.000 ;
        RECT 1267.460 1687.070 1267.600 1700.000 ;
        RECT 1253.600 1686.750 1253.860 1687.070 ;
        RECT 1267.400 1686.750 1267.660 1687.070 ;
        RECT 1253.660 1677.290 1253.800 1686.750 ;
        RECT 1252.280 1677.150 1253.800 1677.290 ;
        RECT 1252.280 20.730 1252.420 1677.150 ;
        RECT 288.060 20.410 288.320 20.730 ;
        RECT 1252.220 20.410 1252.480 20.730 ;
        RECT 288.120 2.400 288.260 20.410 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 496.945 1684.105 497.115 1685.635 ;
        RECT 544.785 1684.105 544.955 1686.315 ;
        RECT 565.945 1683.765 566.115 1686.315 ;
        RECT 613.785 1683.765 613.955 1686.315 ;
      LAYER mcon ;
        RECT 544.785 1686.145 544.955 1686.315 ;
        RECT 496.945 1685.465 497.115 1685.635 ;
        RECT 565.945 1686.145 566.115 1686.315 ;
        RECT 613.785 1686.145 613.955 1686.315 ;
      LAYER met1 ;
        RECT 389.690 1686.640 390.010 1686.700 ;
        RECT 389.690 1686.500 423.500 1686.640 ;
        RECT 389.690 1686.440 390.010 1686.500 ;
        RECT 423.360 1685.960 423.500 1686.500 ;
        RECT 544.725 1686.300 545.015 1686.345 ;
        RECT 565.885 1686.300 566.175 1686.345 ;
        RECT 544.725 1686.160 566.175 1686.300 ;
        RECT 544.725 1686.115 545.015 1686.160 ;
        RECT 565.885 1686.115 566.175 1686.160 ;
        RECT 613.725 1686.300 614.015 1686.345 ;
        RECT 662.470 1686.300 662.790 1686.360 ;
        RECT 613.725 1686.160 662.790 1686.300 ;
        RECT 613.725 1686.115 614.015 1686.160 ;
        RECT 662.470 1686.100 662.790 1686.160 ;
        RECT 710.310 1686.300 710.630 1686.360 ;
        RECT 759.070 1686.300 759.390 1686.360 ;
        RECT 710.310 1686.160 759.390 1686.300 ;
        RECT 710.310 1686.100 710.630 1686.160 ;
        RECT 759.070 1686.100 759.390 1686.160 ;
        RECT 806.910 1686.300 807.230 1686.360 ;
        RECT 855.670 1686.300 855.990 1686.360 ;
        RECT 806.910 1686.160 855.990 1686.300 ;
        RECT 806.910 1686.100 807.230 1686.160 ;
        RECT 855.670 1686.100 855.990 1686.160 ;
        RECT 903.510 1686.300 903.830 1686.360 ;
        RECT 952.270 1686.300 952.590 1686.360 ;
        RECT 903.510 1686.160 952.590 1686.300 ;
        RECT 903.510 1686.100 903.830 1686.160 ;
        RECT 952.270 1686.100 952.590 1686.160 ;
        RECT 1000.110 1686.300 1000.430 1686.360 ;
        RECT 1048.870 1686.300 1049.190 1686.360 ;
        RECT 1000.110 1686.160 1049.190 1686.300 ;
        RECT 1000.110 1686.100 1000.430 1686.160 ;
        RECT 1048.870 1686.100 1049.190 1686.160 ;
        RECT 1096.710 1686.300 1097.030 1686.360 ;
        RECT 1145.930 1686.300 1146.250 1686.360 ;
        RECT 1096.710 1686.160 1146.250 1686.300 ;
        RECT 1096.710 1686.100 1097.030 1686.160 ;
        RECT 1145.930 1686.100 1146.250 1686.160 ;
        RECT 1173.070 1686.300 1173.390 1686.360 ;
        RECT 1274.730 1686.300 1275.050 1686.360 ;
        RECT 1173.070 1686.160 1275.050 1686.300 ;
        RECT 1173.070 1686.100 1173.390 1686.160 ;
        RECT 1274.730 1686.100 1275.050 1686.160 ;
        RECT 423.360 1685.820 472.720 1685.960 ;
        RECT 472.580 1685.620 472.720 1685.820 ;
        RECT 496.885 1685.620 497.175 1685.665 ;
        RECT 472.580 1685.480 497.175 1685.620 ;
        RECT 496.885 1685.435 497.175 1685.480 ;
        RECT 496.885 1684.260 497.175 1684.305 ;
        RECT 544.725 1684.260 545.015 1684.305 ;
        RECT 496.885 1684.120 545.015 1684.260 ;
        RECT 496.885 1684.075 497.175 1684.120 ;
        RECT 544.725 1684.075 545.015 1684.120 ;
        RECT 565.885 1683.920 566.175 1683.965 ;
        RECT 613.725 1683.920 614.015 1683.965 ;
        RECT 565.885 1683.780 614.015 1683.920 ;
        RECT 565.885 1683.735 566.175 1683.780 ;
        RECT 613.725 1683.735 614.015 1683.780 ;
        RECT 305.970 15.540 306.290 15.600 ;
        RECT 389.690 15.540 390.010 15.600 ;
        RECT 305.970 15.400 390.010 15.540 ;
        RECT 305.970 15.340 306.290 15.400 ;
        RECT 389.690 15.340 390.010 15.400 ;
      LAYER via ;
        RECT 389.720 1686.440 389.980 1686.700 ;
        RECT 662.500 1686.100 662.760 1686.360 ;
        RECT 710.340 1686.100 710.600 1686.360 ;
        RECT 759.100 1686.100 759.360 1686.360 ;
        RECT 806.940 1686.100 807.200 1686.360 ;
        RECT 855.700 1686.100 855.960 1686.360 ;
        RECT 903.540 1686.100 903.800 1686.360 ;
        RECT 952.300 1686.100 952.560 1686.360 ;
        RECT 1000.140 1686.100 1000.400 1686.360 ;
        RECT 1048.900 1686.100 1049.160 1686.360 ;
        RECT 1096.740 1686.100 1097.000 1686.360 ;
        RECT 1145.960 1686.100 1146.220 1686.360 ;
        RECT 1173.100 1686.100 1173.360 1686.360 ;
        RECT 1274.760 1686.100 1275.020 1686.360 ;
        RECT 306.000 15.340 306.260 15.600 ;
        RECT 389.720 15.340 389.980 15.600 ;
      LAYER met2 ;
        RECT 1274.685 1700.000 1274.965 1704.000 ;
        RECT 389.720 1686.410 389.980 1686.730 ;
        RECT 389.780 15.630 389.920 1686.410 ;
        RECT 1274.820 1686.390 1274.960 1700.000 ;
        RECT 662.500 1686.245 662.760 1686.390 ;
        RECT 710.340 1686.245 710.600 1686.390 ;
        RECT 759.100 1686.245 759.360 1686.390 ;
        RECT 806.940 1686.245 807.200 1686.390 ;
        RECT 855.700 1686.245 855.960 1686.390 ;
        RECT 903.540 1686.245 903.800 1686.390 ;
        RECT 952.300 1686.245 952.560 1686.390 ;
        RECT 1000.140 1686.245 1000.400 1686.390 ;
        RECT 1048.900 1686.245 1049.160 1686.390 ;
        RECT 1096.740 1686.245 1097.000 1686.390 ;
        RECT 1145.960 1686.245 1146.220 1686.390 ;
        RECT 1173.100 1686.245 1173.360 1686.390 ;
        RECT 662.490 1685.875 662.770 1686.245 ;
        RECT 710.330 1685.875 710.610 1686.245 ;
        RECT 759.090 1685.875 759.370 1686.245 ;
        RECT 806.930 1685.875 807.210 1686.245 ;
        RECT 855.690 1685.875 855.970 1686.245 ;
        RECT 903.530 1685.875 903.810 1686.245 ;
        RECT 952.290 1685.875 952.570 1686.245 ;
        RECT 1000.130 1685.875 1000.410 1686.245 ;
        RECT 1048.890 1685.875 1049.170 1686.245 ;
        RECT 1096.730 1685.875 1097.010 1686.245 ;
        RECT 1145.950 1685.875 1146.230 1686.245 ;
        RECT 1173.090 1685.875 1173.370 1686.245 ;
        RECT 1274.760 1686.070 1275.020 1686.390 ;
        RECT 306.000 15.310 306.260 15.630 ;
        RECT 389.720 15.310 389.980 15.630 ;
        RECT 306.060 2.400 306.200 15.310 ;
        RECT 305.850 -4.800 306.410 2.400 ;
      LAYER via2 ;
        RECT 662.490 1685.920 662.770 1686.200 ;
        RECT 710.330 1685.920 710.610 1686.200 ;
        RECT 759.090 1685.920 759.370 1686.200 ;
        RECT 806.930 1685.920 807.210 1686.200 ;
        RECT 855.690 1685.920 855.970 1686.200 ;
        RECT 903.530 1685.920 903.810 1686.200 ;
        RECT 952.290 1685.920 952.570 1686.200 ;
        RECT 1000.130 1685.920 1000.410 1686.200 ;
        RECT 1048.890 1685.920 1049.170 1686.200 ;
        RECT 1096.730 1685.920 1097.010 1686.200 ;
        RECT 1145.950 1685.920 1146.230 1686.200 ;
        RECT 1173.090 1685.920 1173.370 1686.200 ;
      LAYER met3 ;
        RECT 662.465 1686.210 662.795 1686.225 ;
        RECT 710.305 1686.210 710.635 1686.225 ;
        RECT 662.465 1685.910 710.635 1686.210 ;
        RECT 662.465 1685.895 662.795 1685.910 ;
        RECT 710.305 1685.895 710.635 1685.910 ;
        RECT 759.065 1686.210 759.395 1686.225 ;
        RECT 806.905 1686.210 807.235 1686.225 ;
        RECT 759.065 1685.910 807.235 1686.210 ;
        RECT 759.065 1685.895 759.395 1685.910 ;
        RECT 806.905 1685.895 807.235 1685.910 ;
        RECT 855.665 1686.210 855.995 1686.225 ;
        RECT 903.505 1686.210 903.835 1686.225 ;
        RECT 855.665 1685.910 903.835 1686.210 ;
        RECT 855.665 1685.895 855.995 1685.910 ;
        RECT 903.505 1685.895 903.835 1685.910 ;
        RECT 952.265 1686.210 952.595 1686.225 ;
        RECT 1000.105 1686.210 1000.435 1686.225 ;
        RECT 952.265 1685.910 1000.435 1686.210 ;
        RECT 952.265 1685.895 952.595 1685.910 ;
        RECT 1000.105 1685.895 1000.435 1685.910 ;
        RECT 1048.865 1686.210 1049.195 1686.225 ;
        RECT 1096.705 1686.210 1097.035 1686.225 ;
        RECT 1048.865 1685.910 1097.035 1686.210 ;
        RECT 1048.865 1685.895 1049.195 1685.910 ;
        RECT 1096.705 1685.895 1097.035 1685.910 ;
        RECT 1145.925 1686.210 1146.255 1686.225 ;
        RECT 1173.065 1686.210 1173.395 1686.225 ;
        RECT 1145.925 1685.910 1173.395 1686.210 ;
        RECT 1145.925 1685.895 1146.255 1685.910 ;
        RECT 1173.065 1685.895 1173.395 1685.910 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1260.930 1688.000 1261.250 1688.060 ;
        RECT 1282.090 1688.000 1282.410 1688.060 ;
        RECT 1260.930 1687.860 1282.410 1688.000 ;
        RECT 1260.930 1687.800 1261.250 1687.860 ;
        RECT 1282.090 1687.800 1282.410 1687.860 ;
        RECT 323.450 16.900 323.770 16.960 ;
        RECT 1259.090 16.900 1259.410 16.960 ;
        RECT 323.450 16.760 1259.410 16.900 ;
        RECT 323.450 16.700 323.770 16.760 ;
        RECT 1259.090 16.700 1259.410 16.760 ;
      LAYER via ;
        RECT 1260.960 1687.800 1261.220 1688.060 ;
        RECT 1282.120 1687.800 1282.380 1688.060 ;
        RECT 323.480 16.700 323.740 16.960 ;
        RECT 1259.120 16.700 1259.380 16.960 ;
      LAYER met2 ;
        RECT 1282.045 1700.000 1282.325 1704.000 ;
        RECT 1282.180 1688.090 1282.320 1700.000 ;
        RECT 1260.960 1687.770 1261.220 1688.090 ;
        RECT 1282.120 1687.770 1282.380 1688.090 ;
        RECT 1261.020 1671.850 1261.160 1687.770 ;
        RECT 1259.180 1671.710 1261.160 1671.850 ;
        RECT 1259.180 16.990 1259.320 1671.710 ;
        RECT 323.480 16.670 323.740 16.990 ;
        RECT 1259.120 16.670 1259.380 16.990 ;
        RECT 323.540 8.570 323.680 16.670 ;
        RECT 323.540 8.430 324.140 8.570 ;
        RECT 324.000 2.400 324.140 8.430 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 396.590 1690.380 396.910 1690.440 ;
        RECT 1289.450 1690.380 1289.770 1690.440 ;
        RECT 396.590 1690.240 1289.770 1690.380 ;
        RECT 396.590 1690.180 396.910 1690.240 ;
        RECT 1289.450 1690.180 1289.770 1690.240 ;
        RECT 341.390 15.200 341.710 15.260 ;
        RECT 341.390 15.060 372.900 15.200 ;
        RECT 341.390 15.000 341.710 15.060 ;
        RECT 372.760 14.520 372.900 15.060 ;
        RECT 396.590 14.520 396.910 14.580 ;
        RECT 372.760 14.380 396.910 14.520 ;
        RECT 396.590 14.320 396.910 14.380 ;
      LAYER via ;
        RECT 396.620 1690.180 396.880 1690.440 ;
        RECT 1289.480 1690.180 1289.740 1690.440 ;
        RECT 341.420 15.000 341.680 15.260 ;
        RECT 396.620 14.320 396.880 14.580 ;
      LAYER met2 ;
        RECT 1289.405 1700.000 1289.685 1704.000 ;
        RECT 1289.540 1690.470 1289.680 1700.000 ;
        RECT 396.620 1690.150 396.880 1690.470 ;
        RECT 1289.480 1690.150 1289.740 1690.470 ;
        RECT 341.420 14.970 341.680 15.290 ;
        RECT 341.480 2.400 341.620 14.970 ;
        RECT 396.680 14.610 396.820 1690.150 ;
        RECT 396.620 14.290 396.880 14.610 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1265.990 1687.660 1266.310 1687.720 ;
        RECT 1296.810 1687.660 1297.130 1687.720 ;
        RECT 1265.990 1687.520 1297.130 1687.660 ;
        RECT 1265.990 1687.460 1266.310 1687.520 ;
        RECT 1296.810 1687.460 1297.130 1687.520 ;
        RECT 359.330 16.560 359.650 16.620 ;
        RECT 1265.990 16.560 1266.310 16.620 ;
        RECT 359.330 16.420 1266.310 16.560 ;
        RECT 359.330 16.360 359.650 16.420 ;
        RECT 1265.990 16.360 1266.310 16.420 ;
      LAYER via ;
        RECT 1266.020 1687.460 1266.280 1687.720 ;
        RECT 1296.840 1687.460 1297.100 1687.720 ;
        RECT 359.360 16.360 359.620 16.620 ;
        RECT 1266.020 16.360 1266.280 16.620 ;
      LAYER met2 ;
        RECT 1296.765 1700.000 1297.045 1704.000 ;
        RECT 1296.900 1687.750 1297.040 1700.000 ;
        RECT 1266.020 1687.430 1266.280 1687.750 ;
        RECT 1296.840 1687.430 1297.100 1687.750 ;
        RECT 1266.080 16.650 1266.220 1687.430 ;
        RECT 359.360 16.330 359.620 16.650 ;
        RECT 1266.020 16.330 1266.280 16.650 ;
        RECT 359.420 2.400 359.560 16.330 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 414.145 15.045 414.315 16.235 ;
      LAYER mcon ;
        RECT 414.145 16.065 414.315 16.235 ;
      LAYER met1 ;
        RECT 424.190 1686.640 424.510 1686.700 ;
        RECT 1304.170 1686.640 1304.490 1686.700 ;
        RECT 424.190 1686.500 1304.490 1686.640 ;
        RECT 424.190 1686.440 424.510 1686.500 ;
        RECT 1304.170 1686.440 1304.490 1686.500 ;
        RECT 414.085 16.220 414.375 16.265 ;
        RECT 424.190 16.220 424.510 16.280 ;
        RECT 414.085 16.080 424.510 16.220 ;
        RECT 414.085 16.035 414.375 16.080 ;
        RECT 424.190 16.020 424.510 16.080 ;
        RECT 377.270 15.200 377.590 15.260 ;
        RECT 414.085 15.200 414.375 15.245 ;
        RECT 377.270 15.060 414.375 15.200 ;
        RECT 377.270 15.000 377.590 15.060 ;
        RECT 414.085 15.015 414.375 15.060 ;
      LAYER via ;
        RECT 424.220 1686.440 424.480 1686.700 ;
        RECT 1304.200 1686.440 1304.460 1686.700 ;
        RECT 424.220 16.020 424.480 16.280 ;
        RECT 377.300 15.000 377.560 15.260 ;
      LAYER met2 ;
        RECT 1304.125 1700.000 1304.405 1704.000 ;
        RECT 1304.260 1686.730 1304.400 1700.000 ;
        RECT 424.220 1686.410 424.480 1686.730 ;
        RECT 1304.200 1686.410 1304.460 1686.730 ;
        RECT 424.280 16.310 424.420 1686.410 ;
        RECT 424.220 15.990 424.480 16.310 ;
        RECT 377.300 14.970 377.560 15.290 ;
        RECT 377.360 2.400 377.500 14.970 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1272.890 1688.680 1273.210 1688.740 ;
        RECT 1311.530 1688.680 1311.850 1688.740 ;
        RECT 1272.890 1688.540 1311.850 1688.680 ;
        RECT 1272.890 1688.480 1273.210 1688.540 ;
        RECT 1311.530 1688.480 1311.850 1688.540 ;
        RECT 1272.890 16.220 1273.210 16.280 ;
        RECT 448.660 16.080 1273.210 16.220 ;
        RECT 395.210 15.880 395.530 15.940 ;
        RECT 448.660 15.880 448.800 16.080 ;
        RECT 1272.890 16.020 1273.210 16.080 ;
        RECT 395.210 15.740 448.800 15.880 ;
        RECT 395.210 15.680 395.530 15.740 ;
      LAYER via ;
        RECT 1272.920 1688.480 1273.180 1688.740 ;
        RECT 1311.560 1688.480 1311.820 1688.740 ;
        RECT 395.240 15.680 395.500 15.940 ;
        RECT 1272.920 16.020 1273.180 16.280 ;
      LAYER met2 ;
        RECT 1311.485 1700.000 1311.765 1704.000 ;
        RECT 1311.620 1688.770 1311.760 1700.000 ;
        RECT 1272.920 1688.450 1273.180 1688.770 ;
        RECT 1311.560 1688.450 1311.820 1688.770 ;
        RECT 1272.980 16.310 1273.120 1688.450 ;
        RECT 1272.920 15.990 1273.180 16.310 ;
        RECT 395.240 15.650 395.500 15.970 ;
        RECT 395.300 2.400 395.440 15.650 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 479.390 1685.280 479.710 1685.340 ;
        RECT 1318.890 1685.280 1319.210 1685.340 ;
        RECT 479.390 1685.140 1319.210 1685.280 ;
        RECT 479.390 1685.080 479.710 1685.140 ;
        RECT 1318.890 1685.080 1319.210 1685.140 ;
        RECT 413.150 15.540 413.470 15.600 ;
        RECT 413.150 15.400 429.480 15.540 ;
        RECT 413.150 15.340 413.470 15.400 ;
        RECT 429.340 14.180 429.480 15.400 ;
        RECT 479.390 14.180 479.710 14.240 ;
        RECT 429.340 14.040 479.710 14.180 ;
        RECT 479.390 13.980 479.710 14.040 ;
      LAYER via ;
        RECT 479.420 1685.080 479.680 1685.340 ;
        RECT 1318.920 1685.080 1319.180 1685.340 ;
        RECT 413.180 15.340 413.440 15.600 ;
        RECT 479.420 13.980 479.680 14.240 ;
      LAYER met2 ;
        RECT 1318.845 1700.000 1319.125 1704.000 ;
        RECT 1318.980 1685.370 1319.120 1700.000 ;
        RECT 479.420 1685.050 479.680 1685.370 ;
        RECT 1318.920 1685.050 1319.180 1685.370 ;
        RECT 413.180 15.310 413.440 15.630 ;
        RECT 413.240 2.400 413.380 15.310 ;
        RECT 479.480 14.270 479.620 1685.050 ;
        RECT 479.420 13.950 479.680 14.270 ;
        RECT 413.030 -4.800 413.590 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1175.445 1558.985 1175.615 1593.835 ;
        RECT 1175.445 1449.165 1175.615 1497.275 ;
        RECT 1175.445 1352.605 1175.615 1400.715 ;
        RECT 1175.445 1256.045 1175.615 1304.155 ;
        RECT 1175.445 772.905 1175.615 821.015 ;
        RECT 1175.445 579.785 1175.615 627.895 ;
        RECT 1175.445 483.225 1175.615 531.335 ;
        RECT 1175.445 386.325 1175.615 434.775 ;
        RECT 1175.445 313.565 1175.615 337.875 ;
      LAYER mcon ;
        RECT 1175.445 1593.665 1175.615 1593.835 ;
        RECT 1175.445 1497.105 1175.615 1497.275 ;
        RECT 1175.445 1400.545 1175.615 1400.715 ;
        RECT 1175.445 1303.985 1175.615 1304.155 ;
        RECT 1175.445 820.845 1175.615 821.015 ;
        RECT 1175.445 627.725 1175.615 627.895 ;
        RECT 1175.445 531.165 1175.615 531.335 ;
        RECT 1175.445 434.605 1175.615 434.775 ;
        RECT 1175.445 337.705 1175.615 337.875 ;
      LAYER met1 ;
        RECT 1175.370 1593.820 1175.690 1593.880 ;
        RECT 1175.175 1593.680 1175.690 1593.820 ;
        RECT 1175.370 1593.620 1175.690 1593.680 ;
        RECT 1175.370 1559.140 1175.690 1559.200 ;
        RECT 1175.175 1559.000 1175.690 1559.140 ;
        RECT 1175.370 1558.940 1175.690 1559.000 ;
        RECT 1175.370 1497.260 1175.690 1497.320 ;
        RECT 1175.175 1497.120 1175.690 1497.260 ;
        RECT 1175.370 1497.060 1175.690 1497.120 ;
        RECT 1175.370 1449.320 1175.690 1449.380 ;
        RECT 1175.175 1449.180 1175.690 1449.320 ;
        RECT 1175.370 1449.120 1175.690 1449.180 ;
        RECT 1175.370 1400.700 1175.690 1400.760 ;
        RECT 1175.175 1400.560 1175.690 1400.700 ;
        RECT 1175.370 1400.500 1175.690 1400.560 ;
        RECT 1175.370 1352.760 1175.690 1352.820 ;
        RECT 1175.175 1352.620 1175.690 1352.760 ;
        RECT 1175.370 1352.560 1175.690 1352.620 ;
        RECT 1175.370 1304.140 1175.690 1304.200 ;
        RECT 1175.175 1304.000 1175.690 1304.140 ;
        RECT 1175.370 1303.940 1175.690 1304.000 ;
        RECT 1175.370 1256.200 1175.690 1256.260 ;
        RECT 1175.175 1256.060 1175.690 1256.200 ;
        RECT 1175.370 1256.000 1175.690 1256.060 ;
        RECT 1174.450 1159.300 1174.770 1159.360 ;
        RECT 1175.370 1159.300 1175.690 1159.360 ;
        RECT 1174.450 1159.160 1175.690 1159.300 ;
        RECT 1174.450 1159.100 1174.770 1159.160 ;
        RECT 1175.370 1159.100 1175.690 1159.160 ;
        RECT 1174.450 1062.740 1174.770 1062.800 ;
        RECT 1175.370 1062.740 1175.690 1062.800 ;
        RECT 1174.450 1062.600 1175.690 1062.740 ;
        RECT 1174.450 1062.540 1174.770 1062.600 ;
        RECT 1175.370 1062.540 1175.690 1062.600 ;
        RECT 1175.370 979.580 1175.690 979.840 ;
        RECT 1175.460 979.160 1175.600 979.580 ;
        RECT 1175.370 978.900 1175.690 979.160 ;
        RECT 1175.370 883.020 1175.690 883.280 ;
        RECT 1175.460 882.600 1175.600 883.020 ;
        RECT 1175.370 882.340 1175.690 882.600 ;
        RECT 1175.370 821.000 1175.690 821.060 ;
        RECT 1175.175 820.860 1175.690 821.000 ;
        RECT 1175.370 820.800 1175.690 820.860 ;
        RECT 1175.370 773.060 1175.690 773.120 ;
        RECT 1175.175 772.920 1175.690 773.060 ;
        RECT 1175.370 772.860 1175.690 772.920 ;
        RECT 1175.370 738.520 1175.690 738.780 ;
        RECT 1175.460 738.100 1175.600 738.520 ;
        RECT 1175.370 737.840 1175.690 738.100 ;
        RECT 1175.370 689.900 1175.690 690.160 ;
        RECT 1175.460 689.480 1175.600 689.900 ;
        RECT 1175.370 689.220 1175.690 689.480 ;
        RECT 1175.370 627.880 1175.690 627.940 ;
        RECT 1175.175 627.740 1175.690 627.880 ;
        RECT 1175.370 627.680 1175.690 627.740 ;
        RECT 1175.370 579.940 1175.690 580.000 ;
        RECT 1175.175 579.800 1175.690 579.940 ;
        RECT 1175.370 579.740 1175.690 579.800 ;
        RECT 1175.370 531.320 1175.690 531.380 ;
        RECT 1175.175 531.180 1175.690 531.320 ;
        RECT 1175.370 531.120 1175.690 531.180 ;
        RECT 1175.370 483.380 1175.690 483.440 ;
        RECT 1175.175 483.240 1175.690 483.380 ;
        RECT 1175.370 483.180 1175.690 483.240 ;
        RECT 1175.370 434.760 1175.690 434.820 ;
        RECT 1175.175 434.620 1175.690 434.760 ;
        RECT 1175.370 434.560 1175.690 434.620 ;
        RECT 1175.370 386.480 1175.690 386.540 ;
        RECT 1175.175 386.340 1175.690 386.480 ;
        RECT 1175.370 386.280 1175.690 386.340 ;
        RECT 1175.370 337.860 1175.690 337.920 ;
        RECT 1175.175 337.720 1175.690 337.860 ;
        RECT 1175.370 337.660 1175.690 337.720 ;
        RECT 1175.370 313.720 1175.690 313.780 ;
        RECT 1175.175 313.580 1175.690 313.720 ;
        RECT 1175.370 313.520 1175.690 313.580 ;
        RECT 74.130 17.580 74.450 17.640 ;
        RECT 1174.450 17.580 1174.770 17.640 ;
        RECT 74.130 17.440 1174.770 17.580 ;
        RECT 74.130 17.380 74.450 17.440 ;
        RECT 1174.450 17.380 1174.770 17.440 ;
      LAYER via ;
        RECT 1175.400 1593.620 1175.660 1593.880 ;
        RECT 1175.400 1558.940 1175.660 1559.200 ;
        RECT 1175.400 1497.060 1175.660 1497.320 ;
        RECT 1175.400 1449.120 1175.660 1449.380 ;
        RECT 1175.400 1400.500 1175.660 1400.760 ;
        RECT 1175.400 1352.560 1175.660 1352.820 ;
        RECT 1175.400 1303.940 1175.660 1304.200 ;
        RECT 1175.400 1256.000 1175.660 1256.260 ;
        RECT 1174.480 1159.100 1174.740 1159.360 ;
        RECT 1175.400 1159.100 1175.660 1159.360 ;
        RECT 1174.480 1062.540 1174.740 1062.800 ;
        RECT 1175.400 1062.540 1175.660 1062.800 ;
        RECT 1175.400 979.580 1175.660 979.840 ;
        RECT 1175.400 978.900 1175.660 979.160 ;
        RECT 1175.400 883.020 1175.660 883.280 ;
        RECT 1175.400 882.340 1175.660 882.600 ;
        RECT 1175.400 820.800 1175.660 821.060 ;
        RECT 1175.400 772.860 1175.660 773.120 ;
        RECT 1175.400 738.520 1175.660 738.780 ;
        RECT 1175.400 737.840 1175.660 738.100 ;
        RECT 1175.400 689.900 1175.660 690.160 ;
        RECT 1175.400 689.220 1175.660 689.480 ;
        RECT 1175.400 627.680 1175.660 627.940 ;
        RECT 1175.400 579.740 1175.660 580.000 ;
        RECT 1175.400 531.120 1175.660 531.380 ;
        RECT 1175.400 483.180 1175.660 483.440 ;
        RECT 1175.400 434.560 1175.660 434.820 ;
        RECT 1175.400 386.280 1175.660 386.540 ;
        RECT 1175.400 337.660 1175.660 337.920 ;
        RECT 1175.400 313.520 1175.660 313.780 ;
        RECT 74.160 17.380 74.420 17.640 ;
        RECT 1174.480 17.380 1174.740 17.640 ;
      LAYER met2 ;
        RECT 1179.005 1700.410 1179.285 1704.000 ;
        RECT 1177.300 1700.270 1179.285 1700.410 ;
        RECT 1177.300 1677.970 1177.440 1700.270 ;
        RECT 1179.005 1700.000 1179.285 1700.270 ;
        RECT 1175.460 1677.830 1177.440 1677.970 ;
        RECT 1175.460 1593.910 1175.600 1677.830 ;
        RECT 1175.400 1593.590 1175.660 1593.910 ;
        RECT 1175.400 1558.910 1175.660 1559.230 ;
        RECT 1175.460 1497.350 1175.600 1558.910 ;
        RECT 1175.400 1497.030 1175.660 1497.350 ;
        RECT 1175.400 1449.090 1175.660 1449.410 ;
        RECT 1175.460 1400.790 1175.600 1449.090 ;
        RECT 1175.400 1400.470 1175.660 1400.790 ;
        RECT 1175.400 1352.530 1175.660 1352.850 ;
        RECT 1175.460 1304.230 1175.600 1352.530 ;
        RECT 1175.400 1303.910 1175.660 1304.230 ;
        RECT 1175.400 1255.970 1175.660 1256.290 ;
        RECT 1175.460 1207.525 1175.600 1255.970 ;
        RECT 1174.470 1207.155 1174.750 1207.525 ;
        RECT 1175.390 1207.155 1175.670 1207.525 ;
        RECT 1174.540 1159.390 1174.680 1207.155 ;
        RECT 1174.480 1159.070 1174.740 1159.390 ;
        RECT 1175.400 1159.070 1175.660 1159.390 ;
        RECT 1175.460 1110.965 1175.600 1159.070 ;
        RECT 1174.470 1110.595 1174.750 1110.965 ;
        RECT 1175.390 1110.595 1175.670 1110.965 ;
        RECT 1174.540 1062.830 1174.680 1110.595 ;
        RECT 1174.480 1062.510 1174.740 1062.830 ;
        RECT 1175.400 1062.510 1175.660 1062.830 ;
        RECT 1175.460 979.870 1175.600 1062.510 ;
        RECT 1175.400 979.550 1175.660 979.870 ;
        RECT 1175.400 978.870 1175.660 979.190 ;
        RECT 1175.460 883.310 1175.600 978.870 ;
        RECT 1175.400 882.990 1175.660 883.310 ;
        RECT 1175.400 882.310 1175.660 882.630 ;
        RECT 1175.460 821.090 1175.600 882.310 ;
        RECT 1175.400 820.770 1175.660 821.090 ;
        RECT 1175.400 772.830 1175.660 773.150 ;
        RECT 1175.460 738.810 1175.600 772.830 ;
        RECT 1175.400 738.490 1175.660 738.810 ;
        RECT 1175.400 737.810 1175.660 738.130 ;
        RECT 1175.460 690.190 1175.600 737.810 ;
        RECT 1175.400 689.870 1175.660 690.190 ;
        RECT 1175.400 689.190 1175.660 689.510 ;
        RECT 1175.460 627.970 1175.600 689.190 ;
        RECT 1175.400 627.650 1175.660 627.970 ;
        RECT 1175.400 579.710 1175.660 580.030 ;
        RECT 1175.460 531.410 1175.600 579.710 ;
        RECT 1175.400 531.090 1175.660 531.410 ;
        RECT 1175.400 483.150 1175.660 483.470 ;
        RECT 1175.460 434.850 1175.600 483.150 ;
        RECT 1175.400 434.530 1175.660 434.850 ;
        RECT 1175.400 386.250 1175.660 386.570 ;
        RECT 1175.460 337.950 1175.600 386.250 ;
        RECT 1175.400 337.630 1175.660 337.950 ;
        RECT 1175.400 313.490 1175.660 313.810 ;
        RECT 1175.460 207.130 1175.600 313.490 ;
        RECT 1175.000 206.990 1175.600 207.130 ;
        RECT 1175.000 206.450 1175.140 206.990 ;
        RECT 1175.000 206.310 1175.600 206.450 ;
        RECT 1175.460 110.570 1175.600 206.310 ;
        RECT 1175.000 110.430 1175.600 110.570 ;
        RECT 1175.000 61.610 1175.140 110.430 ;
        RECT 1174.540 61.470 1175.140 61.610 ;
        RECT 1174.540 17.670 1174.680 61.470 ;
        RECT 74.160 17.350 74.420 17.670 ;
        RECT 1174.480 17.350 1174.740 17.670 ;
        RECT 74.220 2.400 74.360 17.350 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 1174.470 1207.200 1174.750 1207.480 ;
        RECT 1175.390 1207.200 1175.670 1207.480 ;
        RECT 1174.470 1110.640 1174.750 1110.920 ;
        RECT 1175.390 1110.640 1175.670 1110.920 ;
      LAYER met3 ;
        RECT 1174.445 1207.490 1174.775 1207.505 ;
        RECT 1175.365 1207.490 1175.695 1207.505 ;
        RECT 1174.445 1207.190 1175.695 1207.490 ;
        RECT 1174.445 1207.175 1174.775 1207.190 ;
        RECT 1175.365 1207.175 1175.695 1207.190 ;
        RECT 1174.445 1110.930 1174.775 1110.945 ;
        RECT 1175.365 1110.930 1175.695 1110.945 ;
        RECT 1174.445 1110.630 1175.695 1110.930 ;
        RECT 1174.445 1110.615 1174.775 1110.630 ;
        RECT 1175.365 1110.615 1175.695 1110.630 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 513.890 1684.600 514.210 1684.660 ;
        RECT 1326.250 1684.600 1326.570 1684.660 ;
        RECT 513.890 1684.460 1326.570 1684.600 ;
        RECT 513.890 1684.400 514.210 1684.460 ;
        RECT 1326.250 1684.400 1326.570 1684.460 ;
        RECT 430.630 15.200 430.950 15.260 ;
        RECT 430.630 15.060 475.940 15.200 ;
        RECT 430.630 15.000 430.950 15.060 ;
        RECT 475.800 14.860 475.940 15.060 ;
        RECT 475.800 14.720 482.840 14.860 ;
        RECT 482.700 14.180 482.840 14.720 ;
        RECT 512.970 14.180 513.290 14.240 ;
        RECT 482.700 14.040 513.290 14.180 ;
        RECT 512.970 13.980 513.290 14.040 ;
      LAYER via ;
        RECT 513.920 1684.400 514.180 1684.660 ;
        RECT 1326.280 1684.400 1326.540 1684.660 ;
        RECT 430.660 15.000 430.920 15.260 ;
        RECT 513.000 13.980 513.260 14.240 ;
      LAYER met2 ;
        RECT 1326.205 1700.000 1326.485 1704.000 ;
        RECT 1326.340 1684.690 1326.480 1700.000 ;
        RECT 513.920 1684.370 514.180 1684.690 ;
        RECT 1326.280 1684.370 1326.540 1684.690 ;
        RECT 513.980 16.050 514.120 1684.370 ;
        RECT 513.060 15.910 514.120 16.050 ;
        RECT 430.660 14.970 430.920 15.290 ;
        RECT 430.720 2.400 430.860 14.970 ;
        RECT 513.060 14.270 513.200 15.910 ;
        RECT 513.000 13.950 513.260 14.270 ;
        RECT 430.510 -4.800 431.070 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1333.610 1686.980 1333.930 1687.040 ;
        RECT 1304.720 1686.840 1333.930 1686.980 ;
        RECT 1279.790 1686.300 1280.110 1686.360 ;
        RECT 1304.720 1686.300 1304.860 1686.840 ;
        RECT 1333.610 1686.780 1333.930 1686.840 ;
        RECT 1279.790 1686.160 1304.860 1686.300 ;
        RECT 1279.790 1686.100 1280.110 1686.160 ;
        RECT 1279.790 15.880 1280.110 15.940 ;
        RECT 472.120 15.740 1280.110 15.880 ;
        RECT 448.570 15.540 448.890 15.600 ;
        RECT 472.120 15.540 472.260 15.740 ;
        RECT 1279.790 15.680 1280.110 15.740 ;
        RECT 448.570 15.400 472.260 15.540 ;
        RECT 448.570 15.340 448.890 15.400 ;
      LAYER via ;
        RECT 1279.820 1686.100 1280.080 1686.360 ;
        RECT 1333.640 1686.780 1333.900 1687.040 ;
        RECT 448.600 15.340 448.860 15.600 ;
        RECT 1279.820 15.680 1280.080 15.940 ;
      LAYER met2 ;
        RECT 1333.565 1700.000 1333.845 1704.000 ;
        RECT 1333.700 1687.070 1333.840 1700.000 ;
        RECT 1333.640 1686.750 1333.900 1687.070 ;
        RECT 1279.820 1686.070 1280.080 1686.390 ;
        RECT 1279.880 15.970 1280.020 1686.070 ;
        RECT 1279.820 15.650 1280.080 15.970 ;
        RECT 448.600 15.310 448.860 15.630 ;
        RECT 448.660 2.400 448.800 15.310 ;
        RECT 448.450 -4.800 449.010 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 474.865 15.045 476.415 15.215 ;
        RECT 474.865 14.705 475.035 15.045 ;
      LAYER mcon ;
        RECT 476.245 15.045 476.415 15.215 ;
      LAYER met1 ;
        RECT 486.290 1685.960 486.610 1686.020 ;
        RECT 1340.970 1685.960 1341.290 1686.020 ;
        RECT 486.290 1685.820 1341.290 1685.960 ;
        RECT 486.290 1685.760 486.610 1685.820 ;
        RECT 1340.970 1685.760 1341.290 1685.820 ;
        RECT 476.185 15.200 476.475 15.245 ;
        RECT 486.290 15.200 486.610 15.260 ;
        RECT 476.185 15.060 486.610 15.200 ;
        RECT 476.185 15.015 476.475 15.060 ;
        RECT 486.290 15.000 486.610 15.060 ;
        RECT 466.510 14.860 466.830 14.920 ;
        RECT 474.805 14.860 475.095 14.905 ;
        RECT 466.510 14.720 475.095 14.860 ;
        RECT 466.510 14.660 466.830 14.720 ;
        RECT 474.805 14.675 475.095 14.720 ;
      LAYER via ;
        RECT 486.320 1685.760 486.580 1686.020 ;
        RECT 1341.000 1685.760 1341.260 1686.020 ;
        RECT 486.320 15.000 486.580 15.260 ;
        RECT 466.540 14.660 466.800 14.920 ;
      LAYER met2 ;
        RECT 1340.925 1700.000 1341.205 1704.000 ;
        RECT 1341.060 1686.050 1341.200 1700.000 ;
        RECT 486.320 1685.730 486.580 1686.050 ;
        RECT 1341.000 1685.730 1341.260 1686.050 ;
        RECT 486.380 15.290 486.520 1685.730 ;
        RECT 486.320 14.970 486.580 15.290 ;
        RECT 466.540 14.630 466.800 14.950 ;
        RECT 466.600 2.400 466.740 14.630 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1348.330 1687.320 1348.650 1687.380 ;
        RECT 1301.960 1687.180 1348.650 1687.320 ;
        RECT 1286.690 1686.980 1287.010 1687.040 ;
        RECT 1301.960 1686.980 1302.100 1687.180 ;
        RECT 1348.330 1687.120 1348.650 1687.180 ;
        RECT 1286.690 1686.840 1302.100 1686.980 ;
        RECT 1286.690 1686.780 1287.010 1686.840 ;
        RECT 1286.690 15.540 1287.010 15.600 ;
        RECT 541.580 15.400 1287.010 15.540 ;
        RECT 484.450 14.860 484.770 14.920 ;
        RECT 541.580 14.860 541.720 15.400 ;
        RECT 1286.690 15.340 1287.010 15.400 ;
        RECT 484.450 14.720 541.720 14.860 ;
        RECT 484.450 14.660 484.770 14.720 ;
      LAYER via ;
        RECT 1286.720 1686.780 1286.980 1687.040 ;
        RECT 1348.360 1687.120 1348.620 1687.380 ;
        RECT 484.480 14.660 484.740 14.920 ;
        RECT 1286.720 15.340 1286.980 15.600 ;
      LAYER met2 ;
        RECT 1348.285 1700.000 1348.565 1704.000 ;
        RECT 1348.420 1687.410 1348.560 1700.000 ;
        RECT 1348.360 1687.090 1348.620 1687.410 ;
        RECT 1286.720 1686.750 1286.980 1687.070 ;
        RECT 1286.780 15.630 1286.920 1686.750 ;
        RECT 1286.720 15.310 1286.980 15.630 ;
        RECT 484.480 14.630 484.740 14.950 ;
        RECT 484.540 2.400 484.680 14.630 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 503.310 1685.620 503.630 1685.680 ;
        RECT 1355.690 1685.620 1356.010 1685.680 ;
        RECT 503.310 1685.480 1356.010 1685.620 ;
        RECT 503.310 1685.420 503.630 1685.480 ;
        RECT 1355.690 1685.420 1356.010 1685.480 ;
      LAYER via ;
        RECT 503.340 1685.420 503.600 1685.680 ;
        RECT 1355.720 1685.420 1355.980 1685.680 ;
      LAYER met2 ;
        RECT 1355.645 1700.000 1355.925 1704.000 ;
        RECT 1355.780 1685.710 1355.920 1700.000 ;
        RECT 503.340 1685.390 503.600 1685.710 ;
        RECT 1355.720 1685.390 1355.980 1685.710 ;
        RECT 503.400 16.730 503.540 1685.390 ;
        RECT 502.480 16.590 503.540 16.730 ;
        RECT 502.480 2.400 502.620 16.590 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1294.050 1689.360 1294.370 1689.420 ;
        RECT 1363.050 1689.360 1363.370 1689.420 ;
        RECT 1294.050 1689.220 1363.370 1689.360 ;
        RECT 1294.050 1689.160 1294.370 1689.220 ;
        RECT 1363.050 1689.160 1363.370 1689.220 ;
        RECT 1294.050 15.200 1294.370 15.260 ;
        RECT 542.040 15.060 1294.370 15.200 ;
        RECT 519.870 14.520 520.190 14.580 ;
        RECT 542.040 14.520 542.180 15.060 ;
        RECT 1294.050 15.000 1294.370 15.060 ;
        RECT 519.870 14.380 542.180 14.520 ;
        RECT 519.870 14.320 520.190 14.380 ;
      LAYER via ;
        RECT 1294.080 1689.160 1294.340 1689.420 ;
        RECT 1363.080 1689.160 1363.340 1689.420 ;
        RECT 519.900 14.320 520.160 14.580 ;
        RECT 1294.080 15.000 1294.340 15.260 ;
      LAYER met2 ;
        RECT 1363.005 1700.000 1363.285 1704.000 ;
        RECT 1363.140 1689.450 1363.280 1700.000 ;
        RECT 1294.080 1689.130 1294.340 1689.450 ;
        RECT 1363.080 1689.130 1363.340 1689.450 ;
        RECT 1294.140 15.290 1294.280 1689.130 ;
        RECT 1294.080 14.970 1294.340 15.290 ;
        RECT 519.900 14.290 520.160 14.610 ;
        RECT 519.960 2.400 520.100 14.290 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 537.810 1684.940 538.130 1685.000 ;
        RECT 1370.410 1684.940 1370.730 1685.000 ;
        RECT 537.810 1684.800 1370.730 1684.940 ;
        RECT 537.810 1684.740 538.130 1684.800 ;
        RECT 1370.410 1684.740 1370.730 1684.800 ;
      LAYER via ;
        RECT 537.840 1684.740 538.100 1685.000 ;
        RECT 1370.440 1684.740 1370.700 1685.000 ;
      LAYER met2 ;
        RECT 1370.365 1700.000 1370.645 1704.000 ;
        RECT 1370.500 1685.030 1370.640 1700.000 ;
        RECT 537.840 1684.710 538.100 1685.030 ;
        RECT 1370.440 1684.710 1370.700 1685.030 ;
        RECT 537.900 2.400 538.040 1684.710 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1377.770 1687.660 1378.090 1687.720 ;
        RECT 1301.500 1687.520 1378.090 1687.660 ;
        RECT 1293.590 1687.320 1293.910 1687.380 ;
        RECT 1301.500 1687.320 1301.640 1687.520 ;
        RECT 1377.770 1687.460 1378.090 1687.520 ;
        RECT 1293.590 1687.180 1301.640 1687.320 ;
        RECT 1293.590 1687.120 1293.910 1687.180 ;
        RECT 1293.590 14.860 1293.910 14.920 ;
        RECT 607.360 14.720 1293.910 14.860 ;
        RECT 555.750 14.520 556.070 14.580 ;
        RECT 607.360 14.520 607.500 14.720 ;
        RECT 1293.590 14.660 1293.910 14.720 ;
        RECT 555.750 14.380 607.500 14.520 ;
        RECT 555.750 14.320 556.070 14.380 ;
      LAYER via ;
        RECT 1293.620 1687.120 1293.880 1687.380 ;
        RECT 1377.800 1687.460 1378.060 1687.720 ;
        RECT 555.780 14.320 556.040 14.580 ;
        RECT 1293.620 14.660 1293.880 14.920 ;
      LAYER met2 ;
        RECT 1377.725 1700.000 1378.005 1704.000 ;
        RECT 1377.860 1687.750 1378.000 1700.000 ;
        RECT 1377.800 1687.430 1378.060 1687.750 ;
        RECT 1293.620 1687.090 1293.880 1687.410 ;
        RECT 1293.680 14.950 1293.820 1687.090 ;
        RECT 1293.620 14.630 1293.880 14.950 ;
        RECT 555.780 14.290 556.040 14.610 ;
        RECT 555.840 2.400 555.980 14.290 ;
        RECT 555.630 -4.800 556.190 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1300.490 1688.340 1300.810 1688.400 ;
        RECT 1385.130 1688.340 1385.450 1688.400 ;
        RECT 1300.490 1688.200 1385.450 1688.340 ;
        RECT 1300.490 1688.140 1300.810 1688.200 ;
        RECT 1385.130 1688.140 1385.450 1688.200 ;
        RECT 1300.490 14.520 1300.810 14.580 ;
        RECT 607.820 14.380 1300.810 14.520 ;
        RECT 573.690 14.180 574.010 14.240 ;
        RECT 607.820 14.180 607.960 14.380 ;
        RECT 1300.490 14.320 1300.810 14.380 ;
        RECT 573.690 14.040 607.960 14.180 ;
        RECT 573.690 13.980 574.010 14.040 ;
      LAYER via ;
        RECT 1300.520 1688.140 1300.780 1688.400 ;
        RECT 1385.160 1688.140 1385.420 1688.400 ;
        RECT 573.720 13.980 573.980 14.240 ;
        RECT 1300.520 14.320 1300.780 14.580 ;
      LAYER met2 ;
        RECT 1385.085 1700.000 1385.365 1704.000 ;
        RECT 1385.220 1688.430 1385.360 1700.000 ;
        RECT 1300.520 1688.110 1300.780 1688.430 ;
        RECT 1385.160 1688.110 1385.420 1688.430 ;
        RECT 1300.580 14.610 1300.720 1688.110 ;
        RECT 1300.520 14.290 1300.780 14.610 ;
        RECT 573.720 13.950 573.980 14.270 ;
        RECT 573.780 2.400 573.920 13.950 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 593.010 1684.260 593.330 1684.320 ;
        RECT 1392.490 1684.260 1392.810 1684.320 ;
        RECT 593.010 1684.120 1392.810 1684.260 ;
        RECT 593.010 1684.060 593.330 1684.120 ;
        RECT 1392.490 1684.060 1392.810 1684.120 ;
      LAYER via ;
        RECT 593.040 1684.060 593.300 1684.320 ;
        RECT 1392.520 1684.060 1392.780 1684.320 ;
      LAYER met2 ;
        RECT 1392.445 1700.000 1392.725 1704.000 ;
        RECT 1392.580 1684.350 1392.720 1700.000 ;
        RECT 593.040 1684.030 593.300 1684.350 ;
        RECT 1392.520 1684.030 1392.780 1684.350 ;
        RECT 593.100 16.730 593.240 1684.030 ;
        RECT 591.260 16.590 593.240 16.730 ;
        RECT 591.260 2.400 591.400 16.590 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 141.290 1687.660 141.610 1687.720 ;
        RECT 141.290 1687.520 1172.380 1687.660 ;
        RECT 141.290 1687.460 141.610 1687.520 ;
        RECT 1172.240 1687.320 1172.380 1687.520 ;
        RECT 1189.170 1687.320 1189.490 1687.380 ;
        RECT 1172.240 1687.180 1189.490 1687.320 ;
        RECT 1189.170 1687.120 1189.490 1687.180 ;
        RECT 97.590 16.900 97.910 16.960 ;
        RECT 141.290 16.900 141.610 16.960 ;
        RECT 97.590 16.760 141.610 16.900 ;
        RECT 97.590 16.700 97.910 16.760 ;
        RECT 141.290 16.700 141.610 16.760 ;
      LAYER via ;
        RECT 141.320 1687.460 141.580 1687.720 ;
        RECT 1189.200 1687.120 1189.460 1687.380 ;
        RECT 97.620 16.700 97.880 16.960 ;
        RECT 141.320 16.700 141.580 16.960 ;
      LAYER met2 ;
        RECT 1189.125 1700.000 1189.405 1704.000 ;
        RECT 141.320 1687.430 141.580 1687.750 ;
        RECT 141.380 16.990 141.520 1687.430 ;
        RECT 1189.260 1687.410 1189.400 1700.000 ;
        RECT 1189.200 1687.090 1189.460 1687.410 ;
        RECT 97.620 16.670 97.880 16.990 ;
        RECT 141.320 16.670 141.580 16.990 ;
        RECT 97.680 2.400 97.820 16.670 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1306.930 1688.000 1307.250 1688.060 ;
        RECT 1399.850 1688.000 1400.170 1688.060 ;
        RECT 1306.930 1687.860 1400.170 1688.000 ;
        RECT 1306.930 1687.800 1307.250 1687.860 ;
        RECT 1399.850 1687.800 1400.170 1687.860 ;
        RECT 609.110 14.180 609.430 14.240 ;
        RECT 1307.390 14.180 1307.710 14.240 ;
        RECT 609.110 14.040 1307.710 14.180 ;
        RECT 609.110 13.980 609.430 14.040 ;
        RECT 1307.390 13.980 1307.710 14.040 ;
      LAYER via ;
        RECT 1306.960 1687.800 1307.220 1688.060 ;
        RECT 1399.880 1687.800 1400.140 1688.060 ;
        RECT 609.140 13.980 609.400 14.240 ;
        RECT 1307.420 13.980 1307.680 14.240 ;
      LAYER met2 ;
        RECT 1399.805 1700.000 1400.085 1704.000 ;
        RECT 1399.940 1688.090 1400.080 1700.000 ;
        RECT 1306.960 1687.770 1307.220 1688.090 ;
        RECT 1399.880 1687.770 1400.140 1688.090 ;
        RECT 1307.020 1671.850 1307.160 1687.770 ;
        RECT 1307.020 1671.710 1307.620 1671.850 ;
        RECT 1307.480 14.270 1307.620 1671.710 ;
        RECT 609.140 13.950 609.400 14.270 ;
        RECT 1307.420 13.950 1307.680 14.270 ;
        RECT 609.200 2.400 609.340 13.950 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 627.510 1683.920 627.830 1683.980 ;
        RECT 1405.830 1683.920 1406.150 1683.980 ;
        RECT 627.510 1683.780 1406.150 1683.920 ;
        RECT 627.510 1683.720 627.830 1683.780 ;
        RECT 1405.830 1683.720 1406.150 1683.780 ;
      LAYER via ;
        RECT 627.540 1683.720 627.800 1683.980 ;
        RECT 1405.860 1683.720 1406.120 1683.980 ;
      LAYER met2 ;
        RECT 1407.165 1700.410 1407.445 1704.000 ;
        RECT 1405.920 1700.270 1407.445 1700.410 ;
        RECT 1405.920 1684.010 1406.060 1700.270 ;
        RECT 1407.165 1700.000 1407.445 1700.270 ;
        RECT 627.540 1683.690 627.800 1684.010 ;
        RECT 1405.860 1683.690 1406.120 1684.010 ;
        RECT 627.600 17.410 627.740 1683.690 ;
        RECT 627.140 17.270 627.740 17.410 ;
        RECT 627.140 2.400 627.280 17.270 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1195.610 1558.260 1195.930 1558.520 ;
        RECT 1195.700 1557.840 1195.840 1558.260 ;
        RECT 1195.610 1557.580 1195.930 1557.840 ;
        RECT 1195.610 1462.380 1195.930 1462.640 ;
        RECT 1195.700 1461.960 1195.840 1462.380 ;
        RECT 1195.610 1461.700 1195.930 1461.960 ;
        RECT 1195.610 1365.820 1195.930 1366.080 ;
        RECT 1195.700 1365.400 1195.840 1365.820 ;
        RECT 1195.610 1365.140 1195.930 1365.400 ;
        RECT 1195.610 1269.260 1195.930 1269.520 ;
        RECT 1195.700 1268.840 1195.840 1269.260 ;
        RECT 1195.610 1268.580 1195.930 1268.840 ;
        RECT 1195.610 1172.700 1195.930 1172.960 ;
        RECT 1195.700 1172.280 1195.840 1172.700 ;
        RECT 1195.610 1172.020 1195.930 1172.280 ;
        RECT 1195.610 1076.140 1195.930 1076.400 ;
        RECT 1195.700 1075.720 1195.840 1076.140 ;
        RECT 1195.610 1075.460 1195.930 1075.720 ;
        RECT 1195.610 882.340 1195.930 882.600 ;
        RECT 1195.700 881.920 1195.840 882.340 ;
        RECT 1195.610 881.660 1195.930 881.920 ;
        RECT 121.510 18.260 121.830 18.320 ;
        RECT 1195.150 18.260 1195.470 18.320 ;
        RECT 121.510 18.120 1195.470 18.260 ;
        RECT 121.510 18.060 121.830 18.120 ;
        RECT 1195.150 18.060 1195.470 18.120 ;
      LAYER via ;
        RECT 1195.640 1558.260 1195.900 1558.520 ;
        RECT 1195.640 1557.580 1195.900 1557.840 ;
        RECT 1195.640 1462.380 1195.900 1462.640 ;
        RECT 1195.640 1461.700 1195.900 1461.960 ;
        RECT 1195.640 1365.820 1195.900 1366.080 ;
        RECT 1195.640 1365.140 1195.900 1365.400 ;
        RECT 1195.640 1269.260 1195.900 1269.520 ;
        RECT 1195.640 1268.580 1195.900 1268.840 ;
        RECT 1195.640 1172.700 1195.900 1172.960 ;
        RECT 1195.640 1172.020 1195.900 1172.280 ;
        RECT 1195.640 1076.140 1195.900 1076.400 ;
        RECT 1195.640 1075.460 1195.900 1075.720 ;
        RECT 1195.640 882.340 1195.900 882.600 ;
        RECT 1195.640 881.660 1195.900 881.920 ;
        RECT 121.540 18.060 121.800 18.320 ;
        RECT 1195.180 18.060 1195.440 18.320 ;
      LAYER met2 ;
        RECT 1198.785 1700.410 1199.065 1704.000 ;
        RECT 1197.540 1700.270 1199.065 1700.410 ;
        RECT 1197.540 1656.210 1197.680 1700.270 ;
        RECT 1198.785 1700.000 1199.065 1700.270 ;
        RECT 1195.700 1656.070 1197.680 1656.210 ;
        RECT 1195.700 1558.550 1195.840 1656.070 ;
        RECT 1195.640 1558.230 1195.900 1558.550 ;
        RECT 1195.640 1557.550 1195.900 1557.870 ;
        RECT 1195.700 1462.670 1195.840 1557.550 ;
        RECT 1195.640 1462.350 1195.900 1462.670 ;
        RECT 1195.640 1461.670 1195.900 1461.990 ;
        RECT 1195.700 1366.110 1195.840 1461.670 ;
        RECT 1195.640 1365.790 1195.900 1366.110 ;
        RECT 1195.640 1365.110 1195.900 1365.430 ;
        RECT 1195.700 1269.550 1195.840 1365.110 ;
        RECT 1195.640 1269.230 1195.900 1269.550 ;
        RECT 1195.640 1268.550 1195.900 1268.870 ;
        RECT 1195.700 1172.990 1195.840 1268.550 ;
        RECT 1195.640 1172.670 1195.900 1172.990 ;
        RECT 1195.640 1171.990 1195.900 1172.310 ;
        RECT 1195.700 1076.430 1195.840 1171.990 ;
        RECT 1195.640 1076.110 1195.900 1076.430 ;
        RECT 1195.640 1075.430 1195.900 1075.750 ;
        RECT 1195.700 882.630 1195.840 1075.430 ;
        RECT 1195.640 882.310 1195.900 882.630 ;
        RECT 1195.640 881.630 1195.900 881.950 ;
        RECT 1195.700 642.330 1195.840 881.630 ;
        RECT 1195.240 642.190 1195.840 642.330 ;
        RECT 1195.240 641.650 1195.380 642.190 ;
        RECT 1195.240 641.510 1195.840 641.650 ;
        RECT 1195.700 497.490 1195.840 641.510 ;
        RECT 1195.240 497.350 1195.840 497.490 ;
        RECT 1195.240 496.810 1195.380 497.350 ;
        RECT 1195.240 496.670 1195.840 496.810 ;
        RECT 1195.700 303.690 1195.840 496.670 ;
        RECT 1195.240 303.550 1195.840 303.690 ;
        RECT 1195.240 303.010 1195.380 303.550 ;
        RECT 1195.240 302.870 1195.840 303.010 ;
        RECT 1195.700 207.130 1195.840 302.870 ;
        RECT 1195.240 206.990 1195.840 207.130 ;
        RECT 1195.240 206.450 1195.380 206.990 ;
        RECT 1195.240 206.310 1195.840 206.450 ;
        RECT 1195.700 62.290 1195.840 206.310 ;
        RECT 1195.700 62.150 1196.300 62.290 ;
        RECT 1196.160 61.610 1196.300 62.150 ;
        RECT 1195.240 61.470 1196.300 61.610 ;
        RECT 1195.240 18.350 1195.380 61.470 ;
        RECT 121.540 18.030 121.800 18.350 ;
        RECT 1195.180 18.030 1195.440 18.350 ;
        RECT 121.600 2.400 121.740 18.030 ;
        RECT 121.390 -4.800 121.950 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 161.990 1688.000 162.310 1688.060 ;
        RECT 1208.490 1688.000 1208.810 1688.060 ;
        RECT 161.990 1687.860 1208.810 1688.000 ;
        RECT 161.990 1687.800 162.310 1687.860 ;
        RECT 1208.490 1687.800 1208.810 1687.860 ;
        RECT 145.430 16.900 145.750 16.960 ;
        RECT 161.990 16.900 162.310 16.960 ;
        RECT 145.430 16.760 162.310 16.900 ;
        RECT 145.430 16.700 145.750 16.760 ;
        RECT 161.990 16.700 162.310 16.760 ;
      LAYER via ;
        RECT 162.020 1687.800 162.280 1688.060 ;
        RECT 1208.520 1687.800 1208.780 1688.060 ;
        RECT 145.460 16.700 145.720 16.960 ;
        RECT 162.020 16.700 162.280 16.960 ;
      LAYER met2 ;
        RECT 1208.445 1700.000 1208.725 1704.000 ;
        RECT 1208.580 1688.090 1208.720 1700.000 ;
        RECT 162.020 1687.770 162.280 1688.090 ;
        RECT 1208.520 1687.770 1208.780 1688.090 ;
        RECT 162.080 16.990 162.220 1687.770 ;
        RECT 145.460 16.670 145.720 16.990 ;
        RECT 162.020 16.670 162.280 16.990 ;
        RECT 145.520 2.400 145.660 16.670 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 163.370 18.600 163.690 18.660 ;
        RECT 1215.390 18.600 1215.710 18.660 ;
        RECT 163.370 18.460 1215.710 18.600 ;
        RECT 163.370 18.400 163.690 18.460 ;
        RECT 1215.390 18.400 1215.710 18.460 ;
      LAYER via ;
        RECT 163.400 18.400 163.660 18.660 ;
        RECT 1215.420 18.400 1215.680 18.660 ;
      LAYER met2 ;
        RECT 1215.805 1700.410 1216.085 1704.000 ;
        RECT 1215.480 1700.270 1216.085 1700.410 ;
        RECT 1215.480 18.690 1215.620 1700.270 ;
        RECT 1215.805 1700.000 1216.085 1700.270 ;
        RECT 163.400 18.370 163.660 18.690 ;
        RECT 1215.420 18.370 1215.680 18.690 ;
        RECT 163.460 2.400 163.600 18.370 ;
        RECT 163.250 -4.800 163.810 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 196.490 1688.340 196.810 1688.400 ;
        RECT 1223.210 1688.340 1223.530 1688.400 ;
        RECT 196.490 1688.200 1223.530 1688.340 ;
        RECT 196.490 1688.140 196.810 1688.200 ;
        RECT 1223.210 1688.140 1223.530 1688.200 ;
        RECT 180.850 15.200 181.170 15.260 ;
        RECT 196.490 15.200 196.810 15.260 ;
        RECT 180.850 15.060 196.810 15.200 ;
        RECT 180.850 15.000 181.170 15.060 ;
        RECT 196.490 15.000 196.810 15.060 ;
      LAYER via ;
        RECT 196.520 1688.140 196.780 1688.400 ;
        RECT 1223.240 1688.140 1223.500 1688.400 ;
        RECT 180.880 15.000 181.140 15.260 ;
        RECT 196.520 15.000 196.780 15.260 ;
      LAYER met2 ;
        RECT 1223.165 1700.000 1223.445 1704.000 ;
        RECT 1223.300 1688.430 1223.440 1700.000 ;
        RECT 196.520 1688.110 196.780 1688.430 ;
        RECT 1223.240 1688.110 1223.500 1688.430 ;
        RECT 196.580 15.290 196.720 1688.110 ;
        RECT 180.880 14.970 181.140 15.290 ;
        RECT 196.520 14.970 196.780 15.290 ;
        RECT 180.940 2.400 181.080 14.970 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1228.805 897.005 1228.975 904.655 ;
        RECT 1228.805 172.465 1228.975 220.575 ;
      LAYER mcon ;
        RECT 1228.805 904.485 1228.975 904.655 ;
        RECT 1228.805 220.405 1228.975 220.575 ;
      LAYER met1 ;
        RECT 1228.730 904.640 1229.050 904.700 ;
        RECT 1228.535 904.500 1229.050 904.640 ;
        RECT 1228.730 904.440 1229.050 904.500 ;
        RECT 1228.730 897.160 1229.050 897.220 ;
        RECT 1228.535 897.020 1229.050 897.160 ;
        RECT 1228.730 896.960 1229.050 897.020 ;
        RECT 1228.730 752.320 1229.050 752.380 ;
        RECT 1230.570 752.320 1230.890 752.380 ;
        RECT 1228.730 752.180 1230.890 752.320 ;
        RECT 1228.730 752.120 1229.050 752.180 ;
        RECT 1230.570 752.120 1230.890 752.180 ;
        RECT 1228.730 655.760 1229.050 655.820 ;
        RECT 1229.650 655.760 1229.970 655.820 ;
        RECT 1228.730 655.620 1229.970 655.760 ;
        RECT 1228.730 655.560 1229.050 655.620 ;
        RECT 1229.650 655.560 1229.970 655.620 ;
        RECT 1228.730 462.640 1229.050 462.700 ;
        RECT 1229.190 462.640 1229.510 462.700 ;
        RECT 1228.730 462.500 1229.510 462.640 ;
        RECT 1228.730 462.440 1229.050 462.500 ;
        RECT 1229.190 462.440 1229.510 462.500 ;
        RECT 1228.730 366.080 1229.050 366.140 ;
        RECT 1229.190 366.080 1229.510 366.140 ;
        RECT 1228.730 365.940 1229.510 366.080 ;
        RECT 1228.730 365.880 1229.050 365.940 ;
        RECT 1229.190 365.880 1229.510 365.940 ;
        RECT 1228.730 220.560 1229.050 220.620 ;
        RECT 1228.535 220.420 1229.050 220.560 ;
        RECT 1228.730 220.360 1229.050 220.420 ;
        RECT 1228.730 172.620 1229.050 172.680 ;
        RECT 1228.535 172.480 1229.050 172.620 ;
        RECT 1228.730 172.420 1229.050 172.480 ;
        RECT 198.790 19.280 199.110 19.340 ;
        RECT 1190.550 19.280 1190.870 19.340 ;
        RECT 198.790 19.140 1190.870 19.280 ;
        RECT 198.790 19.080 199.110 19.140 ;
        RECT 1190.550 19.080 1190.870 19.140 ;
      LAYER via ;
        RECT 1228.760 904.440 1229.020 904.700 ;
        RECT 1228.760 896.960 1229.020 897.220 ;
        RECT 1228.760 752.120 1229.020 752.380 ;
        RECT 1230.600 752.120 1230.860 752.380 ;
        RECT 1228.760 655.560 1229.020 655.820 ;
        RECT 1229.680 655.560 1229.940 655.820 ;
        RECT 1228.760 462.440 1229.020 462.700 ;
        RECT 1229.220 462.440 1229.480 462.700 ;
        RECT 1228.760 365.880 1229.020 366.140 ;
        RECT 1229.220 365.880 1229.480 366.140 ;
        RECT 1228.760 220.360 1229.020 220.620 ;
        RECT 1228.760 172.420 1229.020 172.680 ;
        RECT 198.820 19.080 199.080 19.340 ;
        RECT 1190.580 19.080 1190.840 19.340 ;
      LAYER met2 ;
        RECT 1230.525 1700.410 1230.805 1704.000 ;
        RECT 1228.820 1700.270 1230.805 1700.410 ;
        RECT 1228.820 904.730 1228.960 1700.270 ;
        RECT 1230.525 1700.000 1230.805 1700.270 ;
        RECT 1228.760 904.410 1229.020 904.730 ;
        RECT 1228.760 896.930 1229.020 897.250 ;
        RECT 1228.820 800.205 1228.960 896.930 ;
        RECT 1228.750 799.835 1229.030 800.205 ;
        RECT 1230.590 799.835 1230.870 800.205 ;
        RECT 1230.660 752.410 1230.800 799.835 ;
        RECT 1228.760 752.090 1229.020 752.410 ;
        RECT 1230.600 752.090 1230.860 752.410 ;
        RECT 1228.820 703.645 1228.960 752.090 ;
        RECT 1228.750 703.275 1229.030 703.645 ;
        RECT 1229.670 703.275 1229.950 703.645 ;
        RECT 1229.740 655.850 1229.880 703.275 ;
        RECT 1228.760 655.530 1229.020 655.850 ;
        RECT 1229.680 655.530 1229.940 655.850 ;
        RECT 1228.820 510.410 1228.960 655.530 ;
        RECT 1228.820 510.270 1229.420 510.410 ;
        RECT 1229.280 462.730 1229.420 510.270 ;
        RECT 1228.760 462.410 1229.020 462.730 ;
        RECT 1229.220 462.410 1229.480 462.730 ;
        RECT 1228.820 413.850 1228.960 462.410 ;
        RECT 1228.820 413.710 1229.420 413.850 ;
        RECT 1229.280 366.170 1229.420 413.710 ;
        RECT 1228.760 365.850 1229.020 366.170 ;
        RECT 1229.220 365.850 1229.480 366.170 ;
        RECT 1228.820 220.650 1228.960 365.850 ;
        RECT 1228.760 220.330 1229.020 220.650 ;
        RECT 1228.760 172.390 1229.020 172.710 ;
        RECT 1228.820 27.725 1228.960 172.390 ;
        RECT 1228.750 27.355 1229.030 27.725 ;
        RECT 1190.570 26.675 1190.850 27.045 ;
        RECT 1190.640 19.370 1190.780 26.675 ;
        RECT 198.820 19.050 199.080 19.370 ;
        RECT 1190.580 19.050 1190.840 19.370 ;
        RECT 198.880 2.400 199.020 19.050 ;
        RECT 198.670 -4.800 199.230 2.400 ;
      LAYER via2 ;
        RECT 1228.750 799.880 1229.030 800.160 ;
        RECT 1230.590 799.880 1230.870 800.160 ;
        RECT 1228.750 703.320 1229.030 703.600 ;
        RECT 1229.670 703.320 1229.950 703.600 ;
        RECT 1228.750 27.400 1229.030 27.680 ;
        RECT 1190.570 26.720 1190.850 27.000 ;
      LAYER met3 ;
        RECT 1228.725 800.170 1229.055 800.185 ;
        RECT 1230.565 800.170 1230.895 800.185 ;
        RECT 1228.725 799.870 1230.895 800.170 ;
        RECT 1228.725 799.855 1229.055 799.870 ;
        RECT 1230.565 799.855 1230.895 799.870 ;
        RECT 1228.725 703.610 1229.055 703.625 ;
        RECT 1229.645 703.610 1229.975 703.625 ;
        RECT 1228.725 703.310 1229.975 703.610 ;
        RECT 1228.725 703.295 1229.055 703.310 ;
        RECT 1229.645 703.295 1229.975 703.310 ;
        RECT 1228.725 27.690 1229.055 27.705 ;
        RECT 1228.725 27.390 1229.730 27.690 ;
        RECT 1228.725 27.375 1229.055 27.390 ;
        RECT 1190.545 27.010 1190.875 27.025 ;
        RECT 1229.430 27.010 1229.730 27.390 ;
        RECT 1190.545 26.710 1229.730 27.010 ;
        RECT 1190.545 26.695 1190.875 26.710 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 306.890 1689.360 307.210 1689.420 ;
        RECT 1237.930 1689.360 1238.250 1689.420 ;
        RECT 306.890 1689.220 1238.250 1689.360 ;
        RECT 306.890 1689.160 307.210 1689.220 ;
        RECT 1237.930 1689.160 1238.250 1689.220 ;
        RECT 216.730 16.220 217.050 16.280 ;
        RECT 306.890 16.220 307.210 16.280 ;
        RECT 216.730 16.080 307.210 16.220 ;
        RECT 216.730 16.020 217.050 16.080 ;
        RECT 306.890 16.020 307.210 16.080 ;
      LAYER via ;
        RECT 306.920 1689.160 307.180 1689.420 ;
        RECT 1237.960 1689.160 1238.220 1689.420 ;
        RECT 216.760 16.020 217.020 16.280 ;
        RECT 306.920 16.020 307.180 16.280 ;
      LAYER met2 ;
        RECT 1237.885 1700.000 1238.165 1704.000 ;
        RECT 1238.020 1689.450 1238.160 1700.000 ;
        RECT 306.920 1689.130 307.180 1689.450 ;
        RECT 1237.960 1689.130 1238.220 1689.450 ;
        RECT 306.980 16.310 307.120 1689.130 ;
        RECT 216.760 15.990 217.020 16.310 ;
        RECT 306.920 15.990 307.180 16.310 ;
        RECT 216.820 2.400 216.960 15.990 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 234.670 19.960 234.990 20.020 ;
        RECT 1243.450 19.960 1243.770 20.020 ;
        RECT 234.670 19.820 1243.770 19.960 ;
        RECT 234.670 19.760 234.990 19.820 ;
        RECT 1243.450 19.760 1243.770 19.820 ;
      LAYER via ;
        RECT 234.700 19.760 234.960 20.020 ;
        RECT 1243.480 19.760 1243.740 20.020 ;
      LAYER met2 ;
        RECT 1245.245 1700.410 1245.525 1704.000 ;
        RECT 1243.540 1700.270 1245.525 1700.410 ;
        RECT 1243.540 20.050 1243.680 1700.270 ;
        RECT 1245.245 1700.000 1245.525 1700.270 ;
        RECT 234.700 19.730 234.960 20.050 ;
        RECT 1243.480 19.730 1243.740 20.050 ;
        RECT 234.760 2.400 234.900 19.730 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 99.890 1687.320 100.210 1687.380 ;
        RECT 1171.690 1687.320 1172.010 1687.380 ;
        RECT 99.890 1687.180 1172.010 1687.320 ;
        RECT 99.890 1687.120 100.210 1687.180 ;
        RECT 1171.690 1687.120 1172.010 1687.180 ;
        RECT 56.190 17.920 56.510 17.980 ;
        RECT 99.890 17.920 100.210 17.980 ;
        RECT 56.190 17.780 100.210 17.920 ;
        RECT 56.190 17.720 56.510 17.780 ;
        RECT 99.890 17.720 100.210 17.780 ;
      LAYER via ;
        RECT 99.920 1687.120 100.180 1687.380 ;
        RECT 1171.720 1687.120 1171.980 1687.380 ;
        RECT 56.220 17.720 56.480 17.980 ;
        RECT 99.920 17.720 100.180 17.980 ;
      LAYER met2 ;
        RECT 1171.645 1700.000 1171.925 1704.000 ;
        RECT 1171.780 1687.410 1171.920 1700.000 ;
        RECT 99.920 1687.090 100.180 1687.410 ;
        RECT 1171.720 1687.090 1171.980 1687.410 ;
        RECT 99.980 18.010 100.120 1687.090 ;
        RECT 56.220 17.690 56.480 18.010 ;
        RECT 99.920 17.690 100.180 18.010 ;
        RECT 56.280 2.400 56.420 17.690 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1181.425 1545.725 1181.595 1593.835 ;
        RECT 1181.425 1449.165 1181.595 1497.275 ;
        RECT 1181.425 1352.605 1181.595 1400.715 ;
        RECT 1181.425 1256.045 1181.595 1304.155 ;
        RECT 1181.425 386.325 1181.595 434.775 ;
        RECT 1181.425 289.765 1181.595 337.875 ;
        RECT 1181.425 193.205 1181.595 241.315 ;
      LAYER mcon ;
        RECT 1181.425 1593.665 1181.595 1593.835 ;
        RECT 1181.425 1497.105 1181.595 1497.275 ;
        RECT 1181.425 1400.545 1181.595 1400.715 ;
        RECT 1181.425 1303.985 1181.595 1304.155 ;
        RECT 1181.425 434.605 1181.595 434.775 ;
        RECT 1181.425 337.705 1181.595 337.875 ;
        RECT 1181.425 241.145 1181.595 241.315 ;
      LAYER met1 ;
        RECT 1181.350 1593.820 1181.670 1593.880 ;
        RECT 1181.155 1593.680 1181.670 1593.820 ;
        RECT 1181.350 1593.620 1181.670 1593.680 ;
        RECT 1181.350 1545.880 1181.670 1545.940 ;
        RECT 1181.155 1545.740 1181.670 1545.880 ;
        RECT 1181.350 1545.680 1181.670 1545.740 ;
        RECT 1181.350 1497.260 1181.670 1497.320 ;
        RECT 1181.155 1497.120 1181.670 1497.260 ;
        RECT 1181.350 1497.060 1181.670 1497.120 ;
        RECT 1181.350 1449.320 1181.670 1449.380 ;
        RECT 1181.155 1449.180 1181.670 1449.320 ;
        RECT 1181.350 1449.120 1181.670 1449.180 ;
        RECT 1181.350 1400.700 1181.670 1400.760 ;
        RECT 1181.155 1400.560 1181.670 1400.700 ;
        RECT 1181.350 1400.500 1181.670 1400.560 ;
        RECT 1181.350 1352.760 1181.670 1352.820 ;
        RECT 1181.155 1352.620 1181.670 1352.760 ;
        RECT 1181.350 1352.560 1181.670 1352.620 ;
        RECT 1181.350 1304.140 1181.670 1304.200 ;
        RECT 1181.155 1304.000 1181.670 1304.140 ;
        RECT 1181.350 1303.940 1181.670 1304.000 ;
        RECT 1181.350 1256.200 1181.670 1256.260 ;
        RECT 1181.155 1256.060 1181.670 1256.200 ;
        RECT 1181.350 1256.000 1181.670 1256.060 ;
        RECT 1181.350 1159.300 1181.670 1159.360 ;
        RECT 1182.270 1159.300 1182.590 1159.360 ;
        RECT 1181.350 1159.160 1182.590 1159.300 ;
        RECT 1181.350 1159.100 1181.670 1159.160 ;
        RECT 1182.270 1159.100 1182.590 1159.160 ;
        RECT 1181.350 1062.740 1181.670 1062.800 ;
        RECT 1182.270 1062.740 1182.590 1062.800 ;
        RECT 1181.350 1062.600 1182.590 1062.740 ;
        RECT 1181.350 1062.540 1181.670 1062.600 ;
        RECT 1182.270 1062.540 1182.590 1062.600 ;
        RECT 1181.350 966.180 1181.670 966.240 ;
        RECT 1182.270 966.180 1182.590 966.240 ;
        RECT 1181.350 966.040 1182.590 966.180 ;
        RECT 1181.350 965.980 1181.670 966.040 ;
        RECT 1182.270 965.980 1182.590 966.040 ;
        RECT 1181.350 869.620 1181.670 869.680 ;
        RECT 1182.270 869.620 1182.590 869.680 ;
        RECT 1181.350 869.480 1182.590 869.620 ;
        RECT 1181.350 869.420 1181.670 869.480 ;
        RECT 1182.270 869.420 1182.590 869.480 ;
        RECT 1181.350 821.000 1181.670 821.060 ;
        RECT 1182.270 821.000 1182.590 821.060 ;
        RECT 1181.350 820.860 1182.590 821.000 ;
        RECT 1181.350 820.800 1181.670 820.860 ;
        RECT 1182.270 820.800 1182.590 820.860 ;
        RECT 1181.350 627.880 1181.670 627.940 ;
        RECT 1182.270 627.880 1182.590 627.940 ;
        RECT 1181.350 627.740 1182.590 627.880 ;
        RECT 1181.350 627.680 1181.670 627.740 ;
        RECT 1182.270 627.680 1182.590 627.740 ;
        RECT 1181.350 531.320 1181.670 531.380 ;
        RECT 1182.270 531.320 1182.590 531.380 ;
        RECT 1181.350 531.180 1182.590 531.320 ;
        RECT 1181.350 531.120 1181.670 531.180 ;
        RECT 1182.270 531.120 1182.590 531.180 ;
        RECT 1181.350 434.760 1181.670 434.820 ;
        RECT 1181.155 434.620 1181.670 434.760 ;
        RECT 1181.350 434.560 1181.670 434.620 ;
        RECT 1181.350 386.480 1181.670 386.540 ;
        RECT 1181.155 386.340 1181.670 386.480 ;
        RECT 1181.350 386.280 1181.670 386.340 ;
        RECT 1181.350 337.860 1181.670 337.920 ;
        RECT 1181.155 337.720 1181.670 337.860 ;
        RECT 1181.350 337.660 1181.670 337.720 ;
        RECT 1181.350 289.920 1181.670 289.980 ;
        RECT 1181.155 289.780 1181.670 289.920 ;
        RECT 1181.350 289.720 1181.670 289.780 ;
        RECT 1181.350 241.300 1181.670 241.360 ;
        RECT 1181.155 241.160 1181.670 241.300 ;
        RECT 1181.350 241.100 1181.670 241.160 ;
        RECT 1181.350 193.360 1181.670 193.420 ;
        RECT 1181.155 193.220 1181.670 193.360 ;
        RECT 1181.350 193.160 1181.670 193.220 ;
        RECT 80.110 17.240 80.430 17.300 ;
        RECT 1181.350 17.240 1181.670 17.300 ;
        RECT 80.110 17.100 1181.670 17.240 ;
        RECT 80.110 17.040 80.430 17.100 ;
        RECT 1181.350 17.040 1181.670 17.100 ;
      LAYER via ;
        RECT 1181.380 1593.620 1181.640 1593.880 ;
        RECT 1181.380 1545.680 1181.640 1545.940 ;
        RECT 1181.380 1497.060 1181.640 1497.320 ;
        RECT 1181.380 1449.120 1181.640 1449.380 ;
        RECT 1181.380 1400.500 1181.640 1400.760 ;
        RECT 1181.380 1352.560 1181.640 1352.820 ;
        RECT 1181.380 1303.940 1181.640 1304.200 ;
        RECT 1181.380 1256.000 1181.640 1256.260 ;
        RECT 1181.380 1159.100 1181.640 1159.360 ;
        RECT 1182.300 1159.100 1182.560 1159.360 ;
        RECT 1181.380 1062.540 1181.640 1062.800 ;
        RECT 1182.300 1062.540 1182.560 1062.800 ;
        RECT 1181.380 965.980 1181.640 966.240 ;
        RECT 1182.300 965.980 1182.560 966.240 ;
        RECT 1181.380 869.420 1181.640 869.680 ;
        RECT 1182.300 869.420 1182.560 869.680 ;
        RECT 1181.380 820.800 1181.640 821.060 ;
        RECT 1182.300 820.800 1182.560 821.060 ;
        RECT 1181.380 627.680 1181.640 627.940 ;
        RECT 1182.300 627.680 1182.560 627.940 ;
        RECT 1181.380 531.120 1181.640 531.380 ;
        RECT 1182.300 531.120 1182.560 531.380 ;
        RECT 1181.380 434.560 1181.640 434.820 ;
        RECT 1181.380 386.280 1181.640 386.540 ;
        RECT 1181.380 337.660 1181.640 337.920 ;
        RECT 1181.380 289.720 1181.640 289.980 ;
        RECT 1181.380 241.100 1181.640 241.360 ;
        RECT 1181.380 193.160 1181.640 193.420 ;
        RECT 80.140 17.040 80.400 17.300 ;
        RECT 1181.380 17.040 1181.640 17.300 ;
      LAYER met2 ;
        RECT 1181.765 1700.410 1182.045 1704.000 ;
        RECT 1181.765 1700.270 1182.500 1700.410 ;
        RECT 1181.765 1700.000 1182.045 1700.270 ;
        RECT 1182.360 1607.930 1182.500 1700.270 ;
        RECT 1181.440 1607.790 1182.500 1607.930 ;
        RECT 1181.440 1593.910 1181.580 1607.790 ;
        RECT 1181.380 1593.590 1181.640 1593.910 ;
        RECT 1181.380 1545.650 1181.640 1545.970 ;
        RECT 1181.440 1497.350 1181.580 1545.650 ;
        RECT 1181.380 1497.030 1181.640 1497.350 ;
        RECT 1181.380 1449.090 1181.640 1449.410 ;
        RECT 1181.440 1400.790 1181.580 1449.090 ;
        RECT 1181.380 1400.470 1181.640 1400.790 ;
        RECT 1181.380 1352.530 1181.640 1352.850 ;
        RECT 1181.440 1304.230 1181.580 1352.530 ;
        RECT 1181.380 1303.910 1181.640 1304.230 ;
        RECT 1181.380 1255.970 1181.640 1256.290 ;
        RECT 1181.440 1207.525 1181.580 1255.970 ;
        RECT 1181.370 1207.155 1181.650 1207.525 ;
        RECT 1182.290 1207.155 1182.570 1207.525 ;
        RECT 1182.360 1159.390 1182.500 1207.155 ;
        RECT 1181.380 1159.070 1181.640 1159.390 ;
        RECT 1182.300 1159.070 1182.560 1159.390 ;
        RECT 1181.440 1110.965 1181.580 1159.070 ;
        RECT 1181.370 1110.595 1181.650 1110.965 ;
        RECT 1182.290 1110.595 1182.570 1110.965 ;
        RECT 1182.360 1062.830 1182.500 1110.595 ;
        RECT 1181.380 1062.510 1181.640 1062.830 ;
        RECT 1182.300 1062.510 1182.560 1062.830 ;
        RECT 1181.440 1014.405 1181.580 1062.510 ;
        RECT 1181.370 1014.035 1181.650 1014.405 ;
        RECT 1182.290 1014.035 1182.570 1014.405 ;
        RECT 1182.360 966.270 1182.500 1014.035 ;
        RECT 1181.380 965.950 1181.640 966.270 ;
        RECT 1182.300 965.950 1182.560 966.270 ;
        RECT 1181.440 917.845 1181.580 965.950 ;
        RECT 1181.370 917.475 1181.650 917.845 ;
        RECT 1182.290 917.475 1182.570 917.845 ;
        RECT 1182.360 869.710 1182.500 917.475 ;
        RECT 1181.380 869.390 1181.640 869.710 ;
        RECT 1182.300 869.390 1182.560 869.710 ;
        RECT 1181.440 821.090 1181.580 869.390 ;
        RECT 1181.380 820.770 1181.640 821.090 ;
        RECT 1182.300 820.770 1182.560 821.090 ;
        RECT 1182.360 773.005 1182.500 820.770 ;
        RECT 1181.370 772.635 1181.650 773.005 ;
        RECT 1182.290 772.635 1182.570 773.005 ;
        RECT 1181.440 738.210 1181.580 772.635 ;
        RECT 1181.440 738.070 1182.500 738.210 ;
        RECT 1182.360 676.445 1182.500 738.070 ;
        RECT 1181.370 676.075 1181.650 676.445 ;
        RECT 1182.290 676.075 1182.570 676.445 ;
        RECT 1181.440 627.970 1181.580 676.075 ;
        RECT 1181.380 627.650 1181.640 627.970 ;
        RECT 1182.300 627.650 1182.560 627.970 ;
        RECT 1182.360 579.885 1182.500 627.650 ;
        RECT 1181.370 579.515 1181.650 579.885 ;
        RECT 1182.290 579.515 1182.570 579.885 ;
        RECT 1181.440 531.410 1181.580 579.515 ;
        RECT 1181.380 531.090 1181.640 531.410 ;
        RECT 1182.300 531.090 1182.560 531.410 ;
        RECT 1182.360 483.325 1182.500 531.090 ;
        RECT 1181.370 482.955 1181.650 483.325 ;
        RECT 1182.290 482.955 1182.570 483.325 ;
        RECT 1181.440 434.850 1181.580 482.955 ;
        RECT 1181.380 434.530 1181.640 434.850 ;
        RECT 1181.380 386.250 1181.640 386.570 ;
        RECT 1181.440 337.950 1181.580 386.250 ;
        RECT 1181.380 337.630 1181.640 337.950 ;
        RECT 1181.380 289.690 1181.640 290.010 ;
        RECT 1181.440 241.390 1181.580 289.690 ;
        RECT 1181.380 241.070 1181.640 241.390 ;
        RECT 1181.380 193.130 1181.640 193.450 ;
        RECT 1181.440 158.170 1181.580 193.130 ;
        RECT 1181.440 158.030 1182.040 158.170 ;
        RECT 1181.900 62.290 1182.040 158.030 ;
        RECT 1181.900 62.150 1182.500 62.290 ;
        RECT 1182.360 61.610 1182.500 62.150 ;
        RECT 1181.440 61.470 1182.500 61.610 ;
        RECT 1181.440 17.330 1181.580 61.470 ;
        RECT 80.140 17.010 80.400 17.330 ;
        RECT 1181.380 17.010 1181.640 17.330 ;
        RECT 80.200 2.400 80.340 17.010 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 1181.370 1207.200 1181.650 1207.480 ;
        RECT 1182.290 1207.200 1182.570 1207.480 ;
        RECT 1181.370 1110.640 1181.650 1110.920 ;
        RECT 1182.290 1110.640 1182.570 1110.920 ;
        RECT 1181.370 1014.080 1181.650 1014.360 ;
        RECT 1182.290 1014.080 1182.570 1014.360 ;
        RECT 1181.370 917.520 1181.650 917.800 ;
        RECT 1182.290 917.520 1182.570 917.800 ;
        RECT 1181.370 772.680 1181.650 772.960 ;
        RECT 1182.290 772.680 1182.570 772.960 ;
        RECT 1181.370 676.120 1181.650 676.400 ;
        RECT 1182.290 676.120 1182.570 676.400 ;
        RECT 1181.370 579.560 1181.650 579.840 ;
        RECT 1182.290 579.560 1182.570 579.840 ;
        RECT 1181.370 483.000 1181.650 483.280 ;
        RECT 1182.290 483.000 1182.570 483.280 ;
      LAYER met3 ;
        RECT 1181.345 1207.490 1181.675 1207.505 ;
        RECT 1182.265 1207.490 1182.595 1207.505 ;
        RECT 1181.345 1207.190 1182.595 1207.490 ;
        RECT 1181.345 1207.175 1181.675 1207.190 ;
        RECT 1182.265 1207.175 1182.595 1207.190 ;
        RECT 1181.345 1110.930 1181.675 1110.945 ;
        RECT 1182.265 1110.930 1182.595 1110.945 ;
        RECT 1181.345 1110.630 1182.595 1110.930 ;
        RECT 1181.345 1110.615 1181.675 1110.630 ;
        RECT 1182.265 1110.615 1182.595 1110.630 ;
        RECT 1181.345 1014.370 1181.675 1014.385 ;
        RECT 1182.265 1014.370 1182.595 1014.385 ;
        RECT 1181.345 1014.070 1182.595 1014.370 ;
        RECT 1181.345 1014.055 1181.675 1014.070 ;
        RECT 1182.265 1014.055 1182.595 1014.070 ;
        RECT 1181.345 917.810 1181.675 917.825 ;
        RECT 1182.265 917.810 1182.595 917.825 ;
        RECT 1181.345 917.510 1182.595 917.810 ;
        RECT 1181.345 917.495 1181.675 917.510 ;
        RECT 1182.265 917.495 1182.595 917.510 ;
        RECT 1181.345 772.970 1181.675 772.985 ;
        RECT 1182.265 772.970 1182.595 772.985 ;
        RECT 1181.345 772.670 1182.595 772.970 ;
        RECT 1181.345 772.655 1181.675 772.670 ;
        RECT 1182.265 772.655 1182.595 772.670 ;
        RECT 1181.345 676.410 1181.675 676.425 ;
        RECT 1182.265 676.410 1182.595 676.425 ;
        RECT 1181.345 676.110 1182.595 676.410 ;
        RECT 1181.345 676.095 1181.675 676.110 ;
        RECT 1182.265 676.095 1182.595 676.110 ;
        RECT 1181.345 579.850 1181.675 579.865 ;
        RECT 1182.265 579.850 1182.595 579.865 ;
        RECT 1181.345 579.550 1182.595 579.850 ;
        RECT 1181.345 579.535 1181.675 579.550 ;
        RECT 1182.265 579.535 1182.595 579.550 ;
        RECT 1181.345 483.290 1181.675 483.305 ;
        RECT 1182.265 483.290 1182.595 483.305 ;
        RECT 1181.345 482.990 1182.595 483.290 ;
        RECT 1181.345 482.975 1181.675 482.990 ;
        RECT 1182.265 482.975 1182.595 482.990 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 175.790 1688.680 176.110 1688.740 ;
        RECT 1191.470 1688.680 1191.790 1688.740 ;
        RECT 175.790 1688.540 1191.790 1688.680 ;
        RECT 175.790 1688.480 176.110 1688.540 ;
        RECT 1191.470 1688.480 1191.790 1688.540 ;
        RECT 103.570 18.940 103.890 19.000 ;
        RECT 175.790 18.940 176.110 19.000 ;
        RECT 103.570 18.800 176.110 18.940 ;
        RECT 103.570 18.740 103.890 18.800 ;
        RECT 175.790 18.740 176.110 18.800 ;
      LAYER via ;
        RECT 175.820 1688.480 176.080 1688.740 ;
        RECT 1191.500 1688.480 1191.760 1688.740 ;
        RECT 103.600 18.740 103.860 19.000 ;
        RECT 175.820 18.740 176.080 19.000 ;
      LAYER met2 ;
        RECT 1191.425 1700.000 1191.705 1704.000 ;
        RECT 1191.560 1688.770 1191.700 1700.000 ;
        RECT 175.820 1688.450 176.080 1688.770 ;
        RECT 1191.500 1688.450 1191.760 1688.770 ;
        RECT 175.880 19.030 176.020 1688.450 ;
        RECT 103.600 18.710 103.860 19.030 ;
        RECT 175.820 18.710 176.080 19.030 ;
        RECT 103.660 2.400 103.800 18.710 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 127.490 17.920 127.810 17.980 ;
        RECT 1201.590 17.920 1201.910 17.980 ;
        RECT 127.490 17.780 1201.910 17.920 ;
        RECT 127.490 17.720 127.810 17.780 ;
        RECT 1201.590 17.720 1201.910 17.780 ;
      LAYER via ;
        RECT 127.520 17.720 127.780 17.980 ;
        RECT 1201.620 17.720 1201.880 17.980 ;
      LAYER met2 ;
        RECT 1201.085 1700.410 1201.365 1704.000 ;
        RECT 1201.085 1700.270 1201.820 1700.410 ;
        RECT 1201.085 1700.000 1201.365 1700.270 ;
        RECT 1201.680 18.010 1201.820 1700.270 ;
        RECT 127.520 17.690 127.780 18.010 ;
        RECT 1201.620 17.690 1201.880 18.010 ;
        RECT 127.580 2.400 127.720 17.690 ;
        RECT 127.370 -4.800 127.930 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 51.590 17.240 51.910 17.300 ;
        RECT 26.290 17.100 51.910 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 51.590 17.040 51.910 17.100 ;
      LAYER via ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 51.620 17.040 51.880 17.300 ;
      LAYER met2 ;
        RECT 1159.685 1700.000 1159.965 1704.000 ;
        RECT 1159.820 1686.925 1159.960 1700.000 ;
        RECT 51.610 1686.555 51.890 1686.925 ;
        RECT 1159.750 1686.555 1160.030 1686.925 ;
        RECT 51.680 17.330 51.820 1686.555 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 51.620 17.010 51.880 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 26.170 -4.800 26.730 2.400 ;
      LAYER via2 ;
        RECT 51.610 1686.600 51.890 1686.880 ;
        RECT 1159.750 1686.600 1160.030 1686.880 ;
      LAYER met3 ;
        RECT 51.585 1686.890 51.915 1686.905 ;
        RECT 1159.725 1686.890 1160.055 1686.905 ;
        RECT 51.585 1686.590 1160.055 1686.890 ;
        RECT 51.585 1686.575 51.915 1686.590 ;
        RECT 1159.725 1686.575 1160.055 1686.590 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1161.985 1700.410 1162.265 1704.000 ;
        RECT 1160.280 1700.270 1162.265 1700.410 ;
        RECT 1160.280 16.845 1160.420 1700.270 ;
        RECT 1161.985 1700.000 1162.265 1700.270 ;
        RECT 32.290 16.475 32.570 16.845 ;
        RECT 1160.210 16.475 1160.490 16.845 ;
        RECT 32.360 2.400 32.500 16.475 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 32.290 16.520 32.570 16.800 ;
        RECT 1160.210 16.520 1160.490 16.800 ;
      LAYER met3 ;
        RECT 32.265 16.810 32.595 16.825 ;
        RECT 1160.185 16.810 1160.515 16.825 ;
        RECT 32.265 16.510 1160.515 16.810 ;
        RECT 32.265 16.495 32.595 16.510 ;
        RECT 1160.185 16.495 1160.515 16.510 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.320 7.020 3529.000 ;
        RECT 184.020 -9.320 187.020 3529.000 ;
        RECT 364.020 -9.320 367.020 3529.000 ;
        RECT 544.020 -9.320 547.020 3529.000 ;
        RECT 724.020 -9.320 727.020 3529.000 ;
        RECT 904.020 -9.320 907.020 3529.000 ;
        RECT 1084.020 -9.320 1087.020 3529.000 ;
        RECT 1264.020 -9.320 1267.020 3529.000 ;
        RECT 1444.020 -9.320 1447.020 3529.000 ;
        RECT 1624.020 -9.320 1627.020 3529.000 ;
        RECT 1804.020 -9.320 1807.020 3529.000 ;
        RECT 1984.020 -9.320 1987.020 3529.000 ;
        RECT 2164.020 -9.320 2167.020 3529.000 ;
        RECT 2344.020 -9.320 2347.020 3529.000 ;
        RECT 2524.020 -9.320 2527.020 3529.000 ;
        RECT 2704.020 -9.320 2707.020 3529.000 ;
        RECT 2884.020 -9.320 2887.020 3529.000 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.680 3429.380 2934.300 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.680 3249.380 2934.300 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.680 3069.380 2934.300 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.680 2889.380 2934.300 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.680 2709.380 2934.300 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.680 2529.380 2934.300 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.680 2349.380 2934.300 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.680 2169.380 2934.300 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.680 1989.380 2934.300 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.680 1809.380 2934.300 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.680 1629.380 2934.300 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.680 1449.380 2934.300 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.680 1269.380 2934.300 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.680 1089.380 2934.300 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.680 909.380 2934.300 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.680 729.380 2934.300 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.680 549.380 2934.300 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.680 369.380 2934.300 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.680 189.380 2934.300 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.680 9.380 2934.300 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
        RECT 94.020 -9.320 97.020 3529.000 ;
        RECT 274.020 -9.320 277.020 3529.000 ;
        RECT 454.020 -9.320 457.020 3529.000 ;
        RECT 634.020 -9.320 637.020 3529.000 ;
        RECT 814.020 -9.320 817.020 3529.000 ;
        RECT 994.020 -9.320 997.020 3529.000 ;
        RECT 1174.020 -9.320 1177.020 3529.000 ;
        RECT 1354.020 -9.320 1357.020 3529.000 ;
        RECT 1534.020 -9.320 1537.020 3529.000 ;
        RECT 1714.020 -9.320 1717.020 3529.000 ;
        RECT 1894.020 -9.320 1897.020 3529.000 ;
        RECT 2074.020 -9.320 2077.020 3529.000 ;
        RECT 2254.020 -9.320 2257.020 3529.000 ;
        RECT 2434.020 -9.320 2437.020 3529.000 ;
        RECT 2614.020 -9.320 2617.020 3529.000 ;
        RECT 2794.020 -9.320 2797.020 3529.000 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
      LAYER via4 ;
        RECT -13.770 3527.710 -12.590 3528.890 ;
        RECT -13.770 3526.110 -12.590 3527.290 ;
        RECT -13.770 3341.090 -12.590 3342.270 ;
        RECT -13.770 3339.490 -12.590 3340.670 ;
        RECT -13.770 3161.090 -12.590 3162.270 ;
        RECT -13.770 3159.490 -12.590 3160.670 ;
        RECT -13.770 2981.090 -12.590 2982.270 ;
        RECT -13.770 2979.490 -12.590 2980.670 ;
        RECT -13.770 2801.090 -12.590 2802.270 ;
        RECT -13.770 2799.490 -12.590 2800.670 ;
        RECT -13.770 2621.090 -12.590 2622.270 ;
        RECT -13.770 2619.490 -12.590 2620.670 ;
        RECT -13.770 2441.090 -12.590 2442.270 ;
        RECT -13.770 2439.490 -12.590 2440.670 ;
        RECT -13.770 2261.090 -12.590 2262.270 ;
        RECT -13.770 2259.490 -12.590 2260.670 ;
        RECT -13.770 2081.090 -12.590 2082.270 ;
        RECT -13.770 2079.490 -12.590 2080.670 ;
        RECT -13.770 1901.090 -12.590 1902.270 ;
        RECT -13.770 1899.490 -12.590 1900.670 ;
        RECT -13.770 1721.090 -12.590 1722.270 ;
        RECT -13.770 1719.490 -12.590 1720.670 ;
        RECT -13.770 1541.090 -12.590 1542.270 ;
        RECT -13.770 1539.490 -12.590 1540.670 ;
        RECT -13.770 1361.090 -12.590 1362.270 ;
        RECT -13.770 1359.490 -12.590 1360.670 ;
        RECT -13.770 1181.090 -12.590 1182.270 ;
        RECT -13.770 1179.490 -12.590 1180.670 ;
        RECT -13.770 1001.090 -12.590 1002.270 ;
        RECT -13.770 999.490 -12.590 1000.670 ;
        RECT -13.770 821.090 -12.590 822.270 ;
        RECT -13.770 819.490 -12.590 820.670 ;
        RECT -13.770 641.090 -12.590 642.270 ;
        RECT -13.770 639.490 -12.590 640.670 ;
        RECT -13.770 461.090 -12.590 462.270 ;
        RECT -13.770 459.490 -12.590 460.670 ;
        RECT -13.770 281.090 -12.590 282.270 ;
        RECT -13.770 279.490 -12.590 280.670 ;
        RECT -13.770 101.090 -12.590 102.270 ;
        RECT -13.770 99.490 -12.590 100.670 ;
        RECT -13.770 -7.610 -12.590 -6.430 ;
        RECT -13.770 -9.210 -12.590 -8.030 ;
        RECT 94.930 3527.710 96.110 3528.890 ;
        RECT 94.930 3526.110 96.110 3527.290 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.610 96.110 -6.430 ;
        RECT 94.930 -9.210 96.110 -8.030 ;
        RECT 274.930 3527.710 276.110 3528.890 ;
        RECT 274.930 3526.110 276.110 3527.290 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.610 276.110 -6.430 ;
        RECT 274.930 -9.210 276.110 -8.030 ;
        RECT 454.930 3527.710 456.110 3528.890 ;
        RECT 454.930 3526.110 456.110 3527.290 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.610 456.110 -6.430 ;
        RECT 454.930 -9.210 456.110 -8.030 ;
        RECT 634.930 3527.710 636.110 3528.890 ;
        RECT 634.930 3526.110 636.110 3527.290 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.610 636.110 -6.430 ;
        RECT 634.930 -9.210 636.110 -8.030 ;
        RECT 814.930 3527.710 816.110 3528.890 ;
        RECT 814.930 3526.110 816.110 3527.290 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.610 816.110 -6.430 ;
        RECT 814.930 -9.210 816.110 -8.030 ;
        RECT 994.930 3527.710 996.110 3528.890 ;
        RECT 994.930 3526.110 996.110 3527.290 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.610 996.110 -6.430 ;
        RECT 994.930 -9.210 996.110 -8.030 ;
        RECT 1174.930 3527.710 1176.110 3528.890 ;
        RECT 1174.930 3526.110 1176.110 3527.290 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.610 1176.110 -6.430 ;
        RECT 1174.930 -9.210 1176.110 -8.030 ;
        RECT 1354.930 3527.710 1356.110 3528.890 ;
        RECT 1354.930 3526.110 1356.110 3527.290 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.610 1356.110 -6.430 ;
        RECT 1354.930 -9.210 1356.110 -8.030 ;
        RECT 1534.930 3527.710 1536.110 3528.890 ;
        RECT 1534.930 3526.110 1536.110 3527.290 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.610 1536.110 -6.430 ;
        RECT 1534.930 -9.210 1536.110 -8.030 ;
        RECT 1714.930 3527.710 1716.110 3528.890 ;
        RECT 1714.930 3526.110 1716.110 3527.290 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.610 1716.110 -6.430 ;
        RECT 1714.930 -9.210 1716.110 -8.030 ;
        RECT 1894.930 3527.710 1896.110 3528.890 ;
        RECT 1894.930 3526.110 1896.110 3527.290 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.610 1896.110 -6.430 ;
        RECT 1894.930 -9.210 1896.110 -8.030 ;
        RECT 2074.930 3527.710 2076.110 3528.890 ;
        RECT 2074.930 3526.110 2076.110 3527.290 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.610 2076.110 -6.430 ;
        RECT 2074.930 -9.210 2076.110 -8.030 ;
        RECT 2254.930 3527.710 2256.110 3528.890 ;
        RECT 2254.930 3526.110 2256.110 3527.290 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.610 2256.110 -6.430 ;
        RECT 2254.930 -9.210 2256.110 -8.030 ;
        RECT 2434.930 3527.710 2436.110 3528.890 ;
        RECT 2434.930 3526.110 2436.110 3527.290 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.610 2436.110 -6.430 ;
        RECT 2434.930 -9.210 2436.110 -8.030 ;
        RECT 2614.930 3527.710 2616.110 3528.890 ;
        RECT 2614.930 3526.110 2616.110 3527.290 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.610 2616.110 -6.430 ;
        RECT 2614.930 -9.210 2616.110 -8.030 ;
        RECT 2794.930 3527.710 2796.110 3528.890 ;
        RECT 2794.930 3526.110 2796.110 3527.290 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.610 2796.110 -6.430 ;
        RECT 2794.930 -9.210 2796.110 -8.030 ;
        RECT 2932.210 3527.710 2933.390 3528.890 ;
        RECT 2932.210 3526.110 2933.390 3527.290 ;
        RECT 2932.210 3341.090 2933.390 3342.270 ;
        RECT 2932.210 3339.490 2933.390 3340.670 ;
        RECT 2932.210 3161.090 2933.390 3162.270 ;
        RECT 2932.210 3159.490 2933.390 3160.670 ;
        RECT 2932.210 2981.090 2933.390 2982.270 ;
        RECT 2932.210 2979.490 2933.390 2980.670 ;
        RECT 2932.210 2801.090 2933.390 2802.270 ;
        RECT 2932.210 2799.490 2933.390 2800.670 ;
        RECT 2932.210 2621.090 2933.390 2622.270 ;
        RECT 2932.210 2619.490 2933.390 2620.670 ;
        RECT 2932.210 2441.090 2933.390 2442.270 ;
        RECT 2932.210 2439.490 2933.390 2440.670 ;
        RECT 2932.210 2261.090 2933.390 2262.270 ;
        RECT 2932.210 2259.490 2933.390 2260.670 ;
        RECT 2932.210 2081.090 2933.390 2082.270 ;
        RECT 2932.210 2079.490 2933.390 2080.670 ;
        RECT 2932.210 1901.090 2933.390 1902.270 ;
        RECT 2932.210 1899.490 2933.390 1900.670 ;
        RECT 2932.210 1721.090 2933.390 1722.270 ;
        RECT 2932.210 1719.490 2933.390 1720.670 ;
        RECT 2932.210 1541.090 2933.390 1542.270 ;
        RECT 2932.210 1539.490 2933.390 1540.670 ;
        RECT 2932.210 1361.090 2933.390 1362.270 ;
        RECT 2932.210 1359.490 2933.390 1360.670 ;
        RECT 2932.210 1181.090 2933.390 1182.270 ;
        RECT 2932.210 1179.490 2933.390 1180.670 ;
        RECT 2932.210 1001.090 2933.390 1002.270 ;
        RECT 2932.210 999.490 2933.390 1000.670 ;
        RECT 2932.210 821.090 2933.390 822.270 ;
        RECT 2932.210 819.490 2933.390 820.670 ;
        RECT 2932.210 641.090 2933.390 642.270 ;
        RECT 2932.210 639.490 2933.390 640.670 ;
        RECT 2932.210 461.090 2933.390 462.270 ;
        RECT 2932.210 459.490 2933.390 460.670 ;
        RECT 2932.210 281.090 2933.390 282.270 ;
        RECT 2932.210 279.490 2933.390 280.670 ;
        RECT 2932.210 101.090 2933.390 102.270 ;
        RECT 2932.210 99.490 2933.390 100.670 ;
        RECT 2932.210 -7.610 2933.390 -6.430 ;
        RECT 2932.210 -9.210 2933.390 -8.030 ;
      LAYER met5 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 94.020 3529.000 97.020 3529.010 ;
        RECT 274.020 3529.000 277.020 3529.010 ;
        RECT 454.020 3529.000 457.020 3529.010 ;
        RECT 634.020 3529.000 637.020 3529.010 ;
        RECT 814.020 3529.000 817.020 3529.010 ;
        RECT 994.020 3529.000 997.020 3529.010 ;
        RECT 1174.020 3529.000 1177.020 3529.010 ;
        RECT 1354.020 3529.000 1357.020 3529.010 ;
        RECT 1534.020 3529.000 1537.020 3529.010 ;
        RECT 1714.020 3529.000 1717.020 3529.010 ;
        RECT 1894.020 3529.000 1897.020 3529.010 ;
        RECT 2074.020 3529.000 2077.020 3529.010 ;
        RECT 2254.020 3529.000 2257.020 3529.010 ;
        RECT 2434.020 3529.000 2437.020 3529.010 ;
        RECT 2614.020 3529.000 2617.020 3529.010 ;
        RECT 2794.020 3529.000 2797.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 94.020 3525.990 97.020 3526.000 ;
        RECT 274.020 3525.990 277.020 3526.000 ;
        RECT 454.020 3525.990 457.020 3526.000 ;
        RECT 634.020 3525.990 637.020 3526.000 ;
        RECT 814.020 3525.990 817.020 3526.000 ;
        RECT 994.020 3525.990 997.020 3526.000 ;
        RECT 1174.020 3525.990 1177.020 3526.000 ;
        RECT 1354.020 3525.990 1357.020 3526.000 ;
        RECT 1534.020 3525.990 1537.020 3526.000 ;
        RECT 1714.020 3525.990 1717.020 3526.000 ;
        RECT 1894.020 3525.990 1897.020 3526.000 ;
        RECT 2074.020 3525.990 2077.020 3526.000 ;
        RECT 2254.020 3525.990 2257.020 3526.000 ;
        RECT 2434.020 3525.990 2437.020 3526.000 ;
        RECT 2614.020 3525.990 2617.020 3526.000 ;
        RECT 2794.020 3525.990 2797.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -14.680 3342.380 -11.680 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.300 3342.380 2934.300 3342.390 ;
        RECT -14.680 3339.380 2934.300 3342.380 ;
        RECT -14.680 3339.370 -11.680 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.300 3339.370 2934.300 3339.380 ;
        RECT -14.680 3162.380 -11.680 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.300 3162.380 2934.300 3162.390 ;
        RECT -14.680 3159.380 2934.300 3162.380 ;
        RECT -14.680 3159.370 -11.680 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.300 3159.370 2934.300 3159.380 ;
        RECT -14.680 2982.380 -11.680 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.300 2982.380 2934.300 2982.390 ;
        RECT -14.680 2979.380 2934.300 2982.380 ;
        RECT -14.680 2979.370 -11.680 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.300 2979.370 2934.300 2979.380 ;
        RECT -14.680 2802.380 -11.680 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.300 2802.380 2934.300 2802.390 ;
        RECT -14.680 2799.380 2934.300 2802.380 ;
        RECT -14.680 2799.370 -11.680 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.300 2799.370 2934.300 2799.380 ;
        RECT -14.680 2622.380 -11.680 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.300 2622.380 2934.300 2622.390 ;
        RECT -14.680 2619.380 2934.300 2622.380 ;
        RECT -14.680 2619.370 -11.680 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.300 2619.370 2934.300 2619.380 ;
        RECT -14.680 2442.380 -11.680 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.300 2442.380 2934.300 2442.390 ;
        RECT -14.680 2439.380 2934.300 2442.380 ;
        RECT -14.680 2439.370 -11.680 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.300 2439.370 2934.300 2439.380 ;
        RECT -14.680 2262.380 -11.680 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.300 2262.380 2934.300 2262.390 ;
        RECT -14.680 2259.380 2934.300 2262.380 ;
        RECT -14.680 2259.370 -11.680 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.300 2259.370 2934.300 2259.380 ;
        RECT -14.680 2082.380 -11.680 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.300 2082.380 2934.300 2082.390 ;
        RECT -14.680 2079.380 2934.300 2082.380 ;
        RECT -14.680 2079.370 -11.680 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.300 2079.370 2934.300 2079.380 ;
        RECT -14.680 1902.380 -11.680 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.300 1902.380 2934.300 1902.390 ;
        RECT -14.680 1899.380 2934.300 1902.380 ;
        RECT -14.680 1899.370 -11.680 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.300 1899.370 2934.300 1899.380 ;
        RECT -14.680 1722.380 -11.680 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.300 1722.380 2934.300 1722.390 ;
        RECT -14.680 1719.380 2934.300 1722.380 ;
        RECT -14.680 1719.370 -11.680 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.300 1719.370 2934.300 1719.380 ;
        RECT -14.680 1542.380 -11.680 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.300 1542.380 2934.300 1542.390 ;
        RECT -14.680 1539.380 2934.300 1542.380 ;
        RECT -14.680 1539.370 -11.680 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.300 1539.370 2934.300 1539.380 ;
        RECT -14.680 1362.380 -11.680 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.300 1362.380 2934.300 1362.390 ;
        RECT -14.680 1359.380 2934.300 1362.380 ;
        RECT -14.680 1359.370 -11.680 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.300 1359.370 2934.300 1359.380 ;
        RECT -14.680 1182.380 -11.680 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.300 1182.380 2934.300 1182.390 ;
        RECT -14.680 1179.380 2934.300 1182.380 ;
        RECT -14.680 1179.370 -11.680 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.300 1179.370 2934.300 1179.380 ;
        RECT -14.680 1002.380 -11.680 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.300 1002.380 2934.300 1002.390 ;
        RECT -14.680 999.380 2934.300 1002.380 ;
        RECT -14.680 999.370 -11.680 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.300 999.370 2934.300 999.380 ;
        RECT -14.680 822.380 -11.680 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.300 822.380 2934.300 822.390 ;
        RECT -14.680 819.380 2934.300 822.380 ;
        RECT -14.680 819.370 -11.680 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.300 819.370 2934.300 819.380 ;
        RECT -14.680 642.380 -11.680 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.300 642.380 2934.300 642.390 ;
        RECT -14.680 639.380 2934.300 642.380 ;
        RECT -14.680 639.370 -11.680 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.300 639.370 2934.300 639.380 ;
        RECT -14.680 462.380 -11.680 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.300 462.380 2934.300 462.390 ;
        RECT -14.680 459.380 2934.300 462.380 ;
        RECT -14.680 459.370 -11.680 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.300 459.370 2934.300 459.380 ;
        RECT -14.680 282.380 -11.680 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.300 282.380 2934.300 282.390 ;
        RECT -14.680 279.380 2934.300 282.380 ;
        RECT -14.680 279.370 -11.680 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.300 279.370 2934.300 279.380 ;
        RECT -14.680 102.380 -11.680 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.300 102.380 2934.300 102.390 ;
        RECT -14.680 99.380 2934.300 102.380 ;
        RECT -14.680 99.370 -11.680 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.300 99.370 2934.300 99.380 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 94.020 -6.320 97.020 -6.310 ;
        RECT 274.020 -6.320 277.020 -6.310 ;
        RECT 454.020 -6.320 457.020 -6.310 ;
        RECT 634.020 -6.320 637.020 -6.310 ;
        RECT 814.020 -6.320 817.020 -6.310 ;
        RECT 994.020 -6.320 997.020 -6.310 ;
        RECT 1174.020 -6.320 1177.020 -6.310 ;
        RECT 1354.020 -6.320 1357.020 -6.310 ;
        RECT 1534.020 -6.320 1537.020 -6.310 ;
        RECT 1714.020 -6.320 1717.020 -6.310 ;
        RECT 1894.020 -6.320 1897.020 -6.310 ;
        RECT 2074.020 -6.320 2077.020 -6.310 ;
        RECT 2254.020 -6.320 2257.020 -6.310 ;
        RECT 2434.020 -6.320 2437.020 -6.310 ;
        RECT 2614.020 -6.320 2617.020 -6.310 ;
        RECT 2794.020 -6.320 2797.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 94.020 -9.330 97.020 -9.320 ;
        RECT 274.020 -9.330 277.020 -9.320 ;
        RECT 454.020 -9.330 457.020 -9.320 ;
        RECT 634.020 -9.330 637.020 -9.320 ;
        RECT 814.020 -9.330 817.020 -9.320 ;
        RECT 994.020 -9.330 997.020 -9.320 ;
        RECT 1174.020 -9.330 1177.020 -9.320 ;
        RECT 1354.020 -9.330 1357.020 -9.320 ;
        RECT 1534.020 -9.330 1537.020 -9.320 ;
        RECT 1714.020 -9.330 1717.020 -9.320 ;
        RECT 1894.020 -9.330 1897.020 -9.320 ;
        RECT 2074.020 -9.330 2077.020 -9.320 ;
        RECT 2254.020 -9.330 2257.020 -9.320 ;
        RECT 2434.020 -9.330 2437.020 -9.320 ;
        RECT 2614.020 -9.330 2617.020 -9.320 ;
        RECT 2794.020 -9.330 2797.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
        RECT 22.020 -18.720 25.020 3538.400 ;
        RECT 202.020 -18.720 205.020 3538.400 ;
        RECT 382.020 -18.720 385.020 3538.400 ;
        RECT 562.020 -18.720 565.020 3538.400 ;
        RECT 742.020 -18.720 745.020 3538.400 ;
        RECT 922.020 -18.720 925.020 3538.400 ;
        RECT 1102.020 -18.720 1105.020 3538.400 ;
        RECT 1282.020 -18.720 1285.020 3538.400 ;
        RECT 1462.020 -18.720 1465.020 3538.400 ;
        RECT 1642.020 -18.720 1645.020 3538.400 ;
        RECT 1822.020 -18.720 1825.020 3538.400 ;
        RECT 2002.020 -18.720 2005.020 3538.400 ;
        RECT 2182.020 -18.720 2185.020 3538.400 ;
        RECT 2362.020 -18.720 2365.020 3538.400 ;
        RECT 2542.020 -18.720 2545.020 3538.400 ;
        RECT 2722.020 -18.720 2725.020 3538.400 ;
        RECT 2902.020 -18.720 2905.020 3538.400 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
      LAYER via4 ;
        RECT -18.470 3532.410 -17.290 3533.590 ;
        RECT -18.470 3530.810 -17.290 3531.990 ;
        RECT -18.470 3449.090 -17.290 3450.270 ;
        RECT -18.470 3447.490 -17.290 3448.670 ;
        RECT -18.470 3269.090 -17.290 3270.270 ;
        RECT -18.470 3267.490 -17.290 3268.670 ;
        RECT -18.470 3089.090 -17.290 3090.270 ;
        RECT -18.470 3087.490 -17.290 3088.670 ;
        RECT -18.470 2909.090 -17.290 2910.270 ;
        RECT -18.470 2907.490 -17.290 2908.670 ;
        RECT -18.470 2729.090 -17.290 2730.270 ;
        RECT -18.470 2727.490 -17.290 2728.670 ;
        RECT -18.470 2549.090 -17.290 2550.270 ;
        RECT -18.470 2547.490 -17.290 2548.670 ;
        RECT -18.470 2369.090 -17.290 2370.270 ;
        RECT -18.470 2367.490 -17.290 2368.670 ;
        RECT -18.470 2189.090 -17.290 2190.270 ;
        RECT -18.470 2187.490 -17.290 2188.670 ;
        RECT -18.470 2009.090 -17.290 2010.270 ;
        RECT -18.470 2007.490 -17.290 2008.670 ;
        RECT -18.470 1829.090 -17.290 1830.270 ;
        RECT -18.470 1827.490 -17.290 1828.670 ;
        RECT -18.470 1649.090 -17.290 1650.270 ;
        RECT -18.470 1647.490 -17.290 1648.670 ;
        RECT -18.470 1469.090 -17.290 1470.270 ;
        RECT -18.470 1467.490 -17.290 1468.670 ;
        RECT -18.470 1289.090 -17.290 1290.270 ;
        RECT -18.470 1287.490 -17.290 1288.670 ;
        RECT -18.470 1109.090 -17.290 1110.270 ;
        RECT -18.470 1107.490 -17.290 1108.670 ;
        RECT -18.470 929.090 -17.290 930.270 ;
        RECT -18.470 927.490 -17.290 928.670 ;
        RECT -18.470 749.090 -17.290 750.270 ;
        RECT -18.470 747.490 -17.290 748.670 ;
        RECT -18.470 569.090 -17.290 570.270 ;
        RECT -18.470 567.490 -17.290 568.670 ;
        RECT -18.470 389.090 -17.290 390.270 ;
        RECT -18.470 387.490 -17.290 388.670 ;
        RECT -18.470 209.090 -17.290 210.270 ;
        RECT -18.470 207.490 -17.290 208.670 ;
        RECT -18.470 29.090 -17.290 30.270 ;
        RECT -18.470 27.490 -17.290 28.670 ;
        RECT -18.470 -12.310 -17.290 -11.130 ;
        RECT -18.470 -13.910 -17.290 -12.730 ;
        RECT 22.930 3532.410 24.110 3533.590 ;
        RECT 22.930 3530.810 24.110 3531.990 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.310 24.110 -11.130 ;
        RECT 22.930 -13.910 24.110 -12.730 ;
        RECT 202.930 3532.410 204.110 3533.590 ;
        RECT 202.930 3530.810 204.110 3531.990 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.310 204.110 -11.130 ;
        RECT 202.930 -13.910 204.110 -12.730 ;
        RECT 382.930 3532.410 384.110 3533.590 ;
        RECT 382.930 3530.810 384.110 3531.990 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.310 384.110 -11.130 ;
        RECT 382.930 -13.910 384.110 -12.730 ;
        RECT 562.930 3532.410 564.110 3533.590 ;
        RECT 562.930 3530.810 564.110 3531.990 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.310 564.110 -11.130 ;
        RECT 562.930 -13.910 564.110 -12.730 ;
        RECT 742.930 3532.410 744.110 3533.590 ;
        RECT 742.930 3530.810 744.110 3531.990 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.310 744.110 -11.130 ;
        RECT 742.930 -13.910 744.110 -12.730 ;
        RECT 922.930 3532.410 924.110 3533.590 ;
        RECT 922.930 3530.810 924.110 3531.990 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.310 924.110 -11.130 ;
        RECT 922.930 -13.910 924.110 -12.730 ;
        RECT 1102.930 3532.410 1104.110 3533.590 ;
        RECT 1102.930 3530.810 1104.110 3531.990 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.310 1104.110 -11.130 ;
        RECT 1102.930 -13.910 1104.110 -12.730 ;
        RECT 1282.930 3532.410 1284.110 3533.590 ;
        RECT 1282.930 3530.810 1284.110 3531.990 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.310 1284.110 -11.130 ;
        RECT 1282.930 -13.910 1284.110 -12.730 ;
        RECT 1462.930 3532.410 1464.110 3533.590 ;
        RECT 1462.930 3530.810 1464.110 3531.990 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.310 1464.110 -11.130 ;
        RECT 1462.930 -13.910 1464.110 -12.730 ;
        RECT 1642.930 3532.410 1644.110 3533.590 ;
        RECT 1642.930 3530.810 1644.110 3531.990 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.310 1644.110 -11.130 ;
        RECT 1642.930 -13.910 1644.110 -12.730 ;
        RECT 1822.930 3532.410 1824.110 3533.590 ;
        RECT 1822.930 3530.810 1824.110 3531.990 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.310 1824.110 -11.130 ;
        RECT 1822.930 -13.910 1824.110 -12.730 ;
        RECT 2002.930 3532.410 2004.110 3533.590 ;
        RECT 2002.930 3530.810 2004.110 3531.990 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.310 2004.110 -11.130 ;
        RECT 2002.930 -13.910 2004.110 -12.730 ;
        RECT 2182.930 3532.410 2184.110 3533.590 ;
        RECT 2182.930 3530.810 2184.110 3531.990 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.310 2184.110 -11.130 ;
        RECT 2182.930 -13.910 2184.110 -12.730 ;
        RECT 2362.930 3532.410 2364.110 3533.590 ;
        RECT 2362.930 3530.810 2364.110 3531.990 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.310 2364.110 -11.130 ;
        RECT 2362.930 -13.910 2364.110 -12.730 ;
        RECT 2542.930 3532.410 2544.110 3533.590 ;
        RECT 2542.930 3530.810 2544.110 3531.990 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.310 2544.110 -11.130 ;
        RECT 2542.930 -13.910 2544.110 -12.730 ;
        RECT 2722.930 3532.410 2724.110 3533.590 ;
        RECT 2722.930 3530.810 2724.110 3531.990 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.310 2724.110 -11.130 ;
        RECT 2722.930 -13.910 2724.110 -12.730 ;
        RECT 2902.930 3532.410 2904.110 3533.590 ;
        RECT 2902.930 3530.810 2904.110 3531.990 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.310 2904.110 -11.130 ;
        RECT 2902.930 -13.910 2904.110 -12.730 ;
        RECT 2936.910 3532.410 2938.090 3533.590 ;
        RECT 2936.910 3530.810 2938.090 3531.990 ;
        RECT 2936.910 3449.090 2938.090 3450.270 ;
        RECT 2936.910 3447.490 2938.090 3448.670 ;
        RECT 2936.910 3269.090 2938.090 3270.270 ;
        RECT 2936.910 3267.490 2938.090 3268.670 ;
        RECT 2936.910 3089.090 2938.090 3090.270 ;
        RECT 2936.910 3087.490 2938.090 3088.670 ;
        RECT 2936.910 2909.090 2938.090 2910.270 ;
        RECT 2936.910 2907.490 2938.090 2908.670 ;
        RECT 2936.910 2729.090 2938.090 2730.270 ;
        RECT 2936.910 2727.490 2938.090 2728.670 ;
        RECT 2936.910 2549.090 2938.090 2550.270 ;
        RECT 2936.910 2547.490 2938.090 2548.670 ;
        RECT 2936.910 2369.090 2938.090 2370.270 ;
        RECT 2936.910 2367.490 2938.090 2368.670 ;
        RECT 2936.910 2189.090 2938.090 2190.270 ;
        RECT 2936.910 2187.490 2938.090 2188.670 ;
        RECT 2936.910 2009.090 2938.090 2010.270 ;
        RECT 2936.910 2007.490 2938.090 2008.670 ;
        RECT 2936.910 1829.090 2938.090 1830.270 ;
        RECT 2936.910 1827.490 2938.090 1828.670 ;
        RECT 2936.910 1649.090 2938.090 1650.270 ;
        RECT 2936.910 1647.490 2938.090 1648.670 ;
        RECT 2936.910 1469.090 2938.090 1470.270 ;
        RECT 2936.910 1467.490 2938.090 1468.670 ;
        RECT 2936.910 1289.090 2938.090 1290.270 ;
        RECT 2936.910 1287.490 2938.090 1288.670 ;
        RECT 2936.910 1109.090 2938.090 1110.270 ;
        RECT 2936.910 1107.490 2938.090 1108.670 ;
        RECT 2936.910 929.090 2938.090 930.270 ;
        RECT 2936.910 927.490 2938.090 928.670 ;
        RECT 2936.910 749.090 2938.090 750.270 ;
        RECT 2936.910 747.490 2938.090 748.670 ;
        RECT 2936.910 569.090 2938.090 570.270 ;
        RECT 2936.910 567.490 2938.090 568.670 ;
        RECT 2936.910 389.090 2938.090 390.270 ;
        RECT 2936.910 387.490 2938.090 388.670 ;
        RECT 2936.910 209.090 2938.090 210.270 ;
        RECT 2936.910 207.490 2938.090 208.670 ;
        RECT 2936.910 29.090 2938.090 30.270 ;
        RECT 2936.910 27.490 2938.090 28.670 ;
        RECT 2936.910 -12.310 2938.090 -11.130 ;
        RECT 2936.910 -13.910 2938.090 -12.730 ;
      LAYER met5 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 22.020 3533.700 25.020 3533.710 ;
        RECT 202.020 3533.700 205.020 3533.710 ;
        RECT 382.020 3533.700 385.020 3533.710 ;
        RECT 562.020 3533.700 565.020 3533.710 ;
        RECT 742.020 3533.700 745.020 3533.710 ;
        RECT 922.020 3533.700 925.020 3533.710 ;
        RECT 1102.020 3533.700 1105.020 3533.710 ;
        RECT 1282.020 3533.700 1285.020 3533.710 ;
        RECT 1462.020 3533.700 1465.020 3533.710 ;
        RECT 1642.020 3533.700 1645.020 3533.710 ;
        RECT 1822.020 3533.700 1825.020 3533.710 ;
        RECT 2002.020 3533.700 2005.020 3533.710 ;
        RECT 2182.020 3533.700 2185.020 3533.710 ;
        RECT 2362.020 3533.700 2365.020 3533.710 ;
        RECT 2542.020 3533.700 2545.020 3533.710 ;
        RECT 2722.020 3533.700 2725.020 3533.710 ;
        RECT 2902.020 3533.700 2905.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 22.020 3530.690 25.020 3530.700 ;
        RECT 202.020 3530.690 205.020 3530.700 ;
        RECT 382.020 3530.690 385.020 3530.700 ;
        RECT 562.020 3530.690 565.020 3530.700 ;
        RECT 742.020 3530.690 745.020 3530.700 ;
        RECT 922.020 3530.690 925.020 3530.700 ;
        RECT 1102.020 3530.690 1105.020 3530.700 ;
        RECT 1282.020 3530.690 1285.020 3530.700 ;
        RECT 1462.020 3530.690 1465.020 3530.700 ;
        RECT 1642.020 3530.690 1645.020 3530.700 ;
        RECT 1822.020 3530.690 1825.020 3530.700 ;
        RECT 2002.020 3530.690 2005.020 3530.700 ;
        RECT 2182.020 3530.690 2185.020 3530.700 ;
        RECT 2362.020 3530.690 2365.020 3530.700 ;
        RECT 2542.020 3530.690 2545.020 3530.700 ;
        RECT 2722.020 3530.690 2725.020 3530.700 ;
        RECT 2902.020 3530.690 2905.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -19.380 3450.380 -16.380 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2936.000 3450.380 2939.000 3450.390 ;
        RECT -24.080 3447.380 2943.700 3450.380 ;
        RECT -19.380 3447.370 -16.380 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2936.000 3447.370 2939.000 3447.380 ;
        RECT -19.380 3270.380 -16.380 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2936.000 3270.380 2939.000 3270.390 ;
        RECT -24.080 3267.380 2943.700 3270.380 ;
        RECT -19.380 3267.370 -16.380 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2936.000 3267.370 2939.000 3267.380 ;
        RECT -19.380 3090.380 -16.380 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2936.000 3090.380 2939.000 3090.390 ;
        RECT -24.080 3087.380 2943.700 3090.380 ;
        RECT -19.380 3087.370 -16.380 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2936.000 3087.370 2939.000 3087.380 ;
        RECT -19.380 2910.380 -16.380 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2936.000 2910.380 2939.000 2910.390 ;
        RECT -24.080 2907.380 2943.700 2910.380 ;
        RECT -19.380 2907.370 -16.380 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2936.000 2907.370 2939.000 2907.380 ;
        RECT -19.380 2730.380 -16.380 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2936.000 2730.380 2939.000 2730.390 ;
        RECT -24.080 2727.380 2943.700 2730.380 ;
        RECT -19.380 2727.370 -16.380 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2936.000 2727.370 2939.000 2727.380 ;
        RECT -19.380 2550.380 -16.380 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2936.000 2550.380 2939.000 2550.390 ;
        RECT -24.080 2547.380 2943.700 2550.380 ;
        RECT -19.380 2547.370 -16.380 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2936.000 2547.370 2939.000 2547.380 ;
        RECT -19.380 2370.380 -16.380 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2936.000 2370.380 2939.000 2370.390 ;
        RECT -24.080 2367.380 2943.700 2370.380 ;
        RECT -19.380 2367.370 -16.380 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2936.000 2367.370 2939.000 2367.380 ;
        RECT -19.380 2190.380 -16.380 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2936.000 2190.380 2939.000 2190.390 ;
        RECT -24.080 2187.380 2943.700 2190.380 ;
        RECT -19.380 2187.370 -16.380 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2936.000 2187.370 2939.000 2187.380 ;
        RECT -19.380 2010.380 -16.380 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2936.000 2010.380 2939.000 2010.390 ;
        RECT -24.080 2007.380 2943.700 2010.380 ;
        RECT -19.380 2007.370 -16.380 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2936.000 2007.370 2939.000 2007.380 ;
        RECT -19.380 1830.380 -16.380 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2936.000 1830.380 2939.000 1830.390 ;
        RECT -24.080 1827.380 2943.700 1830.380 ;
        RECT -19.380 1827.370 -16.380 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2936.000 1827.370 2939.000 1827.380 ;
        RECT -19.380 1650.380 -16.380 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2936.000 1650.380 2939.000 1650.390 ;
        RECT -24.080 1647.380 2943.700 1650.380 ;
        RECT -19.380 1647.370 -16.380 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2936.000 1647.370 2939.000 1647.380 ;
        RECT -19.380 1470.380 -16.380 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2936.000 1470.380 2939.000 1470.390 ;
        RECT -24.080 1467.380 2943.700 1470.380 ;
        RECT -19.380 1467.370 -16.380 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2936.000 1467.370 2939.000 1467.380 ;
        RECT -19.380 1290.380 -16.380 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2936.000 1290.380 2939.000 1290.390 ;
        RECT -24.080 1287.380 2943.700 1290.380 ;
        RECT -19.380 1287.370 -16.380 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2936.000 1287.370 2939.000 1287.380 ;
        RECT -19.380 1110.380 -16.380 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2936.000 1110.380 2939.000 1110.390 ;
        RECT -24.080 1107.380 2943.700 1110.380 ;
        RECT -19.380 1107.370 -16.380 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2936.000 1107.370 2939.000 1107.380 ;
        RECT -19.380 930.380 -16.380 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2936.000 930.380 2939.000 930.390 ;
        RECT -24.080 927.380 2943.700 930.380 ;
        RECT -19.380 927.370 -16.380 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2936.000 927.370 2939.000 927.380 ;
        RECT -19.380 750.380 -16.380 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2936.000 750.380 2939.000 750.390 ;
        RECT -24.080 747.380 2943.700 750.380 ;
        RECT -19.380 747.370 -16.380 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2936.000 747.370 2939.000 747.380 ;
        RECT -19.380 570.380 -16.380 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2936.000 570.380 2939.000 570.390 ;
        RECT -24.080 567.380 2943.700 570.380 ;
        RECT -19.380 567.370 -16.380 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2936.000 567.370 2939.000 567.380 ;
        RECT -19.380 390.380 -16.380 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2936.000 390.380 2939.000 390.390 ;
        RECT -24.080 387.380 2943.700 390.380 ;
        RECT -19.380 387.370 -16.380 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2936.000 387.370 2939.000 387.380 ;
        RECT -19.380 210.380 -16.380 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2936.000 210.380 2939.000 210.390 ;
        RECT -24.080 207.380 2943.700 210.380 ;
        RECT -19.380 207.370 -16.380 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2936.000 207.370 2939.000 207.380 ;
        RECT -19.380 30.380 -16.380 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2936.000 30.380 2939.000 30.390 ;
        RECT -24.080 27.380 2943.700 30.380 ;
        RECT -19.380 27.370 -16.380 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2936.000 27.370 2939.000 27.380 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 22.020 -11.020 25.020 -11.010 ;
        RECT 202.020 -11.020 205.020 -11.010 ;
        RECT 382.020 -11.020 385.020 -11.010 ;
        RECT 562.020 -11.020 565.020 -11.010 ;
        RECT 742.020 -11.020 745.020 -11.010 ;
        RECT 922.020 -11.020 925.020 -11.010 ;
        RECT 1102.020 -11.020 1105.020 -11.010 ;
        RECT 1282.020 -11.020 1285.020 -11.010 ;
        RECT 1462.020 -11.020 1465.020 -11.010 ;
        RECT 1642.020 -11.020 1645.020 -11.010 ;
        RECT 1822.020 -11.020 1825.020 -11.010 ;
        RECT 2002.020 -11.020 2005.020 -11.010 ;
        RECT 2182.020 -11.020 2185.020 -11.010 ;
        RECT 2362.020 -11.020 2365.020 -11.010 ;
        RECT 2542.020 -11.020 2545.020 -11.010 ;
        RECT 2722.020 -11.020 2725.020 -11.010 ;
        RECT 2902.020 -11.020 2905.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 22.020 -14.030 25.020 -14.020 ;
        RECT 202.020 -14.030 205.020 -14.020 ;
        RECT 382.020 -14.030 385.020 -14.020 ;
        RECT 562.020 -14.030 565.020 -14.020 ;
        RECT 742.020 -14.030 745.020 -14.020 ;
        RECT 922.020 -14.030 925.020 -14.020 ;
        RECT 1102.020 -14.030 1105.020 -14.020 ;
        RECT 1282.020 -14.030 1285.020 -14.020 ;
        RECT 1462.020 -14.030 1465.020 -14.020 ;
        RECT 1642.020 -14.030 1645.020 -14.020 ;
        RECT 1822.020 -14.030 1825.020 -14.020 ;
        RECT 2002.020 -14.030 2005.020 -14.020 ;
        RECT 2182.020 -14.030 2185.020 -14.020 ;
        RECT 2362.020 -14.030 2365.020 -14.020 ;
        RECT 2542.020 -14.030 2545.020 -14.020 ;
        RECT 2722.020 -14.030 2725.020 -14.020 ;
        RECT 2902.020 -14.030 2905.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
        RECT 112.020 -18.720 115.020 3538.400 ;
        RECT 292.020 -18.720 295.020 3538.400 ;
        RECT 472.020 -18.720 475.020 3538.400 ;
        RECT 652.020 -18.720 655.020 3538.400 ;
        RECT 832.020 -18.720 835.020 3538.400 ;
        RECT 1012.020 -18.720 1015.020 3538.400 ;
        RECT 1192.020 -18.720 1195.020 3538.400 ;
        RECT 1372.020 -18.720 1375.020 3538.400 ;
        RECT 1552.020 -18.720 1555.020 3538.400 ;
        RECT 1732.020 -18.720 1735.020 3538.400 ;
        RECT 1912.020 -18.720 1915.020 3538.400 ;
        RECT 2092.020 -18.720 2095.020 3538.400 ;
        RECT 2272.020 -18.720 2275.020 3538.400 ;
        RECT 2452.020 -18.720 2455.020 3538.400 ;
        RECT 2632.020 -18.720 2635.020 3538.400 ;
        RECT 2812.020 -18.720 2815.020 3538.400 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
      LAYER via4 ;
        RECT -23.170 3537.110 -21.990 3538.290 ;
        RECT -23.170 3535.510 -21.990 3536.690 ;
        RECT -23.170 3359.090 -21.990 3360.270 ;
        RECT -23.170 3357.490 -21.990 3358.670 ;
        RECT -23.170 3179.090 -21.990 3180.270 ;
        RECT -23.170 3177.490 -21.990 3178.670 ;
        RECT -23.170 2999.090 -21.990 3000.270 ;
        RECT -23.170 2997.490 -21.990 2998.670 ;
        RECT -23.170 2819.090 -21.990 2820.270 ;
        RECT -23.170 2817.490 -21.990 2818.670 ;
        RECT -23.170 2639.090 -21.990 2640.270 ;
        RECT -23.170 2637.490 -21.990 2638.670 ;
        RECT -23.170 2459.090 -21.990 2460.270 ;
        RECT -23.170 2457.490 -21.990 2458.670 ;
        RECT -23.170 2279.090 -21.990 2280.270 ;
        RECT -23.170 2277.490 -21.990 2278.670 ;
        RECT -23.170 2099.090 -21.990 2100.270 ;
        RECT -23.170 2097.490 -21.990 2098.670 ;
        RECT -23.170 1919.090 -21.990 1920.270 ;
        RECT -23.170 1917.490 -21.990 1918.670 ;
        RECT -23.170 1739.090 -21.990 1740.270 ;
        RECT -23.170 1737.490 -21.990 1738.670 ;
        RECT -23.170 1559.090 -21.990 1560.270 ;
        RECT -23.170 1557.490 -21.990 1558.670 ;
        RECT -23.170 1379.090 -21.990 1380.270 ;
        RECT -23.170 1377.490 -21.990 1378.670 ;
        RECT -23.170 1199.090 -21.990 1200.270 ;
        RECT -23.170 1197.490 -21.990 1198.670 ;
        RECT -23.170 1019.090 -21.990 1020.270 ;
        RECT -23.170 1017.490 -21.990 1018.670 ;
        RECT -23.170 839.090 -21.990 840.270 ;
        RECT -23.170 837.490 -21.990 838.670 ;
        RECT -23.170 659.090 -21.990 660.270 ;
        RECT -23.170 657.490 -21.990 658.670 ;
        RECT -23.170 479.090 -21.990 480.270 ;
        RECT -23.170 477.490 -21.990 478.670 ;
        RECT -23.170 299.090 -21.990 300.270 ;
        RECT -23.170 297.490 -21.990 298.670 ;
        RECT -23.170 119.090 -21.990 120.270 ;
        RECT -23.170 117.490 -21.990 118.670 ;
        RECT -23.170 -17.010 -21.990 -15.830 ;
        RECT -23.170 -18.610 -21.990 -17.430 ;
        RECT 112.930 3537.110 114.110 3538.290 ;
        RECT 112.930 3535.510 114.110 3536.690 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -17.010 114.110 -15.830 ;
        RECT 112.930 -18.610 114.110 -17.430 ;
        RECT 292.930 3537.110 294.110 3538.290 ;
        RECT 292.930 3535.510 294.110 3536.690 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -17.010 294.110 -15.830 ;
        RECT 292.930 -18.610 294.110 -17.430 ;
        RECT 472.930 3537.110 474.110 3538.290 ;
        RECT 472.930 3535.510 474.110 3536.690 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -17.010 474.110 -15.830 ;
        RECT 472.930 -18.610 474.110 -17.430 ;
        RECT 652.930 3537.110 654.110 3538.290 ;
        RECT 652.930 3535.510 654.110 3536.690 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -17.010 654.110 -15.830 ;
        RECT 652.930 -18.610 654.110 -17.430 ;
        RECT 832.930 3537.110 834.110 3538.290 ;
        RECT 832.930 3535.510 834.110 3536.690 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -17.010 834.110 -15.830 ;
        RECT 832.930 -18.610 834.110 -17.430 ;
        RECT 1012.930 3537.110 1014.110 3538.290 ;
        RECT 1012.930 3535.510 1014.110 3536.690 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -17.010 1014.110 -15.830 ;
        RECT 1012.930 -18.610 1014.110 -17.430 ;
        RECT 1192.930 3537.110 1194.110 3538.290 ;
        RECT 1192.930 3535.510 1194.110 3536.690 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -17.010 1194.110 -15.830 ;
        RECT 1192.930 -18.610 1194.110 -17.430 ;
        RECT 1372.930 3537.110 1374.110 3538.290 ;
        RECT 1372.930 3535.510 1374.110 3536.690 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -17.010 1374.110 -15.830 ;
        RECT 1372.930 -18.610 1374.110 -17.430 ;
        RECT 1552.930 3537.110 1554.110 3538.290 ;
        RECT 1552.930 3535.510 1554.110 3536.690 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -17.010 1554.110 -15.830 ;
        RECT 1552.930 -18.610 1554.110 -17.430 ;
        RECT 1732.930 3537.110 1734.110 3538.290 ;
        RECT 1732.930 3535.510 1734.110 3536.690 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -17.010 1734.110 -15.830 ;
        RECT 1732.930 -18.610 1734.110 -17.430 ;
        RECT 1912.930 3537.110 1914.110 3538.290 ;
        RECT 1912.930 3535.510 1914.110 3536.690 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -17.010 1914.110 -15.830 ;
        RECT 1912.930 -18.610 1914.110 -17.430 ;
        RECT 2092.930 3537.110 2094.110 3538.290 ;
        RECT 2092.930 3535.510 2094.110 3536.690 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -17.010 2094.110 -15.830 ;
        RECT 2092.930 -18.610 2094.110 -17.430 ;
        RECT 2272.930 3537.110 2274.110 3538.290 ;
        RECT 2272.930 3535.510 2274.110 3536.690 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -17.010 2274.110 -15.830 ;
        RECT 2272.930 -18.610 2274.110 -17.430 ;
        RECT 2452.930 3537.110 2454.110 3538.290 ;
        RECT 2452.930 3535.510 2454.110 3536.690 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -17.010 2454.110 -15.830 ;
        RECT 2452.930 -18.610 2454.110 -17.430 ;
        RECT 2632.930 3537.110 2634.110 3538.290 ;
        RECT 2632.930 3535.510 2634.110 3536.690 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -17.010 2634.110 -15.830 ;
        RECT 2632.930 -18.610 2634.110 -17.430 ;
        RECT 2812.930 3537.110 2814.110 3538.290 ;
        RECT 2812.930 3535.510 2814.110 3536.690 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -17.010 2814.110 -15.830 ;
        RECT 2812.930 -18.610 2814.110 -17.430 ;
        RECT 2941.610 3537.110 2942.790 3538.290 ;
        RECT 2941.610 3535.510 2942.790 3536.690 ;
        RECT 2941.610 3359.090 2942.790 3360.270 ;
        RECT 2941.610 3357.490 2942.790 3358.670 ;
        RECT 2941.610 3179.090 2942.790 3180.270 ;
        RECT 2941.610 3177.490 2942.790 3178.670 ;
        RECT 2941.610 2999.090 2942.790 3000.270 ;
        RECT 2941.610 2997.490 2942.790 2998.670 ;
        RECT 2941.610 2819.090 2942.790 2820.270 ;
        RECT 2941.610 2817.490 2942.790 2818.670 ;
        RECT 2941.610 2639.090 2942.790 2640.270 ;
        RECT 2941.610 2637.490 2942.790 2638.670 ;
        RECT 2941.610 2459.090 2942.790 2460.270 ;
        RECT 2941.610 2457.490 2942.790 2458.670 ;
        RECT 2941.610 2279.090 2942.790 2280.270 ;
        RECT 2941.610 2277.490 2942.790 2278.670 ;
        RECT 2941.610 2099.090 2942.790 2100.270 ;
        RECT 2941.610 2097.490 2942.790 2098.670 ;
        RECT 2941.610 1919.090 2942.790 1920.270 ;
        RECT 2941.610 1917.490 2942.790 1918.670 ;
        RECT 2941.610 1739.090 2942.790 1740.270 ;
        RECT 2941.610 1737.490 2942.790 1738.670 ;
        RECT 2941.610 1559.090 2942.790 1560.270 ;
        RECT 2941.610 1557.490 2942.790 1558.670 ;
        RECT 2941.610 1379.090 2942.790 1380.270 ;
        RECT 2941.610 1377.490 2942.790 1378.670 ;
        RECT 2941.610 1199.090 2942.790 1200.270 ;
        RECT 2941.610 1197.490 2942.790 1198.670 ;
        RECT 2941.610 1019.090 2942.790 1020.270 ;
        RECT 2941.610 1017.490 2942.790 1018.670 ;
        RECT 2941.610 839.090 2942.790 840.270 ;
        RECT 2941.610 837.490 2942.790 838.670 ;
        RECT 2941.610 659.090 2942.790 660.270 ;
        RECT 2941.610 657.490 2942.790 658.670 ;
        RECT 2941.610 479.090 2942.790 480.270 ;
        RECT 2941.610 477.490 2942.790 478.670 ;
        RECT 2941.610 299.090 2942.790 300.270 ;
        RECT 2941.610 297.490 2942.790 298.670 ;
        RECT 2941.610 119.090 2942.790 120.270 ;
        RECT 2941.610 117.490 2942.790 118.670 ;
        RECT 2941.610 -17.010 2942.790 -15.830 ;
        RECT 2941.610 -18.610 2942.790 -17.430 ;
      LAYER met5 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 112.020 3538.400 115.020 3538.410 ;
        RECT 292.020 3538.400 295.020 3538.410 ;
        RECT 472.020 3538.400 475.020 3538.410 ;
        RECT 652.020 3538.400 655.020 3538.410 ;
        RECT 832.020 3538.400 835.020 3538.410 ;
        RECT 1012.020 3538.400 1015.020 3538.410 ;
        RECT 1192.020 3538.400 1195.020 3538.410 ;
        RECT 1372.020 3538.400 1375.020 3538.410 ;
        RECT 1552.020 3538.400 1555.020 3538.410 ;
        RECT 1732.020 3538.400 1735.020 3538.410 ;
        RECT 1912.020 3538.400 1915.020 3538.410 ;
        RECT 2092.020 3538.400 2095.020 3538.410 ;
        RECT 2272.020 3538.400 2275.020 3538.410 ;
        RECT 2452.020 3538.400 2455.020 3538.410 ;
        RECT 2632.020 3538.400 2635.020 3538.410 ;
        RECT 2812.020 3538.400 2815.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 112.020 3535.390 115.020 3535.400 ;
        RECT 292.020 3535.390 295.020 3535.400 ;
        RECT 472.020 3535.390 475.020 3535.400 ;
        RECT 652.020 3535.390 655.020 3535.400 ;
        RECT 832.020 3535.390 835.020 3535.400 ;
        RECT 1012.020 3535.390 1015.020 3535.400 ;
        RECT 1192.020 3535.390 1195.020 3535.400 ;
        RECT 1372.020 3535.390 1375.020 3535.400 ;
        RECT 1552.020 3535.390 1555.020 3535.400 ;
        RECT 1732.020 3535.390 1735.020 3535.400 ;
        RECT 1912.020 3535.390 1915.020 3535.400 ;
        RECT 2092.020 3535.390 2095.020 3535.400 ;
        RECT 2272.020 3535.390 2275.020 3535.400 ;
        RECT 2452.020 3535.390 2455.020 3535.400 ;
        RECT 2632.020 3535.390 2635.020 3535.400 ;
        RECT 2812.020 3535.390 2815.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -24.080 3360.380 -21.080 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.700 3360.380 2943.700 3360.390 ;
        RECT -24.080 3357.380 2943.700 3360.380 ;
        RECT -24.080 3357.370 -21.080 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.700 3357.370 2943.700 3357.380 ;
        RECT -24.080 3180.380 -21.080 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.700 3180.380 2943.700 3180.390 ;
        RECT -24.080 3177.380 2943.700 3180.380 ;
        RECT -24.080 3177.370 -21.080 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.700 3177.370 2943.700 3177.380 ;
        RECT -24.080 3000.380 -21.080 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.700 3000.380 2943.700 3000.390 ;
        RECT -24.080 2997.380 2943.700 3000.380 ;
        RECT -24.080 2997.370 -21.080 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.700 2997.370 2943.700 2997.380 ;
        RECT -24.080 2820.380 -21.080 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.700 2820.380 2943.700 2820.390 ;
        RECT -24.080 2817.380 2943.700 2820.380 ;
        RECT -24.080 2817.370 -21.080 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.700 2817.370 2943.700 2817.380 ;
        RECT -24.080 2640.380 -21.080 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.700 2640.380 2943.700 2640.390 ;
        RECT -24.080 2637.380 2943.700 2640.380 ;
        RECT -24.080 2637.370 -21.080 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.700 2637.370 2943.700 2637.380 ;
        RECT -24.080 2460.380 -21.080 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.700 2460.380 2943.700 2460.390 ;
        RECT -24.080 2457.380 2943.700 2460.380 ;
        RECT -24.080 2457.370 -21.080 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.700 2457.370 2943.700 2457.380 ;
        RECT -24.080 2280.380 -21.080 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.700 2280.380 2943.700 2280.390 ;
        RECT -24.080 2277.380 2943.700 2280.380 ;
        RECT -24.080 2277.370 -21.080 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.700 2277.370 2943.700 2277.380 ;
        RECT -24.080 2100.380 -21.080 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.700 2100.380 2943.700 2100.390 ;
        RECT -24.080 2097.380 2943.700 2100.380 ;
        RECT -24.080 2097.370 -21.080 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.700 2097.370 2943.700 2097.380 ;
        RECT -24.080 1920.380 -21.080 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.700 1920.380 2943.700 1920.390 ;
        RECT -24.080 1917.380 2943.700 1920.380 ;
        RECT -24.080 1917.370 -21.080 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.700 1917.370 2943.700 1917.380 ;
        RECT -24.080 1740.380 -21.080 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.700 1740.380 2943.700 1740.390 ;
        RECT -24.080 1737.380 2943.700 1740.380 ;
        RECT -24.080 1737.370 -21.080 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.700 1737.370 2943.700 1737.380 ;
        RECT -24.080 1560.380 -21.080 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.700 1560.380 2943.700 1560.390 ;
        RECT -24.080 1557.380 2943.700 1560.380 ;
        RECT -24.080 1557.370 -21.080 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.700 1557.370 2943.700 1557.380 ;
        RECT -24.080 1380.380 -21.080 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.700 1380.380 2943.700 1380.390 ;
        RECT -24.080 1377.380 2943.700 1380.380 ;
        RECT -24.080 1377.370 -21.080 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.700 1377.370 2943.700 1377.380 ;
        RECT -24.080 1200.380 -21.080 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.700 1200.380 2943.700 1200.390 ;
        RECT -24.080 1197.380 2943.700 1200.380 ;
        RECT -24.080 1197.370 -21.080 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.700 1197.370 2943.700 1197.380 ;
        RECT -24.080 1020.380 -21.080 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.700 1020.380 2943.700 1020.390 ;
        RECT -24.080 1017.380 2943.700 1020.380 ;
        RECT -24.080 1017.370 -21.080 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.700 1017.370 2943.700 1017.380 ;
        RECT -24.080 840.380 -21.080 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.700 840.380 2943.700 840.390 ;
        RECT -24.080 837.380 2943.700 840.380 ;
        RECT -24.080 837.370 -21.080 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.700 837.370 2943.700 837.380 ;
        RECT -24.080 660.380 -21.080 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.700 660.380 2943.700 660.390 ;
        RECT -24.080 657.380 2943.700 660.380 ;
        RECT -24.080 657.370 -21.080 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.700 657.370 2943.700 657.380 ;
        RECT -24.080 480.380 -21.080 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.700 480.380 2943.700 480.390 ;
        RECT -24.080 477.380 2943.700 480.380 ;
        RECT -24.080 477.370 -21.080 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.700 477.370 2943.700 477.380 ;
        RECT -24.080 300.380 -21.080 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.700 300.380 2943.700 300.390 ;
        RECT -24.080 297.380 2943.700 300.380 ;
        RECT -24.080 297.370 -21.080 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.700 297.370 2943.700 297.380 ;
        RECT -24.080 120.380 -21.080 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.700 120.380 2943.700 120.390 ;
        RECT -24.080 117.380 2943.700 120.380 ;
        RECT -24.080 117.370 -21.080 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.700 117.370 2943.700 117.380 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 112.020 -15.720 115.020 -15.710 ;
        RECT 292.020 -15.720 295.020 -15.710 ;
        RECT 472.020 -15.720 475.020 -15.710 ;
        RECT 652.020 -15.720 655.020 -15.710 ;
        RECT 832.020 -15.720 835.020 -15.710 ;
        RECT 1012.020 -15.720 1015.020 -15.710 ;
        RECT 1192.020 -15.720 1195.020 -15.710 ;
        RECT 1372.020 -15.720 1375.020 -15.710 ;
        RECT 1552.020 -15.720 1555.020 -15.710 ;
        RECT 1732.020 -15.720 1735.020 -15.710 ;
        RECT 1912.020 -15.720 1915.020 -15.710 ;
        RECT 2092.020 -15.720 2095.020 -15.710 ;
        RECT 2272.020 -15.720 2275.020 -15.710 ;
        RECT 2452.020 -15.720 2455.020 -15.710 ;
        RECT 2632.020 -15.720 2635.020 -15.710 ;
        RECT 2812.020 -15.720 2815.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 112.020 -18.730 115.020 -18.720 ;
        RECT 292.020 -18.730 295.020 -18.720 ;
        RECT 472.020 -18.730 475.020 -18.720 ;
        RECT 652.020 -18.730 655.020 -18.720 ;
        RECT 832.020 -18.730 835.020 -18.720 ;
        RECT 1012.020 -18.730 1015.020 -18.720 ;
        RECT 1192.020 -18.730 1195.020 -18.720 ;
        RECT 1372.020 -18.730 1375.020 -18.720 ;
        RECT 1552.020 -18.730 1555.020 -18.720 ;
        RECT 1732.020 -18.730 1735.020 -18.720 ;
        RECT 1912.020 -18.730 1915.020 -18.720 ;
        RECT 2092.020 -18.730 2095.020 -18.720 ;
        RECT 2272.020 -18.730 2275.020 -18.720 ;
        RECT 2452.020 -18.730 2455.020 -18.720 ;
        RECT 2632.020 -18.730 2635.020 -18.720 ;
        RECT 2812.020 -18.730 2815.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
        RECT 40.020 -28.120 43.020 3547.800 ;
        RECT 220.020 -28.120 223.020 3547.800 ;
        RECT 400.020 -28.120 403.020 3547.800 ;
        RECT 580.020 -28.120 583.020 3547.800 ;
        RECT 760.020 -28.120 763.020 3547.800 ;
        RECT 940.020 -28.120 943.020 3547.800 ;
        RECT 1120.020 -28.120 1123.020 3547.800 ;
        RECT 1300.020 -28.120 1303.020 3547.800 ;
        RECT 1480.020 -28.120 1483.020 3547.800 ;
        RECT 1660.020 -28.120 1663.020 3547.800 ;
        RECT 1840.020 -28.120 1843.020 3547.800 ;
        RECT 2020.020 -28.120 2023.020 3547.800 ;
        RECT 2200.020 -28.120 2203.020 3547.800 ;
        RECT 2380.020 -28.120 2383.020 3547.800 ;
        RECT 2560.020 -28.120 2563.020 3547.800 ;
        RECT 2740.020 -28.120 2743.020 3547.800 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
      LAYER via4 ;
        RECT -27.870 3541.810 -26.690 3542.990 ;
        RECT -27.870 3540.210 -26.690 3541.390 ;
        RECT -27.870 3467.090 -26.690 3468.270 ;
        RECT -27.870 3465.490 -26.690 3466.670 ;
        RECT -27.870 3287.090 -26.690 3288.270 ;
        RECT -27.870 3285.490 -26.690 3286.670 ;
        RECT -27.870 3107.090 -26.690 3108.270 ;
        RECT -27.870 3105.490 -26.690 3106.670 ;
        RECT -27.870 2927.090 -26.690 2928.270 ;
        RECT -27.870 2925.490 -26.690 2926.670 ;
        RECT -27.870 2747.090 -26.690 2748.270 ;
        RECT -27.870 2745.490 -26.690 2746.670 ;
        RECT -27.870 2567.090 -26.690 2568.270 ;
        RECT -27.870 2565.490 -26.690 2566.670 ;
        RECT -27.870 2387.090 -26.690 2388.270 ;
        RECT -27.870 2385.490 -26.690 2386.670 ;
        RECT -27.870 2207.090 -26.690 2208.270 ;
        RECT -27.870 2205.490 -26.690 2206.670 ;
        RECT -27.870 2027.090 -26.690 2028.270 ;
        RECT -27.870 2025.490 -26.690 2026.670 ;
        RECT -27.870 1847.090 -26.690 1848.270 ;
        RECT -27.870 1845.490 -26.690 1846.670 ;
        RECT -27.870 1667.090 -26.690 1668.270 ;
        RECT -27.870 1665.490 -26.690 1666.670 ;
        RECT -27.870 1487.090 -26.690 1488.270 ;
        RECT -27.870 1485.490 -26.690 1486.670 ;
        RECT -27.870 1307.090 -26.690 1308.270 ;
        RECT -27.870 1305.490 -26.690 1306.670 ;
        RECT -27.870 1127.090 -26.690 1128.270 ;
        RECT -27.870 1125.490 -26.690 1126.670 ;
        RECT -27.870 947.090 -26.690 948.270 ;
        RECT -27.870 945.490 -26.690 946.670 ;
        RECT -27.870 767.090 -26.690 768.270 ;
        RECT -27.870 765.490 -26.690 766.670 ;
        RECT -27.870 587.090 -26.690 588.270 ;
        RECT -27.870 585.490 -26.690 586.670 ;
        RECT -27.870 407.090 -26.690 408.270 ;
        RECT -27.870 405.490 -26.690 406.670 ;
        RECT -27.870 227.090 -26.690 228.270 ;
        RECT -27.870 225.490 -26.690 226.670 ;
        RECT -27.870 47.090 -26.690 48.270 ;
        RECT -27.870 45.490 -26.690 46.670 ;
        RECT -27.870 -21.710 -26.690 -20.530 ;
        RECT -27.870 -23.310 -26.690 -22.130 ;
        RECT 40.930 3541.810 42.110 3542.990 ;
        RECT 40.930 3540.210 42.110 3541.390 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.710 42.110 -20.530 ;
        RECT 40.930 -23.310 42.110 -22.130 ;
        RECT 220.930 3541.810 222.110 3542.990 ;
        RECT 220.930 3540.210 222.110 3541.390 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.710 222.110 -20.530 ;
        RECT 220.930 -23.310 222.110 -22.130 ;
        RECT 400.930 3541.810 402.110 3542.990 ;
        RECT 400.930 3540.210 402.110 3541.390 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.710 402.110 -20.530 ;
        RECT 400.930 -23.310 402.110 -22.130 ;
        RECT 580.930 3541.810 582.110 3542.990 ;
        RECT 580.930 3540.210 582.110 3541.390 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.710 582.110 -20.530 ;
        RECT 580.930 -23.310 582.110 -22.130 ;
        RECT 760.930 3541.810 762.110 3542.990 ;
        RECT 760.930 3540.210 762.110 3541.390 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.710 762.110 -20.530 ;
        RECT 760.930 -23.310 762.110 -22.130 ;
        RECT 940.930 3541.810 942.110 3542.990 ;
        RECT 940.930 3540.210 942.110 3541.390 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.710 942.110 -20.530 ;
        RECT 940.930 -23.310 942.110 -22.130 ;
        RECT 1120.930 3541.810 1122.110 3542.990 ;
        RECT 1120.930 3540.210 1122.110 3541.390 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.710 1122.110 -20.530 ;
        RECT 1120.930 -23.310 1122.110 -22.130 ;
        RECT 1300.930 3541.810 1302.110 3542.990 ;
        RECT 1300.930 3540.210 1302.110 3541.390 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.710 1302.110 -20.530 ;
        RECT 1300.930 -23.310 1302.110 -22.130 ;
        RECT 1480.930 3541.810 1482.110 3542.990 ;
        RECT 1480.930 3540.210 1482.110 3541.390 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.710 1482.110 -20.530 ;
        RECT 1480.930 -23.310 1482.110 -22.130 ;
        RECT 1660.930 3541.810 1662.110 3542.990 ;
        RECT 1660.930 3540.210 1662.110 3541.390 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.710 1662.110 -20.530 ;
        RECT 1660.930 -23.310 1662.110 -22.130 ;
        RECT 1840.930 3541.810 1842.110 3542.990 ;
        RECT 1840.930 3540.210 1842.110 3541.390 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.710 1842.110 -20.530 ;
        RECT 1840.930 -23.310 1842.110 -22.130 ;
        RECT 2020.930 3541.810 2022.110 3542.990 ;
        RECT 2020.930 3540.210 2022.110 3541.390 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.710 2022.110 -20.530 ;
        RECT 2020.930 -23.310 2022.110 -22.130 ;
        RECT 2200.930 3541.810 2202.110 3542.990 ;
        RECT 2200.930 3540.210 2202.110 3541.390 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.710 2202.110 -20.530 ;
        RECT 2200.930 -23.310 2202.110 -22.130 ;
        RECT 2380.930 3541.810 2382.110 3542.990 ;
        RECT 2380.930 3540.210 2382.110 3541.390 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.710 2382.110 -20.530 ;
        RECT 2380.930 -23.310 2382.110 -22.130 ;
        RECT 2560.930 3541.810 2562.110 3542.990 ;
        RECT 2560.930 3540.210 2562.110 3541.390 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.710 2562.110 -20.530 ;
        RECT 2560.930 -23.310 2562.110 -22.130 ;
        RECT 2740.930 3541.810 2742.110 3542.990 ;
        RECT 2740.930 3540.210 2742.110 3541.390 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.710 2742.110 -20.530 ;
        RECT 2740.930 -23.310 2742.110 -22.130 ;
        RECT 2946.310 3541.810 2947.490 3542.990 ;
        RECT 2946.310 3540.210 2947.490 3541.390 ;
        RECT 2946.310 3467.090 2947.490 3468.270 ;
        RECT 2946.310 3465.490 2947.490 3466.670 ;
        RECT 2946.310 3287.090 2947.490 3288.270 ;
        RECT 2946.310 3285.490 2947.490 3286.670 ;
        RECT 2946.310 3107.090 2947.490 3108.270 ;
        RECT 2946.310 3105.490 2947.490 3106.670 ;
        RECT 2946.310 2927.090 2947.490 2928.270 ;
        RECT 2946.310 2925.490 2947.490 2926.670 ;
        RECT 2946.310 2747.090 2947.490 2748.270 ;
        RECT 2946.310 2745.490 2947.490 2746.670 ;
        RECT 2946.310 2567.090 2947.490 2568.270 ;
        RECT 2946.310 2565.490 2947.490 2566.670 ;
        RECT 2946.310 2387.090 2947.490 2388.270 ;
        RECT 2946.310 2385.490 2947.490 2386.670 ;
        RECT 2946.310 2207.090 2947.490 2208.270 ;
        RECT 2946.310 2205.490 2947.490 2206.670 ;
        RECT 2946.310 2027.090 2947.490 2028.270 ;
        RECT 2946.310 2025.490 2947.490 2026.670 ;
        RECT 2946.310 1847.090 2947.490 1848.270 ;
        RECT 2946.310 1845.490 2947.490 1846.670 ;
        RECT 2946.310 1667.090 2947.490 1668.270 ;
        RECT 2946.310 1665.490 2947.490 1666.670 ;
        RECT 2946.310 1487.090 2947.490 1488.270 ;
        RECT 2946.310 1485.490 2947.490 1486.670 ;
        RECT 2946.310 1307.090 2947.490 1308.270 ;
        RECT 2946.310 1305.490 2947.490 1306.670 ;
        RECT 2946.310 1127.090 2947.490 1128.270 ;
        RECT 2946.310 1125.490 2947.490 1126.670 ;
        RECT 2946.310 947.090 2947.490 948.270 ;
        RECT 2946.310 945.490 2947.490 946.670 ;
        RECT 2946.310 767.090 2947.490 768.270 ;
        RECT 2946.310 765.490 2947.490 766.670 ;
        RECT 2946.310 587.090 2947.490 588.270 ;
        RECT 2946.310 585.490 2947.490 586.670 ;
        RECT 2946.310 407.090 2947.490 408.270 ;
        RECT 2946.310 405.490 2947.490 406.670 ;
        RECT 2946.310 227.090 2947.490 228.270 ;
        RECT 2946.310 225.490 2947.490 226.670 ;
        RECT 2946.310 47.090 2947.490 48.270 ;
        RECT 2946.310 45.490 2947.490 46.670 ;
        RECT 2946.310 -21.710 2947.490 -20.530 ;
        RECT 2946.310 -23.310 2947.490 -22.130 ;
      LAYER met5 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 40.020 3543.100 43.020 3543.110 ;
        RECT 220.020 3543.100 223.020 3543.110 ;
        RECT 400.020 3543.100 403.020 3543.110 ;
        RECT 580.020 3543.100 583.020 3543.110 ;
        RECT 760.020 3543.100 763.020 3543.110 ;
        RECT 940.020 3543.100 943.020 3543.110 ;
        RECT 1120.020 3543.100 1123.020 3543.110 ;
        RECT 1300.020 3543.100 1303.020 3543.110 ;
        RECT 1480.020 3543.100 1483.020 3543.110 ;
        RECT 1660.020 3543.100 1663.020 3543.110 ;
        RECT 1840.020 3543.100 1843.020 3543.110 ;
        RECT 2020.020 3543.100 2023.020 3543.110 ;
        RECT 2200.020 3543.100 2203.020 3543.110 ;
        RECT 2380.020 3543.100 2383.020 3543.110 ;
        RECT 2560.020 3543.100 2563.020 3543.110 ;
        RECT 2740.020 3543.100 2743.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 40.020 3540.090 43.020 3540.100 ;
        RECT 220.020 3540.090 223.020 3540.100 ;
        RECT 400.020 3540.090 403.020 3540.100 ;
        RECT 580.020 3540.090 583.020 3540.100 ;
        RECT 760.020 3540.090 763.020 3540.100 ;
        RECT 940.020 3540.090 943.020 3540.100 ;
        RECT 1120.020 3540.090 1123.020 3540.100 ;
        RECT 1300.020 3540.090 1303.020 3540.100 ;
        RECT 1480.020 3540.090 1483.020 3540.100 ;
        RECT 1660.020 3540.090 1663.020 3540.100 ;
        RECT 1840.020 3540.090 1843.020 3540.100 ;
        RECT 2020.020 3540.090 2023.020 3540.100 ;
        RECT 2200.020 3540.090 2203.020 3540.100 ;
        RECT 2380.020 3540.090 2383.020 3540.100 ;
        RECT 2560.020 3540.090 2563.020 3540.100 ;
        RECT 2740.020 3540.090 2743.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -28.780 3468.380 -25.780 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.400 3468.380 2948.400 3468.390 ;
        RECT -33.480 3465.380 2953.100 3468.380 ;
        RECT -28.780 3465.370 -25.780 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.400 3465.370 2948.400 3465.380 ;
        RECT -28.780 3288.380 -25.780 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.400 3288.380 2948.400 3288.390 ;
        RECT -33.480 3285.380 2953.100 3288.380 ;
        RECT -28.780 3285.370 -25.780 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.400 3285.370 2948.400 3285.380 ;
        RECT -28.780 3108.380 -25.780 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.400 3108.380 2948.400 3108.390 ;
        RECT -33.480 3105.380 2953.100 3108.380 ;
        RECT -28.780 3105.370 -25.780 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.400 3105.370 2948.400 3105.380 ;
        RECT -28.780 2928.380 -25.780 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.400 2928.380 2948.400 2928.390 ;
        RECT -33.480 2925.380 2953.100 2928.380 ;
        RECT -28.780 2925.370 -25.780 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.400 2925.370 2948.400 2925.380 ;
        RECT -28.780 2748.380 -25.780 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.400 2748.380 2948.400 2748.390 ;
        RECT -33.480 2745.380 2953.100 2748.380 ;
        RECT -28.780 2745.370 -25.780 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.400 2745.370 2948.400 2745.380 ;
        RECT -28.780 2568.380 -25.780 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.400 2568.380 2948.400 2568.390 ;
        RECT -33.480 2565.380 2953.100 2568.380 ;
        RECT -28.780 2565.370 -25.780 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.400 2565.370 2948.400 2565.380 ;
        RECT -28.780 2388.380 -25.780 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.400 2388.380 2948.400 2388.390 ;
        RECT -33.480 2385.380 2953.100 2388.380 ;
        RECT -28.780 2385.370 -25.780 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.400 2385.370 2948.400 2385.380 ;
        RECT -28.780 2208.380 -25.780 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.400 2208.380 2948.400 2208.390 ;
        RECT -33.480 2205.380 2953.100 2208.380 ;
        RECT -28.780 2205.370 -25.780 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.400 2205.370 2948.400 2205.380 ;
        RECT -28.780 2028.380 -25.780 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.400 2028.380 2948.400 2028.390 ;
        RECT -33.480 2025.380 2953.100 2028.380 ;
        RECT -28.780 2025.370 -25.780 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.400 2025.370 2948.400 2025.380 ;
        RECT -28.780 1848.380 -25.780 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.400 1848.380 2948.400 1848.390 ;
        RECT -33.480 1845.380 2953.100 1848.380 ;
        RECT -28.780 1845.370 -25.780 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.400 1845.370 2948.400 1845.380 ;
        RECT -28.780 1668.380 -25.780 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.400 1668.380 2948.400 1668.390 ;
        RECT -33.480 1665.380 2953.100 1668.380 ;
        RECT -28.780 1665.370 -25.780 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.400 1665.370 2948.400 1665.380 ;
        RECT -28.780 1488.380 -25.780 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.400 1488.380 2948.400 1488.390 ;
        RECT -33.480 1485.380 2953.100 1488.380 ;
        RECT -28.780 1485.370 -25.780 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.400 1485.370 2948.400 1485.380 ;
        RECT -28.780 1308.380 -25.780 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.400 1308.380 2948.400 1308.390 ;
        RECT -33.480 1305.380 2953.100 1308.380 ;
        RECT -28.780 1305.370 -25.780 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.400 1305.370 2948.400 1305.380 ;
        RECT -28.780 1128.380 -25.780 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.400 1128.380 2948.400 1128.390 ;
        RECT -33.480 1125.380 2953.100 1128.380 ;
        RECT -28.780 1125.370 -25.780 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.400 1125.370 2948.400 1125.380 ;
        RECT -28.780 948.380 -25.780 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.400 948.380 2948.400 948.390 ;
        RECT -33.480 945.380 2953.100 948.380 ;
        RECT -28.780 945.370 -25.780 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.400 945.370 2948.400 945.380 ;
        RECT -28.780 768.380 -25.780 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.400 768.380 2948.400 768.390 ;
        RECT -33.480 765.380 2953.100 768.380 ;
        RECT -28.780 765.370 -25.780 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.400 765.370 2948.400 765.380 ;
        RECT -28.780 588.380 -25.780 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.400 588.380 2948.400 588.390 ;
        RECT -33.480 585.380 2953.100 588.380 ;
        RECT -28.780 585.370 -25.780 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.400 585.370 2948.400 585.380 ;
        RECT -28.780 408.380 -25.780 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.400 408.380 2948.400 408.390 ;
        RECT -33.480 405.380 2953.100 408.380 ;
        RECT -28.780 405.370 -25.780 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.400 405.370 2948.400 405.380 ;
        RECT -28.780 228.380 -25.780 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.400 228.380 2948.400 228.390 ;
        RECT -33.480 225.380 2953.100 228.380 ;
        RECT -28.780 225.370 -25.780 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.400 225.370 2948.400 225.380 ;
        RECT -28.780 48.380 -25.780 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.400 48.380 2948.400 48.390 ;
        RECT -33.480 45.380 2953.100 48.380 ;
        RECT -28.780 45.370 -25.780 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.400 45.370 2948.400 45.380 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 40.020 -20.420 43.020 -20.410 ;
        RECT 220.020 -20.420 223.020 -20.410 ;
        RECT 400.020 -20.420 403.020 -20.410 ;
        RECT 580.020 -20.420 583.020 -20.410 ;
        RECT 760.020 -20.420 763.020 -20.410 ;
        RECT 940.020 -20.420 943.020 -20.410 ;
        RECT 1120.020 -20.420 1123.020 -20.410 ;
        RECT 1300.020 -20.420 1303.020 -20.410 ;
        RECT 1480.020 -20.420 1483.020 -20.410 ;
        RECT 1660.020 -20.420 1663.020 -20.410 ;
        RECT 1840.020 -20.420 1843.020 -20.410 ;
        RECT 2020.020 -20.420 2023.020 -20.410 ;
        RECT 2200.020 -20.420 2203.020 -20.410 ;
        RECT 2380.020 -20.420 2383.020 -20.410 ;
        RECT 2560.020 -20.420 2563.020 -20.410 ;
        RECT 2740.020 -20.420 2743.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 40.020 -23.430 43.020 -23.420 ;
        RECT 220.020 -23.430 223.020 -23.420 ;
        RECT 400.020 -23.430 403.020 -23.420 ;
        RECT 580.020 -23.430 583.020 -23.420 ;
        RECT 760.020 -23.430 763.020 -23.420 ;
        RECT 940.020 -23.430 943.020 -23.420 ;
        RECT 1120.020 -23.430 1123.020 -23.420 ;
        RECT 1300.020 -23.430 1303.020 -23.420 ;
        RECT 1480.020 -23.430 1483.020 -23.420 ;
        RECT 1660.020 -23.430 1663.020 -23.420 ;
        RECT 1840.020 -23.430 1843.020 -23.420 ;
        RECT 2020.020 -23.430 2023.020 -23.420 ;
        RECT 2200.020 -23.430 2203.020 -23.420 ;
        RECT 2380.020 -23.430 2383.020 -23.420 ;
        RECT 2560.020 -23.430 2563.020 -23.420 ;
        RECT 2740.020 -23.430 2743.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
        RECT 130.020 -28.120 133.020 3547.800 ;
        RECT 310.020 -28.120 313.020 3547.800 ;
        RECT 490.020 -28.120 493.020 3547.800 ;
        RECT 670.020 -28.120 673.020 3547.800 ;
        RECT 850.020 -28.120 853.020 3547.800 ;
        RECT 1030.020 -28.120 1033.020 3547.800 ;
        RECT 1210.020 -28.120 1213.020 3547.800 ;
        RECT 1390.020 -28.120 1393.020 3547.800 ;
        RECT 1570.020 -28.120 1573.020 3547.800 ;
        RECT 1750.020 -28.120 1753.020 3547.800 ;
        RECT 1930.020 -28.120 1933.020 3547.800 ;
        RECT 2110.020 -28.120 2113.020 3547.800 ;
        RECT 2290.020 -28.120 2293.020 3547.800 ;
        RECT 2470.020 -28.120 2473.020 3547.800 ;
        RECT 2650.020 -28.120 2653.020 3547.800 ;
        RECT 2830.020 -28.120 2833.020 3547.800 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
      LAYER via4 ;
        RECT -32.570 3546.510 -31.390 3547.690 ;
        RECT -32.570 3544.910 -31.390 3546.090 ;
        RECT -32.570 3377.090 -31.390 3378.270 ;
        RECT -32.570 3375.490 -31.390 3376.670 ;
        RECT -32.570 3197.090 -31.390 3198.270 ;
        RECT -32.570 3195.490 -31.390 3196.670 ;
        RECT -32.570 3017.090 -31.390 3018.270 ;
        RECT -32.570 3015.490 -31.390 3016.670 ;
        RECT -32.570 2837.090 -31.390 2838.270 ;
        RECT -32.570 2835.490 -31.390 2836.670 ;
        RECT -32.570 2657.090 -31.390 2658.270 ;
        RECT -32.570 2655.490 -31.390 2656.670 ;
        RECT -32.570 2477.090 -31.390 2478.270 ;
        RECT -32.570 2475.490 -31.390 2476.670 ;
        RECT -32.570 2297.090 -31.390 2298.270 ;
        RECT -32.570 2295.490 -31.390 2296.670 ;
        RECT -32.570 2117.090 -31.390 2118.270 ;
        RECT -32.570 2115.490 -31.390 2116.670 ;
        RECT -32.570 1937.090 -31.390 1938.270 ;
        RECT -32.570 1935.490 -31.390 1936.670 ;
        RECT -32.570 1757.090 -31.390 1758.270 ;
        RECT -32.570 1755.490 -31.390 1756.670 ;
        RECT -32.570 1577.090 -31.390 1578.270 ;
        RECT -32.570 1575.490 -31.390 1576.670 ;
        RECT -32.570 1397.090 -31.390 1398.270 ;
        RECT -32.570 1395.490 -31.390 1396.670 ;
        RECT -32.570 1217.090 -31.390 1218.270 ;
        RECT -32.570 1215.490 -31.390 1216.670 ;
        RECT -32.570 1037.090 -31.390 1038.270 ;
        RECT -32.570 1035.490 -31.390 1036.670 ;
        RECT -32.570 857.090 -31.390 858.270 ;
        RECT -32.570 855.490 -31.390 856.670 ;
        RECT -32.570 677.090 -31.390 678.270 ;
        RECT -32.570 675.490 -31.390 676.670 ;
        RECT -32.570 497.090 -31.390 498.270 ;
        RECT -32.570 495.490 -31.390 496.670 ;
        RECT -32.570 317.090 -31.390 318.270 ;
        RECT -32.570 315.490 -31.390 316.670 ;
        RECT -32.570 137.090 -31.390 138.270 ;
        RECT -32.570 135.490 -31.390 136.670 ;
        RECT -32.570 -26.410 -31.390 -25.230 ;
        RECT -32.570 -28.010 -31.390 -26.830 ;
        RECT 130.930 3546.510 132.110 3547.690 ;
        RECT 130.930 3544.910 132.110 3546.090 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -26.410 132.110 -25.230 ;
        RECT 130.930 -28.010 132.110 -26.830 ;
        RECT 310.930 3546.510 312.110 3547.690 ;
        RECT 310.930 3544.910 312.110 3546.090 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -26.410 312.110 -25.230 ;
        RECT 310.930 -28.010 312.110 -26.830 ;
        RECT 490.930 3546.510 492.110 3547.690 ;
        RECT 490.930 3544.910 492.110 3546.090 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -26.410 492.110 -25.230 ;
        RECT 490.930 -28.010 492.110 -26.830 ;
        RECT 670.930 3546.510 672.110 3547.690 ;
        RECT 670.930 3544.910 672.110 3546.090 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -26.410 672.110 -25.230 ;
        RECT 670.930 -28.010 672.110 -26.830 ;
        RECT 850.930 3546.510 852.110 3547.690 ;
        RECT 850.930 3544.910 852.110 3546.090 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -26.410 852.110 -25.230 ;
        RECT 850.930 -28.010 852.110 -26.830 ;
        RECT 1030.930 3546.510 1032.110 3547.690 ;
        RECT 1030.930 3544.910 1032.110 3546.090 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -26.410 1032.110 -25.230 ;
        RECT 1030.930 -28.010 1032.110 -26.830 ;
        RECT 1210.930 3546.510 1212.110 3547.690 ;
        RECT 1210.930 3544.910 1212.110 3546.090 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -26.410 1212.110 -25.230 ;
        RECT 1210.930 -28.010 1212.110 -26.830 ;
        RECT 1390.930 3546.510 1392.110 3547.690 ;
        RECT 1390.930 3544.910 1392.110 3546.090 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -26.410 1392.110 -25.230 ;
        RECT 1390.930 -28.010 1392.110 -26.830 ;
        RECT 1570.930 3546.510 1572.110 3547.690 ;
        RECT 1570.930 3544.910 1572.110 3546.090 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -26.410 1572.110 -25.230 ;
        RECT 1570.930 -28.010 1572.110 -26.830 ;
        RECT 1750.930 3546.510 1752.110 3547.690 ;
        RECT 1750.930 3544.910 1752.110 3546.090 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -26.410 1752.110 -25.230 ;
        RECT 1750.930 -28.010 1752.110 -26.830 ;
        RECT 1930.930 3546.510 1932.110 3547.690 ;
        RECT 1930.930 3544.910 1932.110 3546.090 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -26.410 1932.110 -25.230 ;
        RECT 1930.930 -28.010 1932.110 -26.830 ;
        RECT 2110.930 3546.510 2112.110 3547.690 ;
        RECT 2110.930 3544.910 2112.110 3546.090 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -26.410 2112.110 -25.230 ;
        RECT 2110.930 -28.010 2112.110 -26.830 ;
        RECT 2290.930 3546.510 2292.110 3547.690 ;
        RECT 2290.930 3544.910 2292.110 3546.090 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -26.410 2292.110 -25.230 ;
        RECT 2290.930 -28.010 2292.110 -26.830 ;
        RECT 2470.930 3546.510 2472.110 3547.690 ;
        RECT 2470.930 3544.910 2472.110 3546.090 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -26.410 2472.110 -25.230 ;
        RECT 2470.930 -28.010 2472.110 -26.830 ;
        RECT 2650.930 3546.510 2652.110 3547.690 ;
        RECT 2650.930 3544.910 2652.110 3546.090 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -26.410 2652.110 -25.230 ;
        RECT 2650.930 -28.010 2652.110 -26.830 ;
        RECT 2830.930 3546.510 2832.110 3547.690 ;
        RECT 2830.930 3544.910 2832.110 3546.090 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -26.410 2832.110 -25.230 ;
        RECT 2830.930 -28.010 2832.110 -26.830 ;
        RECT 2951.010 3546.510 2952.190 3547.690 ;
        RECT 2951.010 3544.910 2952.190 3546.090 ;
        RECT 2951.010 3377.090 2952.190 3378.270 ;
        RECT 2951.010 3375.490 2952.190 3376.670 ;
        RECT 2951.010 3197.090 2952.190 3198.270 ;
        RECT 2951.010 3195.490 2952.190 3196.670 ;
        RECT 2951.010 3017.090 2952.190 3018.270 ;
        RECT 2951.010 3015.490 2952.190 3016.670 ;
        RECT 2951.010 2837.090 2952.190 2838.270 ;
        RECT 2951.010 2835.490 2952.190 2836.670 ;
        RECT 2951.010 2657.090 2952.190 2658.270 ;
        RECT 2951.010 2655.490 2952.190 2656.670 ;
        RECT 2951.010 2477.090 2952.190 2478.270 ;
        RECT 2951.010 2475.490 2952.190 2476.670 ;
        RECT 2951.010 2297.090 2952.190 2298.270 ;
        RECT 2951.010 2295.490 2952.190 2296.670 ;
        RECT 2951.010 2117.090 2952.190 2118.270 ;
        RECT 2951.010 2115.490 2952.190 2116.670 ;
        RECT 2951.010 1937.090 2952.190 1938.270 ;
        RECT 2951.010 1935.490 2952.190 1936.670 ;
        RECT 2951.010 1757.090 2952.190 1758.270 ;
        RECT 2951.010 1755.490 2952.190 1756.670 ;
        RECT 2951.010 1577.090 2952.190 1578.270 ;
        RECT 2951.010 1575.490 2952.190 1576.670 ;
        RECT 2951.010 1397.090 2952.190 1398.270 ;
        RECT 2951.010 1395.490 2952.190 1396.670 ;
        RECT 2951.010 1217.090 2952.190 1218.270 ;
        RECT 2951.010 1215.490 2952.190 1216.670 ;
        RECT 2951.010 1037.090 2952.190 1038.270 ;
        RECT 2951.010 1035.490 2952.190 1036.670 ;
        RECT 2951.010 857.090 2952.190 858.270 ;
        RECT 2951.010 855.490 2952.190 856.670 ;
        RECT 2951.010 677.090 2952.190 678.270 ;
        RECT 2951.010 675.490 2952.190 676.670 ;
        RECT 2951.010 497.090 2952.190 498.270 ;
        RECT 2951.010 495.490 2952.190 496.670 ;
        RECT 2951.010 317.090 2952.190 318.270 ;
        RECT 2951.010 315.490 2952.190 316.670 ;
        RECT 2951.010 137.090 2952.190 138.270 ;
        RECT 2951.010 135.490 2952.190 136.670 ;
        RECT 2951.010 -26.410 2952.190 -25.230 ;
        RECT 2951.010 -28.010 2952.190 -26.830 ;
      LAYER met5 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 130.020 3547.800 133.020 3547.810 ;
        RECT 310.020 3547.800 313.020 3547.810 ;
        RECT 490.020 3547.800 493.020 3547.810 ;
        RECT 670.020 3547.800 673.020 3547.810 ;
        RECT 850.020 3547.800 853.020 3547.810 ;
        RECT 1030.020 3547.800 1033.020 3547.810 ;
        RECT 1210.020 3547.800 1213.020 3547.810 ;
        RECT 1390.020 3547.800 1393.020 3547.810 ;
        RECT 1570.020 3547.800 1573.020 3547.810 ;
        RECT 1750.020 3547.800 1753.020 3547.810 ;
        RECT 1930.020 3547.800 1933.020 3547.810 ;
        RECT 2110.020 3547.800 2113.020 3547.810 ;
        RECT 2290.020 3547.800 2293.020 3547.810 ;
        RECT 2470.020 3547.800 2473.020 3547.810 ;
        RECT 2650.020 3547.800 2653.020 3547.810 ;
        RECT 2830.020 3547.800 2833.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 130.020 3544.790 133.020 3544.800 ;
        RECT 310.020 3544.790 313.020 3544.800 ;
        RECT 490.020 3544.790 493.020 3544.800 ;
        RECT 670.020 3544.790 673.020 3544.800 ;
        RECT 850.020 3544.790 853.020 3544.800 ;
        RECT 1030.020 3544.790 1033.020 3544.800 ;
        RECT 1210.020 3544.790 1213.020 3544.800 ;
        RECT 1390.020 3544.790 1393.020 3544.800 ;
        RECT 1570.020 3544.790 1573.020 3544.800 ;
        RECT 1750.020 3544.790 1753.020 3544.800 ;
        RECT 1930.020 3544.790 1933.020 3544.800 ;
        RECT 2110.020 3544.790 2113.020 3544.800 ;
        RECT 2290.020 3544.790 2293.020 3544.800 ;
        RECT 2470.020 3544.790 2473.020 3544.800 ;
        RECT 2650.020 3544.790 2653.020 3544.800 ;
        RECT 2830.020 3544.790 2833.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -33.480 3378.380 -30.480 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2950.100 3378.380 2953.100 3378.390 ;
        RECT -33.480 3375.380 2953.100 3378.380 ;
        RECT -33.480 3375.370 -30.480 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2950.100 3375.370 2953.100 3375.380 ;
        RECT -33.480 3198.380 -30.480 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2950.100 3198.380 2953.100 3198.390 ;
        RECT -33.480 3195.380 2953.100 3198.380 ;
        RECT -33.480 3195.370 -30.480 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2950.100 3195.370 2953.100 3195.380 ;
        RECT -33.480 3018.380 -30.480 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2950.100 3018.380 2953.100 3018.390 ;
        RECT -33.480 3015.380 2953.100 3018.380 ;
        RECT -33.480 3015.370 -30.480 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2950.100 3015.370 2953.100 3015.380 ;
        RECT -33.480 2838.380 -30.480 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2950.100 2838.380 2953.100 2838.390 ;
        RECT -33.480 2835.380 2953.100 2838.380 ;
        RECT -33.480 2835.370 -30.480 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2950.100 2835.370 2953.100 2835.380 ;
        RECT -33.480 2658.380 -30.480 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2950.100 2658.380 2953.100 2658.390 ;
        RECT -33.480 2655.380 2953.100 2658.380 ;
        RECT -33.480 2655.370 -30.480 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2950.100 2655.370 2953.100 2655.380 ;
        RECT -33.480 2478.380 -30.480 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2950.100 2478.380 2953.100 2478.390 ;
        RECT -33.480 2475.380 2953.100 2478.380 ;
        RECT -33.480 2475.370 -30.480 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2950.100 2475.370 2953.100 2475.380 ;
        RECT -33.480 2298.380 -30.480 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2950.100 2298.380 2953.100 2298.390 ;
        RECT -33.480 2295.380 2953.100 2298.380 ;
        RECT -33.480 2295.370 -30.480 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2950.100 2295.370 2953.100 2295.380 ;
        RECT -33.480 2118.380 -30.480 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2950.100 2118.380 2953.100 2118.390 ;
        RECT -33.480 2115.380 2953.100 2118.380 ;
        RECT -33.480 2115.370 -30.480 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2950.100 2115.370 2953.100 2115.380 ;
        RECT -33.480 1938.380 -30.480 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2950.100 1938.380 2953.100 1938.390 ;
        RECT -33.480 1935.380 2953.100 1938.380 ;
        RECT -33.480 1935.370 -30.480 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2950.100 1935.370 2953.100 1935.380 ;
        RECT -33.480 1758.380 -30.480 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2950.100 1758.380 2953.100 1758.390 ;
        RECT -33.480 1755.380 2953.100 1758.380 ;
        RECT -33.480 1755.370 -30.480 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2950.100 1755.370 2953.100 1755.380 ;
        RECT -33.480 1578.380 -30.480 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2950.100 1578.380 2953.100 1578.390 ;
        RECT -33.480 1575.380 2953.100 1578.380 ;
        RECT -33.480 1575.370 -30.480 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2950.100 1575.370 2953.100 1575.380 ;
        RECT -33.480 1398.380 -30.480 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2950.100 1398.380 2953.100 1398.390 ;
        RECT -33.480 1395.380 2953.100 1398.380 ;
        RECT -33.480 1395.370 -30.480 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2950.100 1395.370 2953.100 1395.380 ;
        RECT -33.480 1218.380 -30.480 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2950.100 1218.380 2953.100 1218.390 ;
        RECT -33.480 1215.380 2953.100 1218.380 ;
        RECT -33.480 1215.370 -30.480 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2950.100 1215.370 2953.100 1215.380 ;
        RECT -33.480 1038.380 -30.480 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2950.100 1038.380 2953.100 1038.390 ;
        RECT -33.480 1035.380 2953.100 1038.380 ;
        RECT -33.480 1035.370 -30.480 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2950.100 1035.370 2953.100 1035.380 ;
        RECT -33.480 858.380 -30.480 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2950.100 858.380 2953.100 858.390 ;
        RECT -33.480 855.380 2953.100 858.380 ;
        RECT -33.480 855.370 -30.480 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2950.100 855.370 2953.100 855.380 ;
        RECT -33.480 678.380 -30.480 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2950.100 678.380 2953.100 678.390 ;
        RECT -33.480 675.380 2953.100 678.380 ;
        RECT -33.480 675.370 -30.480 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2950.100 675.370 2953.100 675.380 ;
        RECT -33.480 498.380 -30.480 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2950.100 498.380 2953.100 498.390 ;
        RECT -33.480 495.380 2953.100 498.380 ;
        RECT -33.480 495.370 -30.480 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2950.100 495.370 2953.100 495.380 ;
        RECT -33.480 318.380 -30.480 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2950.100 318.380 2953.100 318.390 ;
        RECT -33.480 315.380 2953.100 318.380 ;
        RECT -33.480 315.370 -30.480 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2950.100 315.370 2953.100 315.380 ;
        RECT -33.480 138.380 -30.480 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2950.100 138.380 2953.100 138.390 ;
        RECT -33.480 135.380 2953.100 138.380 ;
        RECT -33.480 135.370 -30.480 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2950.100 135.370 2953.100 135.380 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 130.020 -25.120 133.020 -25.110 ;
        RECT 310.020 -25.120 313.020 -25.110 ;
        RECT 490.020 -25.120 493.020 -25.110 ;
        RECT 670.020 -25.120 673.020 -25.110 ;
        RECT 850.020 -25.120 853.020 -25.110 ;
        RECT 1030.020 -25.120 1033.020 -25.110 ;
        RECT 1210.020 -25.120 1213.020 -25.110 ;
        RECT 1390.020 -25.120 1393.020 -25.110 ;
        RECT 1570.020 -25.120 1573.020 -25.110 ;
        RECT 1750.020 -25.120 1753.020 -25.110 ;
        RECT 1930.020 -25.120 1933.020 -25.110 ;
        RECT 2110.020 -25.120 2113.020 -25.110 ;
        RECT 2290.020 -25.120 2293.020 -25.110 ;
        RECT 2470.020 -25.120 2473.020 -25.110 ;
        RECT 2650.020 -25.120 2653.020 -25.110 ;
        RECT 2830.020 -25.120 2833.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 130.020 -28.130 133.020 -28.120 ;
        RECT 310.020 -28.130 313.020 -28.120 ;
        RECT 490.020 -28.130 493.020 -28.120 ;
        RECT 670.020 -28.130 673.020 -28.120 ;
        RECT 850.020 -28.130 853.020 -28.120 ;
        RECT 1030.020 -28.130 1033.020 -28.120 ;
        RECT 1210.020 -28.130 1213.020 -28.120 ;
        RECT 1390.020 -28.130 1393.020 -28.120 ;
        RECT 1570.020 -28.130 1573.020 -28.120 ;
        RECT 1750.020 -28.130 1753.020 -28.120 ;
        RECT 1930.020 -28.130 1933.020 -28.120 ;
        RECT 2110.020 -28.130 2113.020 -28.120 ;
        RECT 2290.020 -28.130 2293.020 -28.120 ;
        RECT 2470.020 -28.130 2473.020 -28.120 ;
        RECT 2650.020 -28.130 2653.020 -28.120 ;
        RECT 2830.020 -28.130 2833.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
        RECT 58.020 -37.520 61.020 3557.200 ;
        RECT 238.020 -37.520 241.020 3557.200 ;
        RECT 418.020 -37.520 421.020 3557.200 ;
        RECT 598.020 -37.520 601.020 3557.200 ;
        RECT 778.020 -37.520 781.020 3557.200 ;
        RECT 958.020 -37.520 961.020 3557.200 ;
        RECT 1138.020 -37.520 1141.020 3557.200 ;
        RECT 1318.020 -37.520 1321.020 3557.200 ;
        RECT 1498.020 -37.520 1501.020 3557.200 ;
        RECT 1678.020 -37.520 1681.020 3557.200 ;
        RECT 1858.020 -37.520 1861.020 3557.200 ;
        RECT 2038.020 -37.520 2041.020 3557.200 ;
        RECT 2218.020 -37.520 2221.020 3557.200 ;
        RECT 2398.020 -37.520 2401.020 3557.200 ;
        RECT 2578.020 -37.520 2581.020 3557.200 ;
        RECT 2758.020 -37.520 2761.020 3557.200 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
      LAYER via4 ;
        RECT -37.270 3551.210 -36.090 3552.390 ;
        RECT -37.270 3549.610 -36.090 3550.790 ;
        RECT -37.270 3485.090 -36.090 3486.270 ;
        RECT -37.270 3483.490 -36.090 3484.670 ;
        RECT -37.270 3305.090 -36.090 3306.270 ;
        RECT -37.270 3303.490 -36.090 3304.670 ;
        RECT -37.270 3125.090 -36.090 3126.270 ;
        RECT -37.270 3123.490 -36.090 3124.670 ;
        RECT -37.270 2945.090 -36.090 2946.270 ;
        RECT -37.270 2943.490 -36.090 2944.670 ;
        RECT -37.270 2765.090 -36.090 2766.270 ;
        RECT -37.270 2763.490 -36.090 2764.670 ;
        RECT -37.270 2585.090 -36.090 2586.270 ;
        RECT -37.270 2583.490 -36.090 2584.670 ;
        RECT -37.270 2405.090 -36.090 2406.270 ;
        RECT -37.270 2403.490 -36.090 2404.670 ;
        RECT -37.270 2225.090 -36.090 2226.270 ;
        RECT -37.270 2223.490 -36.090 2224.670 ;
        RECT -37.270 2045.090 -36.090 2046.270 ;
        RECT -37.270 2043.490 -36.090 2044.670 ;
        RECT -37.270 1865.090 -36.090 1866.270 ;
        RECT -37.270 1863.490 -36.090 1864.670 ;
        RECT -37.270 1685.090 -36.090 1686.270 ;
        RECT -37.270 1683.490 -36.090 1684.670 ;
        RECT -37.270 1505.090 -36.090 1506.270 ;
        RECT -37.270 1503.490 -36.090 1504.670 ;
        RECT -37.270 1325.090 -36.090 1326.270 ;
        RECT -37.270 1323.490 -36.090 1324.670 ;
        RECT -37.270 1145.090 -36.090 1146.270 ;
        RECT -37.270 1143.490 -36.090 1144.670 ;
        RECT -37.270 965.090 -36.090 966.270 ;
        RECT -37.270 963.490 -36.090 964.670 ;
        RECT -37.270 785.090 -36.090 786.270 ;
        RECT -37.270 783.490 -36.090 784.670 ;
        RECT -37.270 605.090 -36.090 606.270 ;
        RECT -37.270 603.490 -36.090 604.670 ;
        RECT -37.270 425.090 -36.090 426.270 ;
        RECT -37.270 423.490 -36.090 424.670 ;
        RECT -37.270 245.090 -36.090 246.270 ;
        RECT -37.270 243.490 -36.090 244.670 ;
        RECT -37.270 65.090 -36.090 66.270 ;
        RECT -37.270 63.490 -36.090 64.670 ;
        RECT -37.270 -31.110 -36.090 -29.930 ;
        RECT -37.270 -32.710 -36.090 -31.530 ;
        RECT 58.930 3551.210 60.110 3552.390 ;
        RECT 58.930 3549.610 60.110 3550.790 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -31.110 60.110 -29.930 ;
        RECT 58.930 -32.710 60.110 -31.530 ;
        RECT 238.930 3551.210 240.110 3552.390 ;
        RECT 238.930 3549.610 240.110 3550.790 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -31.110 240.110 -29.930 ;
        RECT 238.930 -32.710 240.110 -31.530 ;
        RECT 418.930 3551.210 420.110 3552.390 ;
        RECT 418.930 3549.610 420.110 3550.790 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -31.110 420.110 -29.930 ;
        RECT 418.930 -32.710 420.110 -31.530 ;
        RECT 598.930 3551.210 600.110 3552.390 ;
        RECT 598.930 3549.610 600.110 3550.790 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -31.110 600.110 -29.930 ;
        RECT 598.930 -32.710 600.110 -31.530 ;
        RECT 778.930 3551.210 780.110 3552.390 ;
        RECT 778.930 3549.610 780.110 3550.790 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -31.110 780.110 -29.930 ;
        RECT 778.930 -32.710 780.110 -31.530 ;
        RECT 958.930 3551.210 960.110 3552.390 ;
        RECT 958.930 3549.610 960.110 3550.790 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -31.110 960.110 -29.930 ;
        RECT 958.930 -32.710 960.110 -31.530 ;
        RECT 1138.930 3551.210 1140.110 3552.390 ;
        RECT 1138.930 3549.610 1140.110 3550.790 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -31.110 1140.110 -29.930 ;
        RECT 1138.930 -32.710 1140.110 -31.530 ;
        RECT 1318.930 3551.210 1320.110 3552.390 ;
        RECT 1318.930 3549.610 1320.110 3550.790 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -31.110 1320.110 -29.930 ;
        RECT 1318.930 -32.710 1320.110 -31.530 ;
        RECT 1498.930 3551.210 1500.110 3552.390 ;
        RECT 1498.930 3549.610 1500.110 3550.790 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -31.110 1500.110 -29.930 ;
        RECT 1498.930 -32.710 1500.110 -31.530 ;
        RECT 1678.930 3551.210 1680.110 3552.390 ;
        RECT 1678.930 3549.610 1680.110 3550.790 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -31.110 1680.110 -29.930 ;
        RECT 1678.930 -32.710 1680.110 -31.530 ;
        RECT 1858.930 3551.210 1860.110 3552.390 ;
        RECT 1858.930 3549.610 1860.110 3550.790 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -31.110 1860.110 -29.930 ;
        RECT 1858.930 -32.710 1860.110 -31.530 ;
        RECT 2038.930 3551.210 2040.110 3552.390 ;
        RECT 2038.930 3549.610 2040.110 3550.790 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -31.110 2040.110 -29.930 ;
        RECT 2038.930 -32.710 2040.110 -31.530 ;
        RECT 2218.930 3551.210 2220.110 3552.390 ;
        RECT 2218.930 3549.610 2220.110 3550.790 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -31.110 2220.110 -29.930 ;
        RECT 2218.930 -32.710 2220.110 -31.530 ;
        RECT 2398.930 3551.210 2400.110 3552.390 ;
        RECT 2398.930 3549.610 2400.110 3550.790 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -31.110 2400.110 -29.930 ;
        RECT 2398.930 -32.710 2400.110 -31.530 ;
        RECT 2578.930 3551.210 2580.110 3552.390 ;
        RECT 2578.930 3549.610 2580.110 3550.790 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -31.110 2580.110 -29.930 ;
        RECT 2578.930 -32.710 2580.110 -31.530 ;
        RECT 2758.930 3551.210 2760.110 3552.390 ;
        RECT 2758.930 3549.610 2760.110 3550.790 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -31.110 2760.110 -29.930 ;
        RECT 2758.930 -32.710 2760.110 -31.530 ;
        RECT 2955.710 3551.210 2956.890 3552.390 ;
        RECT 2955.710 3549.610 2956.890 3550.790 ;
        RECT 2955.710 3485.090 2956.890 3486.270 ;
        RECT 2955.710 3483.490 2956.890 3484.670 ;
        RECT 2955.710 3305.090 2956.890 3306.270 ;
        RECT 2955.710 3303.490 2956.890 3304.670 ;
        RECT 2955.710 3125.090 2956.890 3126.270 ;
        RECT 2955.710 3123.490 2956.890 3124.670 ;
        RECT 2955.710 2945.090 2956.890 2946.270 ;
        RECT 2955.710 2943.490 2956.890 2944.670 ;
        RECT 2955.710 2765.090 2956.890 2766.270 ;
        RECT 2955.710 2763.490 2956.890 2764.670 ;
        RECT 2955.710 2585.090 2956.890 2586.270 ;
        RECT 2955.710 2583.490 2956.890 2584.670 ;
        RECT 2955.710 2405.090 2956.890 2406.270 ;
        RECT 2955.710 2403.490 2956.890 2404.670 ;
        RECT 2955.710 2225.090 2956.890 2226.270 ;
        RECT 2955.710 2223.490 2956.890 2224.670 ;
        RECT 2955.710 2045.090 2956.890 2046.270 ;
        RECT 2955.710 2043.490 2956.890 2044.670 ;
        RECT 2955.710 1865.090 2956.890 1866.270 ;
        RECT 2955.710 1863.490 2956.890 1864.670 ;
        RECT 2955.710 1685.090 2956.890 1686.270 ;
        RECT 2955.710 1683.490 2956.890 1684.670 ;
        RECT 2955.710 1505.090 2956.890 1506.270 ;
        RECT 2955.710 1503.490 2956.890 1504.670 ;
        RECT 2955.710 1325.090 2956.890 1326.270 ;
        RECT 2955.710 1323.490 2956.890 1324.670 ;
        RECT 2955.710 1145.090 2956.890 1146.270 ;
        RECT 2955.710 1143.490 2956.890 1144.670 ;
        RECT 2955.710 965.090 2956.890 966.270 ;
        RECT 2955.710 963.490 2956.890 964.670 ;
        RECT 2955.710 785.090 2956.890 786.270 ;
        RECT 2955.710 783.490 2956.890 784.670 ;
        RECT 2955.710 605.090 2956.890 606.270 ;
        RECT 2955.710 603.490 2956.890 604.670 ;
        RECT 2955.710 425.090 2956.890 426.270 ;
        RECT 2955.710 423.490 2956.890 424.670 ;
        RECT 2955.710 245.090 2956.890 246.270 ;
        RECT 2955.710 243.490 2956.890 244.670 ;
        RECT 2955.710 65.090 2956.890 66.270 ;
        RECT 2955.710 63.490 2956.890 64.670 ;
        RECT 2955.710 -31.110 2956.890 -29.930 ;
        RECT 2955.710 -32.710 2956.890 -31.530 ;
      LAYER met5 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 58.020 3552.500 61.020 3552.510 ;
        RECT 238.020 3552.500 241.020 3552.510 ;
        RECT 418.020 3552.500 421.020 3552.510 ;
        RECT 598.020 3552.500 601.020 3552.510 ;
        RECT 778.020 3552.500 781.020 3552.510 ;
        RECT 958.020 3552.500 961.020 3552.510 ;
        RECT 1138.020 3552.500 1141.020 3552.510 ;
        RECT 1318.020 3552.500 1321.020 3552.510 ;
        RECT 1498.020 3552.500 1501.020 3552.510 ;
        RECT 1678.020 3552.500 1681.020 3552.510 ;
        RECT 1858.020 3552.500 1861.020 3552.510 ;
        RECT 2038.020 3552.500 2041.020 3552.510 ;
        RECT 2218.020 3552.500 2221.020 3552.510 ;
        RECT 2398.020 3552.500 2401.020 3552.510 ;
        RECT 2578.020 3552.500 2581.020 3552.510 ;
        RECT 2758.020 3552.500 2761.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 58.020 3549.490 61.020 3549.500 ;
        RECT 238.020 3549.490 241.020 3549.500 ;
        RECT 418.020 3549.490 421.020 3549.500 ;
        RECT 598.020 3549.490 601.020 3549.500 ;
        RECT 778.020 3549.490 781.020 3549.500 ;
        RECT 958.020 3549.490 961.020 3549.500 ;
        RECT 1138.020 3549.490 1141.020 3549.500 ;
        RECT 1318.020 3549.490 1321.020 3549.500 ;
        RECT 1498.020 3549.490 1501.020 3549.500 ;
        RECT 1678.020 3549.490 1681.020 3549.500 ;
        RECT 1858.020 3549.490 1861.020 3549.500 ;
        RECT 2038.020 3549.490 2041.020 3549.500 ;
        RECT 2218.020 3549.490 2221.020 3549.500 ;
        RECT 2398.020 3549.490 2401.020 3549.500 ;
        RECT 2578.020 3549.490 2581.020 3549.500 ;
        RECT 2758.020 3549.490 2761.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -38.180 3486.380 -35.180 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.800 3486.380 2957.800 3486.390 ;
        RECT -42.880 3483.380 2962.500 3486.380 ;
        RECT -38.180 3483.370 -35.180 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.800 3483.370 2957.800 3483.380 ;
        RECT -38.180 3306.380 -35.180 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.800 3306.380 2957.800 3306.390 ;
        RECT -42.880 3303.380 2962.500 3306.380 ;
        RECT -38.180 3303.370 -35.180 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.800 3303.370 2957.800 3303.380 ;
        RECT -38.180 3126.380 -35.180 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.800 3126.380 2957.800 3126.390 ;
        RECT -42.880 3123.380 2962.500 3126.380 ;
        RECT -38.180 3123.370 -35.180 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.800 3123.370 2957.800 3123.380 ;
        RECT -38.180 2946.380 -35.180 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.800 2946.380 2957.800 2946.390 ;
        RECT -42.880 2943.380 2962.500 2946.380 ;
        RECT -38.180 2943.370 -35.180 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.800 2943.370 2957.800 2943.380 ;
        RECT -38.180 2766.380 -35.180 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.800 2766.380 2957.800 2766.390 ;
        RECT -42.880 2763.380 2962.500 2766.380 ;
        RECT -38.180 2763.370 -35.180 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.800 2763.370 2957.800 2763.380 ;
        RECT -38.180 2586.380 -35.180 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.800 2586.380 2957.800 2586.390 ;
        RECT -42.880 2583.380 2962.500 2586.380 ;
        RECT -38.180 2583.370 -35.180 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.800 2583.370 2957.800 2583.380 ;
        RECT -38.180 2406.380 -35.180 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.800 2406.380 2957.800 2406.390 ;
        RECT -42.880 2403.380 2962.500 2406.380 ;
        RECT -38.180 2403.370 -35.180 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.800 2403.370 2957.800 2403.380 ;
        RECT -38.180 2226.380 -35.180 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.800 2226.380 2957.800 2226.390 ;
        RECT -42.880 2223.380 2962.500 2226.380 ;
        RECT -38.180 2223.370 -35.180 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.800 2223.370 2957.800 2223.380 ;
        RECT -38.180 2046.380 -35.180 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.800 2046.380 2957.800 2046.390 ;
        RECT -42.880 2043.380 2962.500 2046.380 ;
        RECT -38.180 2043.370 -35.180 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.800 2043.370 2957.800 2043.380 ;
        RECT -38.180 1866.380 -35.180 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.800 1866.380 2957.800 1866.390 ;
        RECT -42.880 1863.380 2962.500 1866.380 ;
        RECT -38.180 1863.370 -35.180 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.800 1863.370 2957.800 1863.380 ;
        RECT -38.180 1686.380 -35.180 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.800 1686.380 2957.800 1686.390 ;
        RECT -42.880 1683.380 2962.500 1686.380 ;
        RECT -38.180 1683.370 -35.180 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.800 1683.370 2957.800 1683.380 ;
        RECT -38.180 1506.380 -35.180 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.800 1506.380 2957.800 1506.390 ;
        RECT -42.880 1503.380 2962.500 1506.380 ;
        RECT -38.180 1503.370 -35.180 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.800 1503.370 2957.800 1503.380 ;
        RECT -38.180 1326.380 -35.180 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.800 1326.380 2957.800 1326.390 ;
        RECT -42.880 1323.380 2962.500 1326.380 ;
        RECT -38.180 1323.370 -35.180 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.800 1323.370 2957.800 1323.380 ;
        RECT -38.180 1146.380 -35.180 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.800 1146.380 2957.800 1146.390 ;
        RECT -42.880 1143.380 2962.500 1146.380 ;
        RECT -38.180 1143.370 -35.180 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.800 1143.370 2957.800 1143.380 ;
        RECT -38.180 966.380 -35.180 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.800 966.380 2957.800 966.390 ;
        RECT -42.880 963.380 2962.500 966.380 ;
        RECT -38.180 963.370 -35.180 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.800 963.370 2957.800 963.380 ;
        RECT -38.180 786.380 -35.180 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.800 786.380 2957.800 786.390 ;
        RECT -42.880 783.380 2962.500 786.380 ;
        RECT -38.180 783.370 -35.180 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.800 783.370 2957.800 783.380 ;
        RECT -38.180 606.380 -35.180 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.800 606.380 2957.800 606.390 ;
        RECT -42.880 603.380 2962.500 606.380 ;
        RECT -38.180 603.370 -35.180 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.800 603.370 2957.800 603.380 ;
        RECT -38.180 426.380 -35.180 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.800 426.380 2957.800 426.390 ;
        RECT -42.880 423.380 2962.500 426.380 ;
        RECT -38.180 423.370 -35.180 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.800 423.370 2957.800 423.380 ;
        RECT -38.180 246.380 -35.180 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.800 246.380 2957.800 246.390 ;
        RECT -42.880 243.380 2962.500 246.380 ;
        RECT -38.180 243.370 -35.180 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.800 243.370 2957.800 243.380 ;
        RECT -38.180 66.380 -35.180 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.800 66.380 2957.800 66.390 ;
        RECT -42.880 63.380 2962.500 66.380 ;
        RECT -38.180 63.370 -35.180 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.800 63.370 2957.800 63.380 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 58.020 -29.820 61.020 -29.810 ;
        RECT 238.020 -29.820 241.020 -29.810 ;
        RECT 418.020 -29.820 421.020 -29.810 ;
        RECT 598.020 -29.820 601.020 -29.810 ;
        RECT 778.020 -29.820 781.020 -29.810 ;
        RECT 958.020 -29.820 961.020 -29.810 ;
        RECT 1138.020 -29.820 1141.020 -29.810 ;
        RECT 1318.020 -29.820 1321.020 -29.810 ;
        RECT 1498.020 -29.820 1501.020 -29.810 ;
        RECT 1678.020 -29.820 1681.020 -29.810 ;
        RECT 1858.020 -29.820 1861.020 -29.810 ;
        RECT 2038.020 -29.820 2041.020 -29.810 ;
        RECT 2218.020 -29.820 2221.020 -29.810 ;
        RECT 2398.020 -29.820 2401.020 -29.810 ;
        RECT 2578.020 -29.820 2581.020 -29.810 ;
        RECT 2758.020 -29.820 2761.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 58.020 -32.830 61.020 -32.820 ;
        RECT 238.020 -32.830 241.020 -32.820 ;
        RECT 418.020 -32.830 421.020 -32.820 ;
        RECT 598.020 -32.830 601.020 -32.820 ;
        RECT 778.020 -32.830 781.020 -32.820 ;
        RECT 958.020 -32.830 961.020 -32.820 ;
        RECT 1138.020 -32.830 1141.020 -32.820 ;
        RECT 1318.020 -32.830 1321.020 -32.820 ;
        RECT 1498.020 -32.830 1501.020 -32.820 ;
        RECT 1678.020 -32.830 1681.020 -32.820 ;
        RECT 1858.020 -32.830 1861.020 -32.820 ;
        RECT 2038.020 -32.830 2041.020 -32.820 ;
        RECT 2218.020 -32.830 2221.020 -32.820 ;
        RECT 2398.020 -32.830 2401.020 -32.820 ;
        RECT 2578.020 -32.830 2581.020 -32.820 ;
        RECT 2758.020 -32.830 2761.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
        RECT 148.020 -37.520 151.020 3557.200 ;
        RECT 328.020 -37.520 331.020 3557.200 ;
        RECT 508.020 -37.520 511.020 3557.200 ;
        RECT 688.020 -37.520 691.020 3557.200 ;
        RECT 868.020 -37.520 871.020 3557.200 ;
        RECT 1048.020 -37.520 1051.020 3557.200 ;
        RECT 1228.020 -37.520 1231.020 3557.200 ;
        RECT 1408.020 -37.520 1411.020 3557.200 ;
        RECT 1588.020 -37.520 1591.020 3557.200 ;
        RECT 1768.020 -37.520 1771.020 3557.200 ;
        RECT 1948.020 -37.520 1951.020 3557.200 ;
        RECT 2128.020 -37.520 2131.020 3557.200 ;
        RECT 2308.020 -37.520 2311.020 3557.200 ;
        RECT 2488.020 -37.520 2491.020 3557.200 ;
        RECT 2668.020 -37.520 2671.020 3557.200 ;
        RECT 2848.020 -37.520 2851.020 3557.200 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
      LAYER via4 ;
        RECT -41.970 3555.910 -40.790 3557.090 ;
        RECT -41.970 3554.310 -40.790 3555.490 ;
        RECT -41.970 3395.090 -40.790 3396.270 ;
        RECT -41.970 3393.490 -40.790 3394.670 ;
        RECT -41.970 3215.090 -40.790 3216.270 ;
        RECT -41.970 3213.490 -40.790 3214.670 ;
        RECT -41.970 3035.090 -40.790 3036.270 ;
        RECT -41.970 3033.490 -40.790 3034.670 ;
        RECT -41.970 2855.090 -40.790 2856.270 ;
        RECT -41.970 2853.490 -40.790 2854.670 ;
        RECT -41.970 2675.090 -40.790 2676.270 ;
        RECT -41.970 2673.490 -40.790 2674.670 ;
        RECT -41.970 2495.090 -40.790 2496.270 ;
        RECT -41.970 2493.490 -40.790 2494.670 ;
        RECT -41.970 2315.090 -40.790 2316.270 ;
        RECT -41.970 2313.490 -40.790 2314.670 ;
        RECT -41.970 2135.090 -40.790 2136.270 ;
        RECT -41.970 2133.490 -40.790 2134.670 ;
        RECT -41.970 1955.090 -40.790 1956.270 ;
        RECT -41.970 1953.490 -40.790 1954.670 ;
        RECT -41.970 1775.090 -40.790 1776.270 ;
        RECT -41.970 1773.490 -40.790 1774.670 ;
        RECT -41.970 1595.090 -40.790 1596.270 ;
        RECT -41.970 1593.490 -40.790 1594.670 ;
        RECT -41.970 1415.090 -40.790 1416.270 ;
        RECT -41.970 1413.490 -40.790 1414.670 ;
        RECT -41.970 1235.090 -40.790 1236.270 ;
        RECT -41.970 1233.490 -40.790 1234.670 ;
        RECT -41.970 1055.090 -40.790 1056.270 ;
        RECT -41.970 1053.490 -40.790 1054.670 ;
        RECT -41.970 875.090 -40.790 876.270 ;
        RECT -41.970 873.490 -40.790 874.670 ;
        RECT -41.970 695.090 -40.790 696.270 ;
        RECT -41.970 693.490 -40.790 694.670 ;
        RECT -41.970 515.090 -40.790 516.270 ;
        RECT -41.970 513.490 -40.790 514.670 ;
        RECT -41.970 335.090 -40.790 336.270 ;
        RECT -41.970 333.490 -40.790 334.670 ;
        RECT -41.970 155.090 -40.790 156.270 ;
        RECT -41.970 153.490 -40.790 154.670 ;
        RECT -41.970 -35.810 -40.790 -34.630 ;
        RECT -41.970 -37.410 -40.790 -36.230 ;
        RECT 148.930 3555.910 150.110 3557.090 ;
        RECT 148.930 3554.310 150.110 3555.490 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.810 150.110 -34.630 ;
        RECT 148.930 -37.410 150.110 -36.230 ;
        RECT 328.930 3555.910 330.110 3557.090 ;
        RECT 328.930 3554.310 330.110 3555.490 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.810 330.110 -34.630 ;
        RECT 328.930 -37.410 330.110 -36.230 ;
        RECT 508.930 3555.910 510.110 3557.090 ;
        RECT 508.930 3554.310 510.110 3555.490 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.810 510.110 -34.630 ;
        RECT 508.930 -37.410 510.110 -36.230 ;
        RECT 688.930 3555.910 690.110 3557.090 ;
        RECT 688.930 3554.310 690.110 3555.490 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.810 690.110 -34.630 ;
        RECT 688.930 -37.410 690.110 -36.230 ;
        RECT 868.930 3555.910 870.110 3557.090 ;
        RECT 868.930 3554.310 870.110 3555.490 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.810 870.110 -34.630 ;
        RECT 868.930 -37.410 870.110 -36.230 ;
        RECT 1048.930 3555.910 1050.110 3557.090 ;
        RECT 1048.930 3554.310 1050.110 3555.490 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.810 1050.110 -34.630 ;
        RECT 1048.930 -37.410 1050.110 -36.230 ;
        RECT 1228.930 3555.910 1230.110 3557.090 ;
        RECT 1228.930 3554.310 1230.110 3555.490 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.810 1230.110 -34.630 ;
        RECT 1228.930 -37.410 1230.110 -36.230 ;
        RECT 1408.930 3555.910 1410.110 3557.090 ;
        RECT 1408.930 3554.310 1410.110 3555.490 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.810 1410.110 -34.630 ;
        RECT 1408.930 -37.410 1410.110 -36.230 ;
        RECT 1588.930 3555.910 1590.110 3557.090 ;
        RECT 1588.930 3554.310 1590.110 3555.490 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.810 1590.110 -34.630 ;
        RECT 1588.930 -37.410 1590.110 -36.230 ;
        RECT 1768.930 3555.910 1770.110 3557.090 ;
        RECT 1768.930 3554.310 1770.110 3555.490 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.810 1770.110 -34.630 ;
        RECT 1768.930 -37.410 1770.110 -36.230 ;
        RECT 1948.930 3555.910 1950.110 3557.090 ;
        RECT 1948.930 3554.310 1950.110 3555.490 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.810 1950.110 -34.630 ;
        RECT 1948.930 -37.410 1950.110 -36.230 ;
        RECT 2128.930 3555.910 2130.110 3557.090 ;
        RECT 2128.930 3554.310 2130.110 3555.490 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.810 2130.110 -34.630 ;
        RECT 2128.930 -37.410 2130.110 -36.230 ;
        RECT 2308.930 3555.910 2310.110 3557.090 ;
        RECT 2308.930 3554.310 2310.110 3555.490 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.810 2310.110 -34.630 ;
        RECT 2308.930 -37.410 2310.110 -36.230 ;
        RECT 2488.930 3555.910 2490.110 3557.090 ;
        RECT 2488.930 3554.310 2490.110 3555.490 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.810 2490.110 -34.630 ;
        RECT 2488.930 -37.410 2490.110 -36.230 ;
        RECT 2668.930 3555.910 2670.110 3557.090 ;
        RECT 2668.930 3554.310 2670.110 3555.490 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.810 2670.110 -34.630 ;
        RECT 2668.930 -37.410 2670.110 -36.230 ;
        RECT 2848.930 3555.910 2850.110 3557.090 ;
        RECT 2848.930 3554.310 2850.110 3555.490 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.810 2850.110 -34.630 ;
        RECT 2848.930 -37.410 2850.110 -36.230 ;
        RECT 2960.410 3555.910 2961.590 3557.090 ;
        RECT 2960.410 3554.310 2961.590 3555.490 ;
        RECT 2960.410 3395.090 2961.590 3396.270 ;
        RECT 2960.410 3393.490 2961.590 3394.670 ;
        RECT 2960.410 3215.090 2961.590 3216.270 ;
        RECT 2960.410 3213.490 2961.590 3214.670 ;
        RECT 2960.410 3035.090 2961.590 3036.270 ;
        RECT 2960.410 3033.490 2961.590 3034.670 ;
        RECT 2960.410 2855.090 2961.590 2856.270 ;
        RECT 2960.410 2853.490 2961.590 2854.670 ;
        RECT 2960.410 2675.090 2961.590 2676.270 ;
        RECT 2960.410 2673.490 2961.590 2674.670 ;
        RECT 2960.410 2495.090 2961.590 2496.270 ;
        RECT 2960.410 2493.490 2961.590 2494.670 ;
        RECT 2960.410 2315.090 2961.590 2316.270 ;
        RECT 2960.410 2313.490 2961.590 2314.670 ;
        RECT 2960.410 2135.090 2961.590 2136.270 ;
        RECT 2960.410 2133.490 2961.590 2134.670 ;
        RECT 2960.410 1955.090 2961.590 1956.270 ;
        RECT 2960.410 1953.490 2961.590 1954.670 ;
        RECT 2960.410 1775.090 2961.590 1776.270 ;
        RECT 2960.410 1773.490 2961.590 1774.670 ;
        RECT 2960.410 1595.090 2961.590 1596.270 ;
        RECT 2960.410 1593.490 2961.590 1594.670 ;
        RECT 2960.410 1415.090 2961.590 1416.270 ;
        RECT 2960.410 1413.490 2961.590 1414.670 ;
        RECT 2960.410 1235.090 2961.590 1236.270 ;
        RECT 2960.410 1233.490 2961.590 1234.670 ;
        RECT 2960.410 1055.090 2961.590 1056.270 ;
        RECT 2960.410 1053.490 2961.590 1054.670 ;
        RECT 2960.410 875.090 2961.590 876.270 ;
        RECT 2960.410 873.490 2961.590 874.670 ;
        RECT 2960.410 695.090 2961.590 696.270 ;
        RECT 2960.410 693.490 2961.590 694.670 ;
        RECT 2960.410 515.090 2961.590 516.270 ;
        RECT 2960.410 513.490 2961.590 514.670 ;
        RECT 2960.410 335.090 2961.590 336.270 ;
        RECT 2960.410 333.490 2961.590 334.670 ;
        RECT 2960.410 155.090 2961.590 156.270 ;
        RECT 2960.410 153.490 2961.590 154.670 ;
        RECT 2960.410 -35.810 2961.590 -34.630 ;
        RECT 2960.410 -37.410 2961.590 -36.230 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 148.020 3557.200 151.020 3557.210 ;
        RECT 328.020 3557.200 331.020 3557.210 ;
        RECT 508.020 3557.200 511.020 3557.210 ;
        RECT 688.020 3557.200 691.020 3557.210 ;
        RECT 868.020 3557.200 871.020 3557.210 ;
        RECT 1048.020 3557.200 1051.020 3557.210 ;
        RECT 1228.020 3557.200 1231.020 3557.210 ;
        RECT 1408.020 3557.200 1411.020 3557.210 ;
        RECT 1588.020 3557.200 1591.020 3557.210 ;
        RECT 1768.020 3557.200 1771.020 3557.210 ;
        RECT 1948.020 3557.200 1951.020 3557.210 ;
        RECT 2128.020 3557.200 2131.020 3557.210 ;
        RECT 2308.020 3557.200 2311.020 3557.210 ;
        RECT 2488.020 3557.200 2491.020 3557.210 ;
        RECT 2668.020 3557.200 2671.020 3557.210 ;
        RECT 2848.020 3557.200 2851.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 148.020 3554.190 151.020 3554.200 ;
        RECT 328.020 3554.190 331.020 3554.200 ;
        RECT 508.020 3554.190 511.020 3554.200 ;
        RECT 688.020 3554.190 691.020 3554.200 ;
        RECT 868.020 3554.190 871.020 3554.200 ;
        RECT 1048.020 3554.190 1051.020 3554.200 ;
        RECT 1228.020 3554.190 1231.020 3554.200 ;
        RECT 1408.020 3554.190 1411.020 3554.200 ;
        RECT 1588.020 3554.190 1591.020 3554.200 ;
        RECT 1768.020 3554.190 1771.020 3554.200 ;
        RECT 1948.020 3554.190 1951.020 3554.200 ;
        RECT 2128.020 3554.190 2131.020 3554.200 ;
        RECT 2308.020 3554.190 2311.020 3554.200 ;
        RECT 2488.020 3554.190 2491.020 3554.200 ;
        RECT 2668.020 3554.190 2671.020 3554.200 ;
        RECT 2848.020 3554.190 2851.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -42.880 3396.380 -39.880 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2959.500 3396.380 2962.500 3396.390 ;
        RECT -42.880 3393.380 2962.500 3396.380 ;
        RECT -42.880 3393.370 -39.880 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2959.500 3393.370 2962.500 3393.380 ;
        RECT -42.880 3216.380 -39.880 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2959.500 3216.380 2962.500 3216.390 ;
        RECT -42.880 3213.380 2962.500 3216.380 ;
        RECT -42.880 3213.370 -39.880 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2959.500 3213.370 2962.500 3213.380 ;
        RECT -42.880 3036.380 -39.880 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2959.500 3036.380 2962.500 3036.390 ;
        RECT -42.880 3033.380 2962.500 3036.380 ;
        RECT -42.880 3033.370 -39.880 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2959.500 3033.370 2962.500 3033.380 ;
        RECT -42.880 2856.380 -39.880 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2959.500 2856.380 2962.500 2856.390 ;
        RECT -42.880 2853.380 2962.500 2856.380 ;
        RECT -42.880 2853.370 -39.880 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2959.500 2853.370 2962.500 2853.380 ;
        RECT -42.880 2676.380 -39.880 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2959.500 2676.380 2962.500 2676.390 ;
        RECT -42.880 2673.380 2962.500 2676.380 ;
        RECT -42.880 2673.370 -39.880 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2959.500 2673.370 2962.500 2673.380 ;
        RECT -42.880 2496.380 -39.880 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2959.500 2496.380 2962.500 2496.390 ;
        RECT -42.880 2493.380 2962.500 2496.380 ;
        RECT -42.880 2493.370 -39.880 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2959.500 2493.370 2962.500 2493.380 ;
        RECT -42.880 2316.380 -39.880 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2959.500 2316.380 2962.500 2316.390 ;
        RECT -42.880 2313.380 2962.500 2316.380 ;
        RECT -42.880 2313.370 -39.880 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2959.500 2313.370 2962.500 2313.380 ;
        RECT -42.880 2136.380 -39.880 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2959.500 2136.380 2962.500 2136.390 ;
        RECT -42.880 2133.380 2962.500 2136.380 ;
        RECT -42.880 2133.370 -39.880 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2959.500 2133.370 2962.500 2133.380 ;
        RECT -42.880 1956.380 -39.880 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2959.500 1956.380 2962.500 1956.390 ;
        RECT -42.880 1953.380 2962.500 1956.380 ;
        RECT -42.880 1953.370 -39.880 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2959.500 1953.370 2962.500 1953.380 ;
        RECT -42.880 1776.380 -39.880 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2959.500 1776.380 2962.500 1776.390 ;
        RECT -42.880 1773.380 2962.500 1776.380 ;
        RECT -42.880 1773.370 -39.880 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2959.500 1773.370 2962.500 1773.380 ;
        RECT -42.880 1596.380 -39.880 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2959.500 1596.380 2962.500 1596.390 ;
        RECT -42.880 1593.380 2962.500 1596.380 ;
        RECT -42.880 1593.370 -39.880 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2959.500 1593.370 2962.500 1593.380 ;
        RECT -42.880 1416.380 -39.880 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2959.500 1416.380 2962.500 1416.390 ;
        RECT -42.880 1413.380 2962.500 1416.380 ;
        RECT -42.880 1413.370 -39.880 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2959.500 1413.370 2962.500 1413.380 ;
        RECT -42.880 1236.380 -39.880 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2959.500 1236.380 2962.500 1236.390 ;
        RECT -42.880 1233.380 2962.500 1236.380 ;
        RECT -42.880 1233.370 -39.880 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2959.500 1233.370 2962.500 1233.380 ;
        RECT -42.880 1056.380 -39.880 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2959.500 1056.380 2962.500 1056.390 ;
        RECT -42.880 1053.380 2962.500 1056.380 ;
        RECT -42.880 1053.370 -39.880 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2959.500 1053.370 2962.500 1053.380 ;
        RECT -42.880 876.380 -39.880 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2959.500 876.380 2962.500 876.390 ;
        RECT -42.880 873.380 2962.500 876.380 ;
        RECT -42.880 873.370 -39.880 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2959.500 873.370 2962.500 873.380 ;
        RECT -42.880 696.380 -39.880 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2959.500 696.380 2962.500 696.390 ;
        RECT -42.880 693.380 2962.500 696.380 ;
        RECT -42.880 693.370 -39.880 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2959.500 693.370 2962.500 693.380 ;
        RECT -42.880 516.380 -39.880 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2959.500 516.380 2962.500 516.390 ;
        RECT -42.880 513.380 2962.500 516.380 ;
        RECT -42.880 513.370 -39.880 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2959.500 513.370 2962.500 513.380 ;
        RECT -42.880 336.380 -39.880 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2959.500 336.380 2962.500 336.390 ;
        RECT -42.880 333.380 2962.500 336.380 ;
        RECT -42.880 333.370 -39.880 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2959.500 333.370 2962.500 333.380 ;
        RECT -42.880 156.380 -39.880 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2959.500 156.380 2962.500 156.390 ;
        RECT -42.880 153.380 2962.500 156.380 ;
        RECT -42.880 153.370 -39.880 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2959.500 153.370 2962.500 153.380 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 148.020 -34.520 151.020 -34.510 ;
        RECT 328.020 -34.520 331.020 -34.510 ;
        RECT 508.020 -34.520 511.020 -34.510 ;
        RECT 688.020 -34.520 691.020 -34.510 ;
        RECT 868.020 -34.520 871.020 -34.510 ;
        RECT 1048.020 -34.520 1051.020 -34.510 ;
        RECT 1228.020 -34.520 1231.020 -34.510 ;
        RECT 1408.020 -34.520 1411.020 -34.510 ;
        RECT 1588.020 -34.520 1591.020 -34.510 ;
        RECT 1768.020 -34.520 1771.020 -34.510 ;
        RECT 1948.020 -34.520 1951.020 -34.510 ;
        RECT 2128.020 -34.520 2131.020 -34.510 ;
        RECT 2308.020 -34.520 2311.020 -34.510 ;
        RECT 2488.020 -34.520 2491.020 -34.510 ;
        RECT 2668.020 -34.520 2671.020 -34.510 ;
        RECT 2848.020 -34.520 2851.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 148.020 -37.530 151.020 -37.520 ;
        RECT 328.020 -37.530 331.020 -37.520 ;
        RECT 508.020 -37.530 511.020 -37.520 ;
        RECT 688.020 -37.530 691.020 -37.520 ;
        RECT 868.020 -37.530 871.020 -37.520 ;
        RECT 1048.020 -37.530 1051.020 -37.520 ;
        RECT 1228.020 -37.530 1231.020 -37.520 ;
        RECT 1408.020 -37.530 1411.020 -37.520 ;
        RECT 1588.020 -37.530 1591.020 -37.520 ;
        RECT 1768.020 -37.530 1771.020 -37.520 ;
        RECT 1948.020 -37.530 1951.020 -37.520 ;
        RECT 2128.020 -37.530 2131.020 -37.520 ;
        RECT 2308.020 -37.530 2311.020 -37.520 ;
        RECT 2488.020 -37.530 2491.020 -37.520 ;
        RECT 2668.020 -37.530 2671.020 -37.520 ;
        RECT 2848.020 -37.530 2851.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 1154.535 1710.795 2343.175 2888.725 ;
      LAYER met1 ;
        RECT 1154.535 1705.480 2347.705 2888.880 ;
      LAYER met2 ;
        RECT 1150.025 2895.720 1153.885 2896.000 ;
        RECT 1154.725 2895.720 1164.005 2896.000 ;
        RECT 1164.845 2895.720 1174.585 2896.000 ;
        RECT 1175.425 2895.720 1185.165 2896.000 ;
        RECT 1186.005 2895.720 1195.745 2896.000 ;
        RECT 1196.585 2895.720 1206.325 2896.000 ;
        RECT 1207.165 2895.720 1216.905 2896.000 ;
        RECT 1217.745 2895.720 1227.485 2896.000 ;
        RECT 1228.325 2895.720 1238.065 2896.000 ;
        RECT 1238.905 2895.720 1248.185 2896.000 ;
        RECT 1249.025 2895.720 1258.765 2896.000 ;
        RECT 1259.605 2895.720 1269.345 2896.000 ;
        RECT 1270.185 2895.720 1279.925 2896.000 ;
        RECT 1280.765 2895.720 1290.505 2896.000 ;
        RECT 1291.345 2895.720 1301.085 2896.000 ;
        RECT 1301.925 2895.720 1311.665 2896.000 ;
        RECT 1312.505 2895.720 1322.245 2896.000 ;
        RECT 1323.085 2895.720 1332.825 2896.000 ;
        RECT 1333.665 2895.720 1342.945 2896.000 ;
        RECT 1343.785 2895.720 1353.525 2896.000 ;
        RECT 1354.365 2895.720 1364.105 2896.000 ;
        RECT 1364.945 2895.720 1374.685 2896.000 ;
        RECT 1375.525 2895.720 1385.265 2896.000 ;
        RECT 1386.105 2895.720 1395.845 2896.000 ;
        RECT 1396.685 2895.720 1406.425 2896.000 ;
        RECT 1407.265 2895.720 1417.005 2896.000 ;
        RECT 1417.845 2895.720 1427.585 2896.000 ;
        RECT 1428.425 2895.720 1437.705 2896.000 ;
        RECT 1438.545 2895.720 1448.285 2896.000 ;
        RECT 1449.125 2895.720 1458.865 2896.000 ;
        RECT 1459.705 2895.720 1469.445 2896.000 ;
        RECT 1470.285 2895.720 1480.025 2896.000 ;
        RECT 1480.865 2895.720 1490.605 2896.000 ;
        RECT 1491.445 2895.720 1501.185 2896.000 ;
        RECT 1502.025 2895.720 1511.765 2896.000 ;
        RECT 1512.605 2895.720 1522.345 2896.000 ;
        RECT 1523.185 2895.720 1532.465 2896.000 ;
        RECT 1533.305 2895.720 1543.045 2896.000 ;
        RECT 1543.885 2895.720 1553.625 2896.000 ;
        RECT 1554.465 2895.720 1564.205 2896.000 ;
        RECT 1565.045 2895.720 1574.785 2896.000 ;
        RECT 1575.625 2895.720 1585.365 2896.000 ;
        RECT 1586.205 2895.720 1595.945 2896.000 ;
        RECT 1596.785 2895.720 1606.525 2896.000 ;
        RECT 1607.365 2895.720 1616.645 2896.000 ;
        RECT 1617.485 2895.720 1627.225 2896.000 ;
        RECT 1628.065 2895.720 1637.805 2896.000 ;
        RECT 1638.645 2895.720 1648.385 2896.000 ;
        RECT 1649.225 2895.720 1658.965 2896.000 ;
        RECT 1659.805 2895.720 1669.545 2896.000 ;
        RECT 1670.385 2895.720 1680.125 2896.000 ;
        RECT 1680.965 2895.720 1690.705 2896.000 ;
        RECT 1691.545 2895.720 1701.285 2896.000 ;
        RECT 1702.125 2895.720 1711.405 2896.000 ;
        RECT 1712.245 2895.720 1721.985 2896.000 ;
        RECT 1722.825 2895.720 1732.565 2896.000 ;
        RECT 1733.405 2895.720 1743.145 2896.000 ;
        RECT 1743.985 2895.720 1753.725 2896.000 ;
        RECT 1754.565 2895.720 1764.305 2896.000 ;
        RECT 1765.145 2895.720 1774.885 2896.000 ;
        RECT 1775.725 2895.720 1785.465 2896.000 ;
        RECT 1786.305 2895.720 1796.045 2896.000 ;
        RECT 1796.885 2895.720 1806.165 2896.000 ;
        RECT 1807.005 2895.720 1816.745 2896.000 ;
        RECT 1817.585 2895.720 1827.325 2896.000 ;
        RECT 1828.165 2895.720 1837.905 2896.000 ;
        RECT 1838.745 2895.720 1848.485 2896.000 ;
        RECT 1849.325 2895.720 1859.065 2896.000 ;
        RECT 1859.905 2895.720 1869.645 2896.000 ;
        RECT 1870.485 2895.720 1880.225 2896.000 ;
        RECT 1881.065 2895.720 1890.805 2896.000 ;
        RECT 1891.645 2895.720 1900.925 2896.000 ;
        RECT 1901.765 2895.720 1911.505 2896.000 ;
        RECT 1912.345 2895.720 1922.085 2896.000 ;
        RECT 1922.925 2895.720 1932.665 2896.000 ;
        RECT 1933.505 2895.720 1943.245 2896.000 ;
        RECT 1944.085 2895.720 1953.825 2896.000 ;
        RECT 1954.665 2895.720 1964.405 2896.000 ;
        RECT 1965.245 2895.720 1974.985 2896.000 ;
        RECT 1975.825 2895.720 1985.105 2896.000 ;
        RECT 1985.945 2895.720 1995.685 2896.000 ;
        RECT 1996.525 2895.720 2006.265 2896.000 ;
        RECT 2007.105 2895.720 2016.845 2896.000 ;
        RECT 2017.685 2895.720 2027.425 2896.000 ;
        RECT 2028.265 2895.720 2038.005 2896.000 ;
        RECT 2038.845 2895.720 2048.585 2896.000 ;
        RECT 2049.425 2895.720 2059.165 2896.000 ;
        RECT 2060.005 2895.720 2069.745 2896.000 ;
        RECT 2070.585 2895.720 2079.865 2896.000 ;
        RECT 2080.705 2895.720 2090.445 2896.000 ;
        RECT 2091.285 2895.720 2101.025 2896.000 ;
        RECT 2101.865 2895.720 2111.605 2896.000 ;
        RECT 2112.445 2895.720 2122.185 2896.000 ;
        RECT 2123.025 2895.720 2132.765 2896.000 ;
        RECT 2133.605 2895.720 2143.345 2896.000 ;
        RECT 2144.185 2895.720 2153.925 2896.000 ;
        RECT 2154.765 2895.720 2164.505 2896.000 ;
        RECT 2165.345 2895.720 2174.625 2896.000 ;
        RECT 2175.465 2895.720 2185.205 2896.000 ;
        RECT 2186.045 2895.720 2195.785 2896.000 ;
        RECT 2196.625 2895.720 2206.365 2896.000 ;
        RECT 2207.205 2895.720 2216.945 2896.000 ;
        RECT 2217.785 2895.720 2227.525 2896.000 ;
        RECT 2228.365 2895.720 2238.105 2896.000 ;
        RECT 2238.945 2895.720 2248.685 2896.000 ;
        RECT 2249.525 2895.720 2259.265 2896.000 ;
        RECT 2260.105 2895.720 2269.385 2896.000 ;
        RECT 2270.225 2895.720 2279.965 2896.000 ;
        RECT 2280.805 2895.720 2290.545 2896.000 ;
        RECT 2291.385 2895.720 2301.125 2896.000 ;
        RECT 2301.965 2895.720 2311.705 2896.000 ;
        RECT 2312.545 2895.720 2322.285 2896.000 ;
        RECT 2323.125 2895.720 2332.865 2896.000 ;
        RECT 2333.705 2895.720 2343.445 2896.000 ;
        RECT 2344.285 2895.720 2347.675 2896.000 ;
        RECT 1150.025 1704.280 2347.675 2895.720 ;
        RECT 1150.585 1704.000 1152.045 1704.280 ;
        RECT 1152.885 1704.000 1154.345 1704.280 ;
        RECT 1155.185 1704.000 1156.645 1704.280 ;
        RECT 1157.485 1704.000 1159.405 1704.280 ;
        RECT 1160.245 1704.000 1161.705 1704.280 ;
        RECT 1162.545 1704.000 1164.005 1704.280 ;
        RECT 1164.845 1704.000 1166.765 1704.280 ;
        RECT 1167.605 1704.000 1169.065 1704.280 ;
        RECT 1169.905 1704.000 1171.365 1704.280 ;
        RECT 1172.205 1704.000 1174.125 1704.280 ;
        RECT 1174.965 1704.000 1176.425 1704.280 ;
        RECT 1177.265 1704.000 1178.725 1704.280 ;
        RECT 1179.565 1704.000 1181.485 1704.280 ;
        RECT 1182.325 1704.000 1183.785 1704.280 ;
        RECT 1184.625 1704.000 1186.085 1704.280 ;
        RECT 1186.925 1704.000 1188.845 1704.280 ;
        RECT 1189.685 1704.000 1191.145 1704.280 ;
        RECT 1191.985 1704.000 1193.445 1704.280 ;
        RECT 1194.285 1704.000 1196.205 1704.280 ;
        RECT 1197.045 1704.000 1198.505 1704.280 ;
        RECT 1199.345 1704.000 1200.805 1704.280 ;
        RECT 1201.645 1704.000 1203.565 1704.280 ;
        RECT 1204.405 1704.000 1205.865 1704.280 ;
        RECT 1206.705 1704.000 1208.165 1704.280 ;
        RECT 1209.005 1704.000 1210.925 1704.280 ;
        RECT 1211.765 1704.000 1213.225 1704.280 ;
        RECT 1214.065 1704.000 1215.525 1704.280 ;
        RECT 1216.365 1704.000 1218.285 1704.280 ;
        RECT 1219.125 1704.000 1220.585 1704.280 ;
        RECT 1221.425 1704.000 1222.885 1704.280 ;
        RECT 1223.725 1704.000 1225.645 1704.280 ;
        RECT 1226.485 1704.000 1227.945 1704.280 ;
        RECT 1228.785 1704.000 1230.245 1704.280 ;
        RECT 1231.085 1704.000 1233.005 1704.280 ;
        RECT 1233.845 1704.000 1235.305 1704.280 ;
        RECT 1236.145 1704.000 1237.605 1704.280 ;
        RECT 1238.445 1704.000 1240.365 1704.280 ;
        RECT 1241.205 1704.000 1242.665 1704.280 ;
        RECT 1243.505 1704.000 1244.965 1704.280 ;
        RECT 1245.805 1704.000 1247.265 1704.280 ;
        RECT 1248.105 1704.000 1250.025 1704.280 ;
        RECT 1250.865 1704.000 1252.325 1704.280 ;
        RECT 1253.165 1704.000 1254.625 1704.280 ;
        RECT 1255.465 1704.000 1257.385 1704.280 ;
        RECT 1258.225 1704.000 1259.685 1704.280 ;
        RECT 1260.525 1704.000 1261.985 1704.280 ;
        RECT 1262.825 1704.000 1264.745 1704.280 ;
        RECT 1265.585 1704.000 1267.045 1704.280 ;
        RECT 1267.885 1704.000 1269.345 1704.280 ;
        RECT 1270.185 1704.000 1272.105 1704.280 ;
        RECT 1272.945 1704.000 1274.405 1704.280 ;
        RECT 1275.245 1704.000 1276.705 1704.280 ;
        RECT 1277.545 1704.000 1279.465 1704.280 ;
        RECT 1280.305 1704.000 1281.765 1704.280 ;
        RECT 1282.605 1704.000 1284.065 1704.280 ;
        RECT 1284.905 1704.000 1286.825 1704.280 ;
        RECT 1287.665 1704.000 1289.125 1704.280 ;
        RECT 1289.965 1704.000 1291.425 1704.280 ;
        RECT 1292.265 1704.000 1294.185 1704.280 ;
        RECT 1295.025 1704.000 1296.485 1704.280 ;
        RECT 1297.325 1704.000 1298.785 1704.280 ;
        RECT 1299.625 1704.000 1301.545 1704.280 ;
        RECT 1302.385 1704.000 1303.845 1704.280 ;
        RECT 1304.685 1704.000 1306.145 1704.280 ;
        RECT 1306.985 1704.000 1308.905 1704.280 ;
        RECT 1309.745 1704.000 1311.205 1704.280 ;
        RECT 1312.045 1704.000 1313.505 1704.280 ;
        RECT 1314.345 1704.000 1316.265 1704.280 ;
        RECT 1317.105 1704.000 1318.565 1704.280 ;
        RECT 1319.405 1704.000 1320.865 1704.280 ;
        RECT 1321.705 1704.000 1323.625 1704.280 ;
        RECT 1324.465 1704.000 1325.925 1704.280 ;
        RECT 1326.765 1704.000 1328.225 1704.280 ;
        RECT 1329.065 1704.000 1330.985 1704.280 ;
        RECT 1331.825 1704.000 1333.285 1704.280 ;
        RECT 1334.125 1704.000 1335.585 1704.280 ;
        RECT 1336.425 1704.000 1337.885 1704.280 ;
        RECT 1338.725 1704.000 1340.645 1704.280 ;
        RECT 1341.485 1704.000 1342.945 1704.280 ;
        RECT 1343.785 1704.000 1345.245 1704.280 ;
        RECT 1346.085 1704.000 1348.005 1704.280 ;
        RECT 1348.845 1704.000 1350.305 1704.280 ;
        RECT 1351.145 1704.000 1352.605 1704.280 ;
        RECT 1353.445 1704.000 1355.365 1704.280 ;
        RECT 1356.205 1704.000 1357.665 1704.280 ;
        RECT 1358.505 1704.000 1359.965 1704.280 ;
        RECT 1360.805 1704.000 1362.725 1704.280 ;
        RECT 1363.565 1704.000 1365.025 1704.280 ;
        RECT 1365.865 1704.000 1367.325 1704.280 ;
        RECT 1368.165 1704.000 1370.085 1704.280 ;
        RECT 1370.925 1704.000 1372.385 1704.280 ;
        RECT 1373.225 1704.000 1374.685 1704.280 ;
        RECT 1375.525 1704.000 1377.445 1704.280 ;
        RECT 1378.285 1704.000 1379.745 1704.280 ;
        RECT 1380.585 1704.000 1382.045 1704.280 ;
        RECT 1382.885 1704.000 1384.805 1704.280 ;
        RECT 1385.645 1704.000 1387.105 1704.280 ;
        RECT 1387.945 1704.000 1389.405 1704.280 ;
        RECT 1390.245 1704.000 1392.165 1704.280 ;
        RECT 1393.005 1704.000 1394.465 1704.280 ;
        RECT 1395.305 1704.000 1396.765 1704.280 ;
        RECT 1397.605 1704.000 1399.525 1704.280 ;
        RECT 1400.365 1704.000 1401.825 1704.280 ;
        RECT 1402.665 1704.000 1404.125 1704.280 ;
        RECT 1404.965 1704.000 1406.885 1704.280 ;
        RECT 1407.725 1704.000 1409.185 1704.280 ;
        RECT 1410.025 1704.000 1411.485 1704.280 ;
        RECT 1412.325 1704.000 1414.245 1704.280 ;
        RECT 1415.085 1704.000 1416.545 1704.280 ;
        RECT 1417.385 1704.000 1418.845 1704.280 ;
        RECT 1419.685 1704.000 1421.605 1704.280 ;
        RECT 1422.445 1704.000 1423.905 1704.280 ;
        RECT 1424.745 1704.000 1426.205 1704.280 ;
        RECT 1427.045 1704.000 1428.505 1704.280 ;
        RECT 1429.345 1704.000 1431.265 1704.280 ;
        RECT 1432.105 1704.000 1433.565 1704.280 ;
        RECT 1434.405 1704.000 1435.865 1704.280 ;
        RECT 1436.705 1704.000 1438.625 1704.280 ;
        RECT 1439.465 1704.000 1440.925 1704.280 ;
        RECT 1441.765 1704.000 1443.225 1704.280 ;
        RECT 1444.065 1704.000 1445.985 1704.280 ;
        RECT 1446.825 1704.000 1448.285 1704.280 ;
        RECT 1449.125 1704.000 1450.585 1704.280 ;
        RECT 1451.425 1704.000 1453.345 1704.280 ;
        RECT 1454.185 1704.000 1455.645 1704.280 ;
        RECT 1456.485 1704.000 1457.945 1704.280 ;
        RECT 1458.785 1704.000 1460.705 1704.280 ;
        RECT 1461.545 1704.000 1463.005 1704.280 ;
        RECT 1463.845 1704.000 1465.305 1704.280 ;
        RECT 1466.145 1704.000 1468.065 1704.280 ;
        RECT 1468.905 1704.000 1470.365 1704.280 ;
        RECT 1471.205 1704.000 1472.665 1704.280 ;
        RECT 1473.505 1704.000 1475.425 1704.280 ;
        RECT 1476.265 1704.000 1477.725 1704.280 ;
        RECT 1478.565 1704.000 1480.025 1704.280 ;
        RECT 1480.865 1704.000 1482.785 1704.280 ;
        RECT 1483.625 1704.000 1485.085 1704.280 ;
        RECT 1485.925 1704.000 1487.385 1704.280 ;
        RECT 1488.225 1704.000 1490.145 1704.280 ;
        RECT 1490.985 1704.000 1492.445 1704.280 ;
        RECT 1493.285 1704.000 1494.745 1704.280 ;
        RECT 1495.585 1704.000 1497.505 1704.280 ;
        RECT 1498.345 1704.000 1499.805 1704.280 ;
        RECT 1500.645 1704.000 1502.105 1704.280 ;
        RECT 1502.945 1704.000 1504.865 1704.280 ;
        RECT 1505.705 1704.000 1507.165 1704.280 ;
        RECT 1508.005 1704.000 1509.465 1704.280 ;
        RECT 1510.305 1704.000 1512.225 1704.280 ;
        RECT 1513.065 1704.000 1514.525 1704.280 ;
        RECT 1515.365 1704.000 1516.825 1704.280 ;
        RECT 1517.665 1704.000 1519.125 1704.280 ;
        RECT 1519.965 1704.000 1521.885 1704.280 ;
        RECT 1522.725 1704.000 1524.185 1704.280 ;
        RECT 1525.025 1704.000 1526.485 1704.280 ;
        RECT 1527.325 1704.000 1529.245 1704.280 ;
        RECT 1530.085 1704.000 1531.545 1704.280 ;
        RECT 1532.385 1704.000 1533.845 1704.280 ;
        RECT 1534.685 1704.000 1536.605 1704.280 ;
        RECT 1537.445 1704.000 1538.905 1704.280 ;
        RECT 1539.745 1704.000 1541.205 1704.280 ;
        RECT 1542.045 1704.000 1543.965 1704.280 ;
        RECT 1544.805 1704.000 1546.265 1704.280 ;
        RECT 1547.105 1704.000 1548.565 1704.280 ;
        RECT 1549.405 1704.000 1551.325 1704.280 ;
        RECT 1552.165 1704.000 1553.625 1704.280 ;
        RECT 1554.465 1704.000 1555.925 1704.280 ;
        RECT 1556.765 1704.000 1558.685 1704.280 ;
        RECT 1559.525 1704.000 1560.985 1704.280 ;
        RECT 1561.825 1704.000 1563.285 1704.280 ;
        RECT 1564.125 1704.000 1566.045 1704.280 ;
        RECT 1566.885 1704.000 1568.345 1704.280 ;
        RECT 1569.185 1704.000 1570.645 1704.280 ;
        RECT 1571.485 1704.000 1573.405 1704.280 ;
        RECT 1574.245 1704.000 1575.705 1704.280 ;
        RECT 1576.545 1704.000 1578.005 1704.280 ;
        RECT 1578.845 1704.000 1580.765 1704.280 ;
        RECT 1581.605 1704.000 1583.065 1704.280 ;
        RECT 1583.905 1704.000 1585.365 1704.280 ;
        RECT 1586.205 1704.000 1588.125 1704.280 ;
        RECT 1588.965 1704.000 1590.425 1704.280 ;
        RECT 1591.265 1704.000 1592.725 1704.280 ;
        RECT 1593.565 1704.000 1595.485 1704.280 ;
        RECT 1596.325 1704.000 1597.785 1704.280 ;
        RECT 1598.625 1704.000 1600.085 1704.280 ;
        RECT 1600.925 1704.000 1602.845 1704.280 ;
        RECT 1603.685 1704.000 1605.145 1704.280 ;
        RECT 1605.985 1704.000 1607.445 1704.280 ;
        RECT 1608.285 1704.000 1610.205 1704.280 ;
        RECT 1611.045 1704.000 1612.505 1704.280 ;
        RECT 1613.345 1704.000 1614.805 1704.280 ;
        RECT 1615.645 1704.000 1617.105 1704.280 ;
        RECT 1617.945 1704.000 1619.865 1704.280 ;
        RECT 1620.705 1704.000 1622.165 1704.280 ;
        RECT 1623.005 1704.000 1624.465 1704.280 ;
        RECT 1625.305 1704.000 1627.225 1704.280 ;
        RECT 1628.065 1704.000 1629.525 1704.280 ;
        RECT 1630.365 1704.000 1631.825 1704.280 ;
        RECT 1632.665 1704.000 1634.585 1704.280 ;
        RECT 1635.425 1704.000 1636.885 1704.280 ;
        RECT 1637.725 1704.000 1639.185 1704.280 ;
        RECT 1640.025 1704.000 1641.945 1704.280 ;
        RECT 1642.785 1704.000 1644.245 1704.280 ;
        RECT 1645.085 1704.000 1646.545 1704.280 ;
        RECT 1647.385 1704.000 1649.305 1704.280 ;
        RECT 1650.145 1704.000 1651.605 1704.280 ;
        RECT 1652.445 1704.000 1653.905 1704.280 ;
        RECT 1654.745 1704.000 1656.665 1704.280 ;
        RECT 1657.505 1704.000 1658.965 1704.280 ;
        RECT 1659.805 1704.000 1661.265 1704.280 ;
        RECT 1662.105 1704.000 1664.025 1704.280 ;
        RECT 1664.865 1704.000 1666.325 1704.280 ;
        RECT 1667.165 1704.000 1668.625 1704.280 ;
        RECT 1669.465 1704.000 1671.385 1704.280 ;
        RECT 1672.225 1704.000 1673.685 1704.280 ;
        RECT 1674.525 1704.000 1675.985 1704.280 ;
        RECT 1676.825 1704.000 1678.745 1704.280 ;
        RECT 1679.585 1704.000 1681.045 1704.280 ;
        RECT 1681.885 1704.000 1683.345 1704.280 ;
        RECT 1684.185 1704.000 1686.105 1704.280 ;
        RECT 1686.945 1704.000 1688.405 1704.280 ;
        RECT 1689.245 1704.000 1690.705 1704.280 ;
        RECT 1691.545 1704.000 1693.465 1704.280 ;
        RECT 1694.305 1704.000 1695.765 1704.280 ;
        RECT 1696.605 1704.000 1698.065 1704.280 ;
        RECT 1698.905 1704.000 1700.825 1704.280 ;
        RECT 1701.665 1704.000 1703.125 1704.280 ;
        RECT 1703.965 1704.000 1705.425 1704.280 ;
        RECT 1706.265 1704.000 1707.725 1704.280 ;
        RECT 1708.565 1704.000 1710.485 1704.280 ;
        RECT 1711.325 1704.000 1712.785 1704.280 ;
        RECT 1713.625 1704.000 1715.085 1704.280 ;
        RECT 1715.925 1704.000 1717.845 1704.280 ;
        RECT 1718.685 1704.000 1720.145 1704.280 ;
        RECT 1720.985 1704.000 1722.445 1704.280 ;
        RECT 1723.285 1704.000 1725.205 1704.280 ;
        RECT 1726.045 1704.000 1727.505 1704.280 ;
        RECT 1728.345 1704.000 1729.805 1704.280 ;
        RECT 1730.645 1704.000 1732.565 1704.280 ;
        RECT 1733.405 1704.000 1734.865 1704.280 ;
        RECT 1735.705 1704.000 1737.165 1704.280 ;
        RECT 1738.005 1704.000 1739.925 1704.280 ;
        RECT 1740.765 1704.000 1742.225 1704.280 ;
        RECT 1743.065 1704.000 1744.525 1704.280 ;
        RECT 1745.365 1704.000 1747.285 1704.280 ;
        RECT 1748.125 1704.000 1749.585 1704.280 ;
        RECT 1750.425 1704.000 1751.885 1704.280 ;
        RECT 1752.725 1704.000 1754.645 1704.280 ;
        RECT 1755.485 1704.000 1756.945 1704.280 ;
        RECT 1757.785 1704.000 1759.245 1704.280 ;
        RECT 1760.085 1704.000 1762.005 1704.280 ;
        RECT 1762.845 1704.000 1764.305 1704.280 ;
        RECT 1765.145 1704.000 1766.605 1704.280 ;
        RECT 1767.445 1704.000 1769.365 1704.280 ;
        RECT 1770.205 1704.000 1771.665 1704.280 ;
        RECT 1772.505 1704.000 1773.965 1704.280 ;
        RECT 1774.805 1704.000 1776.725 1704.280 ;
        RECT 1777.565 1704.000 1779.025 1704.280 ;
        RECT 1779.865 1704.000 1781.325 1704.280 ;
        RECT 1782.165 1704.000 1784.085 1704.280 ;
        RECT 1784.925 1704.000 1786.385 1704.280 ;
        RECT 1787.225 1704.000 1788.685 1704.280 ;
        RECT 1789.525 1704.000 1791.445 1704.280 ;
        RECT 1792.285 1704.000 1793.745 1704.280 ;
        RECT 1794.585 1704.000 1796.045 1704.280 ;
        RECT 1796.885 1704.000 1798.345 1704.280 ;
        RECT 1799.185 1704.000 1801.105 1704.280 ;
        RECT 1801.945 1704.000 1803.405 1704.280 ;
        RECT 1804.245 1704.000 1805.705 1704.280 ;
        RECT 1806.545 1704.000 1808.465 1704.280 ;
        RECT 1809.305 1704.000 1810.765 1704.280 ;
        RECT 1811.605 1704.000 1813.065 1704.280 ;
        RECT 1813.905 1704.000 1815.825 1704.280 ;
        RECT 1816.665 1704.000 1818.125 1704.280 ;
        RECT 1818.965 1704.000 1820.425 1704.280 ;
        RECT 1821.265 1704.000 1823.185 1704.280 ;
        RECT 1824.025 1704.000 1825.485 1704.280 ;
        RECT 1826.325 1704.000 1827.785 1704.280 ;
        RECT 1828.625 1704.000 1830.545 1704.280 ;
        RECT 1831.385 1704.000 1832.845 1704.280 ;
        RECT 1833.685 1704.000 1835.145 1704.280 ;
        RECT 1835.985 1704.000 1837.905 1704.280 ;
        RECT 1838.745 1704.000 1840.205 1704.280 ;
        RECT 1841.045 1704.000 1842.505 1704.280 ;
        RECT 1843.345 1704.000 1845.265 1704.280 ;
        RECT 1846.105 1704.000 1847.565 1704.280 ;
        RECT 1848.405 1704.000 1849.865 1704.280 ;
        RECT 1850.705 1704.000 1852.625 1704.280 ;
        RECT 1853.465 1704.000 1854.925 1704.280 ;
        RECT 1855.765 1704.000 1857.225 1704.280 ;
        RECT 1858.065 1704.000 1859.985 1704.280 ;
        RECT 1860.825 1704.000 1862.285 1704.280 ;
        RECT 1863.125 1704.000 1864.585 1704.280 ;
        RECT 1865.425 1704.000 1867.345 1704.280 ;
        RECT 1868.185 1704.000 1869.645 1704.280 ;
        RECT 1870.485 1704.000 1871.945 1704.280 ;
        RECT 1872.785 1704.000 1874.705 1704.280 ;
        RECT 1875.545 1704.000 1877.005 1704.280 ;
        RECT 1877.845 1704.000 1879.305 1704.280 ;
        RECT 1880.145 1704.000 1882.065 1704.280 ;
        RECT 1882.905 1704.000 1884.365 1704.280 ;
        RECT 1885.205 1704.000 1886.665 1704.280 ;
        RECT 1887.505 1704.000 1888.965 1704.280 ;
        RECT 1889.805 1704.000 1891.725 1704.280 ;
        RECT 1892.565 1704.000 1894.025 1704.280 ;
        RECT 1894.865 1704.000 1896.325 1704.280 ;
        RECT 1897.165 1704.000 1899.085 1704.280 ;
        RECT 1899.925 1704.000 1901.385 1704.280 ;
        RECT 1902.225 1704.000 1903.685 1704.280 ;
        RECT 1904.525 1704.000 1906.445 1704.280 ;
        RECT 1907.285 1704.000 1908.745 1704.280 ;
        RECT 1909.585 1704.000 1911.045 1704.280 ;
        RECT 1911.885 1704.000 1913.805 1704.280 ;
        RECT 1914.645 1704.000 1916.105 1704.280 ;
        RECT 1916.945 1704.000 1918.405 1704.280 ;
        RECT 1919.245 1704.000 1921.165 1704.280 ;
        RECT 1922.005 1704.000 1923.465 1704.280 ;
        RECT 1924.305 1704.000 1925.765 1704.280 ;
        RECT 1926.605 1704.000 1928.525 1704.280 ;
        RECT 1929.365 1704.000 1930.825 1704.280 ;
        RECT 1931.665 1704.000 1933.125 1704.280 ;
        RECT 1933.965 1704.000 1935.885 1704.280 ;
        RECT 1936.725 1704.000 1938.185 1704.280 ;
        RECT 1939.025 1704.000 1940.485 1704.280 ;
        RECT 1941.325 1704.000 1943.245 1704.280 ;
        RECT 1944.085 1704.000 1945.545 1704.280 ;
        RECT 1946.385 1704.000 1947.845 1704.280 ;
        RECT 1948.685 1704.000 1950.605 1704.280 ;
        RECT 1951.445 1704.000 1952.905 1704.280 ;
        RECT 1953.745 1704.000 1955.205 1704.280 ;
        RECT 1956.045 1704.000 1957.965 1704.280 ;
        RECT 1958.805 1704.000 1960.265 1704.280 ;
        RECT 1961.105 1704.000 1962.565 1704.280 ;
        RECT 1963.405 1704.000 1965.325 1704.280 ;
        RECT 1966.165 1704.000 1967.625 1704.280 ;
        RECT 1968.465 1704.000 1969.925 1704.280 ;
        RECT 1970.765 1704.000 1972.685 1704.280 ;
        RECT 1973.525 1704.000 1974.985 1704.280 ;
        RECT 1975.825 1704.000 1977.285 1704.280 ;
        RECT 1978.125 1704.000 1980.045 1704.280 ;
        RECT 1980.885 1704.000 1982.345 1704.280 ;
        RECT 1983.185 1704.000 1984.645 1704.280 ;
        RECT 1985.485 1704.000 1986.945 1704.280 ;
        RECT 1987.785 1704.000 1989.705 1704.280 ;
        RECT 1990.545 1704.000 1992.005 1704.280 ;
        RECT 1992.845 1704.000 1994.305 1704.280 ;
        RECT 1995.145 1704.000 1997.065 1704.280 ;
        RECT 1997.905 1704.000 1999.365 1704.280 ;
        RECT 2000.205 1704.000 2001.665 1704.280 ;
        RECT 2002.505 1704.000 2004.425 1704.280 ;
        RECT 2005.265 1704.000 2006.725 1704.280 ;
        RECT 2007.565 1704.000 2009.025 1704.280 ;
        RECT 2009.865 1704.000 2011.785 1704.280 ;
        RECT 2012.625 1704.000 2014.085 1704.280 ;
        RECT 2014.925 1704.000 2016.385 1704.280 ;
        RECT 2017.225 1704.000 2019.145 1704.280 ;
        RECT 2019.985 1704.000 2021.445 1704.280 ;
        RECT 2022.285 1704.000 2023.745 1704.280 ;
        RECT 2024.585 1704.000 2026.505 1704.280 ;
        RECT 2027.345 1704.000 2028.805 1704.280 ;
        RECT 2029.645 1704.000 2031.105 1704.280 ;
        RECT 2031.945 1704.000 2033.865 1704.280 ;
        RECT 2034.705 1704.000 2036.165 1704.280 ;
        RECT 2037.005 1704.000 2038.465 1704.280 ;
        RECT 2039.305 1704.000 2041.225 1704.280 ;
        RECT 2042.065 1704.000 2043.525 1704.280 ;
        RECT 2044.365 1704.000 2045.825 1704.280 ;
        RECT 2046.665 1704.000 2048.585 1704.280 ;
        RECT 2049.425 1704.000 2050.885 1704.280 ;
        RECT 2051.725 1704.000 2053.185 1704.280 ;
        RECT 2054.025 1704.000 2055.945 1704.280 ;
        RECT 2056.785 1704.000 2058.245 1704.280 ;
        RECT 2059.085 1704.000 2060.545 1704.280 ;
        RECT 2061.385 1704.000 2063.305 1704.280 ;
        RECT 2064.145 1704.000 2065.605 1704.280 ;
        RECT 2066.445 1704.000 2067.905 1704.280 ;
        RECT 2068.745 1704.000 2070.665 1704.280 ;
        RECT 2071.505 1704.000 2072.965 1704.280 ;
        RECT 2073.805 1704.000 2075.265 1704.280 ;
        RECT 2076.105 1704.000 2077.565 1704.280 ;
        RECT 2078.405 1704.000 2080.325 1704.280 ;
        RECT 2081.165 1704.000 2082.625 1704.280 ;
        RECT 2083.465 1704.000 2084.925 1704.280 ;
        RECT 2085.765 1704.000 2087.685 1704.280 ;
        RECT 2088.525 1704.000 2089.985 1704.280 ;
        RECT 2090.825 1704.000 2092.285 1704.280 ;
        RECT 2093.125 1704.000 2095.045 1704.280 ;
        RECT 2095.885 1704.000 2097.345 1704.280 ;
        RECT 2098.185 1704.000 2099.645 1704.280 ;
        RECT 2100.485 1704.000 2102.405 1704.280 ;
        RECT 2103.245 1704.000 2104.705 1704.280 ;
        RECT 2105.545 1704.000 2107.005 1704.280 ;
        RECT 2107.845 1704.000 2109.765 1704.280 ;
        RECT 2110.605 1704.000 2112.065 1704.280 ;
        RECT 2112.905 1704.000 2114.365 1704.280 ;
        RECT 2115.205 1704.000 2117.125 1704.280 ;
        RECT 2117.965 1704.000 2119.425 1704.280 ;
        RECT 2120.265 1704.000 2121.725 1704.280 ;
        RECT 2122.565 1704.000 2124.485 1704.280 ;
        RECT 2125.325 1704.000 2126.785 1704.280 ;
        RECT 2127.625 1704.000 2129.085 1704.280 ;
        RECT 2129.925 1704.000 2131.845 1704.280 ;
        RECT 2132.685 1704.000 2134.145 1704.280 ;
        RECT 2134.985 1704.000 2136.445 1704.280 ;
        RECT 2137.285 1704.000 2139.205 1704.280 ;
        RECT 2140.045 1704.000 2141.505 1704.280 ;
        RECT 2142.345 1704.000 2143.805 1704.280 ;
        RECT 2144.645 1704.000 2146.565 1704.280 ;
        RECT 2147.405 1704.000 2148.865 1704.280 ;
        RECT 2149.705 1704.000 2151.165 1704.280 ;
        RECT 2152.005 1704.000 2153.925 1704.280 ;
        RECT 2154.765 1704.000 2156.225 1704.280 ;
        RECT 2157.065 1704.000 2158.525 1704.280 ;
        RECT 2159.365 1704.000 2161.285 1704.280 ;
        RECT 2162.125 1704.000 2163.585 1704.280 ;
        RECT 2164.425 1704.000 2165.885 1704.280 ;
        RECT 2166.725 1704.000 2168.185 1704.280 ;
        RECT 2169.025 1704.000 2170.945 1704.280 ;
        RECT 2171.785 1704.000 2173.245 1704.280 ;
        RECT 2174.085 1704.000 2175.545 1704.280 ;
        RECT 2176.385 1704.000 2178.305 1704.280 ;
        RECT 2179.145 1704.000 2180.605 1704.280 ;
        RECT 2181.445 1704.000 2182.905 1704.280 ;
        RECT 2183.745 1704.000 2185.665 1704.280 ;
        RECT 2186.505 1704.000 2187.965 1704.280 ;
        RECT 2188.805 1704.000 2190.265 1704.280 ;
        RECT 2191.105 1704.000 2193.025 1704.280 ;
        RECT 2193.865 1704.000 2195.325 1704.280 ;
        RECT 2196.165 1704.000 2197.625 1704.280 ;
        RECT 2198.465 1704.000 2200.385 1704.280 ;
        RECT 2201.225 1704.000 2202.685 1704.280 ;
        RECT 2203.525 1704.000 2204.985 1704.280 ;
        RECT 2205.825 1704.000 2207.745 1704.280 ;
        RECT 2208.585 1704.000 2210.045 1704.280 ;
        RECT 2210.885 1704.000 2212.345 1704.280 ;
        RECT 2213.185 1704.000 2215.105 1704.280 ;
        RECT 2215.945 1704.000 2217.405 1704.280 ;
        RECT 2218.245 1704.000 2219.705 1704.280 ;
        RECT 2220.545 1704.000 2222.465 1704.280 ;
        RECT 2223.305 1704.000 2224.765 1704.280 ;
        RECT 2225.605 1704.000 2227.065 1704.280 ;
        RECT 2227.905 1704.000 2229.825 1704.280 ;
        RECT 2230.665 1704.000 2232.125 1704.280 ;
        RECT 2232.965 1704.000 2234.425 1704.280 ;
        RECT 2235.265 1704.000 2237.185 1704.280 ;
        RECT 2238.025 1704.000 2239.485 1704.280 ;
        RECT 2240.325 1704.000 2241.785 1704.280 ;
        RECT 2242.625 1704.000 2244.545 1704.280 ;
        RECT 2245.385 1704.000 2246.845 1704.280 ;
        RECT 2247.685 1704.000 2249.145 1704.280 ;
        RECT 2249.985 1704.000 2251.905 1704.280 ;
        RECT 2252.745 1704.000 2254.205 1704.280 ;
        RECT 2255.045 1704.000 2256.505 1704.280 ;
        RECT 2257.345 1704.000 2258.805 1704.280 ;
        RECT 2259.645 1704.000 2261.565 1704.280 ;
        RECT 2262.405 1704.000 2263.865 1704.280 ;
        RECT 2264.705 1704.000 2266.165 1704.280 ;
        RECT 2267.005 1704.000 2268.925 1704.280 ;
        RECT 2269.765 1704.000 2271.225 1704.280 ;
        RECT 2272.065 1704.000 2273.525 1704.280 ;
        RECT 2274.365 1704.000 2276.285 1704.280 ;
        RECT 2277.125 1704.000 2278.585 1704.280 ;
        RECT 2279.425 1704.000 2280.885 1704.280 ;
        RECT 2281.725 1704.000 2283.645 1704.280 ;
        RECT 2284.485 1704.000 2285.945 1704.280 ;
        RECT 2286.785 1704.000 2288.245 1704.280 ;
        RECT 2289.085 1704.000 2291.005 1704.280 ;
        RECT 2291.845 1704.000 2293.305 1704.280 ;
        RECT 2294.145 1704.000 2295.605 1704.280 ;
        RECT 2296.445 1704.000 2298.365 1704.280 ;
        RECT 2299.205 1704.000 2300.665 1704.280 ;
        RECT 2301.505 1704.000 2302.965 1704.280 ;
        RECT 2303.805 1704.000 2305.725 1704.280 ;
        RECT 2306.565 1704.000 2308.025 1704.280 ;
        RECT 2308.865 1704.000 2310.325 1704.280 ;
        RECT 2311.165 1704.000 2313.085 1704.280 ;
        RECT 2313.925 1704.000 2315.385 1704.280 ;
        RECT 2316.225 1704.000 2317.685 1704.280 ;
        RECT 2318.525 1704.000 2320.445 1704.280 ;
        RECT 2321.285 1704.000 2322.745 1704.280 ;
        RECT 2323.585 1704.000 2325.045 1704.280 ;
        RECT 2325.885 1704.000 2327.805 1704.280 ;
        RECT 2328.645 1704.000 2330.105 1704.280 ;
        RECT 2330.945 1704.000 2332.405 1704.280 ;
        RECT 2333.245 1704.000 2335.165 1704.280 ;
        RECT 2336.005 1704.000 2337.465 1704.280 ;
        RECT 2338.305 1704.000 2339.765 1704.280 ;
        RECT 2340.605 1704.000 2342.525 1704.280 ;
        RECT 2343.365 1704.000 2344.825 1704.280 ;
        RECT 2345.665 1704.000 2347.125 1704.280 ;
      LAYER met3 ;
        RECT 1150.000 1704.255 2327.930 2888.805 ;
      LAYER met4 ;
        RECT 1170.055 1710.640 1171.655 2888.880 ;
      LAYER met4 ;
        RECT 1245.910 1710.640 1246.455 2888.880 ;
      LAYER met4 ;
        RECT 1246.855 1710.640 1248.455 2888.880 ;
      LAYER met4 ;
        RECT 1248.855 1710.640 1264.020 2888.880 ;
        RECT 1267.020 1710.640 1282.020 2888.880 ;
        RECT 1285.020 1710.640 1300.020 2888.880 ;
        RECT 1303.020 1710.640 1318.020 2888.880 ;
        RECT 1321.020 1710.640 1354.020 2888.880 ;
        RECT 1357.020 1710.640 1372.020 2888.880 ;
        RECT 1375.020 1710.640 1390.020 2888.880 ;
        RECT 1393.020 1710.640 1408.020 2888.880 ;
        RECT 1411.020 1710.640 1444.020 2888.880 ;
        RECT 1447.020 1710.640 1462.020 2888.880 ;
        RECT 1465.020 1710.640 1480.020 2888.880 ;
        RECT 1483.020 1710.640 1498.020 2888.880 ;
        RECT 1501.020 1710.640 1534.020 2888.880 ;
        RECT 1537.020 1710.640 1552.020 2888.880 ;
        RECT 1555.020 1710.640 1570.020 2888.880 ;
        RECT 1573.020 1710.640 1588.020 2888.880 ;
        RECT 1591.020 1710.640 1624.020 2888.880 ;
        RECT 1627.020 1710.640 1642.020 2888.880 ;
        RECT 1645.020 1710.640 1660.020 2888.880 ;
        RECT 1663.020 1710.640 1678.020 2888.880 ;
        RECT 1681.020 1710.640 1714.020 2888.880 ;
        RECT 1717.020 1710.640 1732.020 2888.880 ;
        RECT 1735.020 1710.640 1750.020 2888.880 ;
        RECT 1753.020 1710.640 1768.020 2888.880 ;
        RECT 1771.020 1710.640 1804.020 2888.880 ;
        RECT 1807.020 1710.640 1822.020 2888.880 ;
        RECT 1825.020 1710.640 1840.020 2888.880 ;
        RECT 1843.020 1710.640 1858.020 2888.880 ;
        RECT 1861.020 1710.640 1894.020 2888.880 ;
        RECT 1897.020 1710.640 1912.020 2888.880 ;
        RECT 1915.020 1710.640 1930.020 2888.880 ;
        RECT 1933.020 1710.640 1948.020 2888.880 ;
        RECT 1951.020 1710.640 1984.020 2888.880 ;
        RECT 1987.020 1710.640 2002.020 2888.880 ;
        RECT 2005.020 1710.640 2020.020 2888.880 ;
        RECT 2023.020 1710.640 2038.020 2888.880 ;
        RECT 2041.020 1710.640 2074.020 2888.880 ;
        RECT 2077.020 1710.640 2092.020 2888.880 ;
        RECT 2095.020 1710.640 2110.020 2888.880 ;
        RECT 2113.020 1710.640 2128.020 2888.880 ;
        RECT 2131.020 1710.640 2164.020 2888.880 ;
        RECT 2167.020 1710.640 2182.020 2888.880 ;
        RECT 2185.020 1710.640 2200.020 2888.880 ;
        RECT 2203.020 1710.640 2218.020 2888.880 ;
        RECT 2221.020 1710.640 2254.020 2888.880 ;
        RECT 2257.020 1710.640 2272.020 2888.880 ;
        RECT 2275.020 1710.640 2290.020 2888.880 ;
        RECT 2293.020 1710.640 2308.020 2888.880 ;
        RECT 2311.020 1710.640 2323.655 2888.880 ;
  END
END user_project_wrapper
END LIBRARY

