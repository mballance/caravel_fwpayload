VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1497.160 BY 1500.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 5.080 1496.000 5.360 1500.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 399.760 1496.000 400.040 1500.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 438.860 1496.000 439.140 1500.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.420 1496.000 478.700 1500.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 517.980 1496.000 518.260 1500.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 557.540 1496.000 557.820 1500.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.100 1496.000 597.380 1500.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 636.660 1496.000 636.940 1500.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 675.760 1496.000 676.040 1500.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 715.320 1496.000 715.600 1500.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 754.880 1496.000 755.160 1500.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.180 1496.000 44.460 1500.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 794.440 1496.000 794.720 1500.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 834.000 1496.000 834.280 1500.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 873.100 1496.000 873.380 1500.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.660 1496.000 912.940 1500.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 952.220 1496.000 952.500 1500.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 991.780 1496.000 992.060 1500.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1031.340 1496.000 1031.620 1500.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1070.900 1496.000 1071.180 1500.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.000 1496.000 1110.280 1500.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1149.560 1496.000 1149.840 1500.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.740 1496.000 84.020 1500.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1189.120 1496.000 1189.400 1500.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1228.680 1496.000 1228.960 1500.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1268.240 1496.000 1268.520 1500.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1307.340 1496.000 1307.620 1500.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.900 1496.000 1347.180 1500.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1386.460 1496.000 1386.740 1500.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1426.020 1496.000 1426.300 1500.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1465.580 1496.000 1465.860 1500.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.300 1496.000 123.580 1500.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 162.860 1496.000 163.140 1500.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.420 1496.000 202.700 1500.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 241.520 1496.000 241.800 1500.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.080 1496.000 281.360 1500.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 320.640 1496.000 320.920 1500.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 360.200 1496.000 360.480 1500.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.960 1496.000 18.240 1500.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 412.640 1496.000 412.920 1500.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 452.200 1496.000 452.480 1500.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 491.760 1496.000 492.040 1500.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 531.320 1496.000 531.600 1500.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 570.880 1496.000 571.160 1500.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 609.980 1496.000 610.260 1500.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 649.540 1496.000 649.820 1500.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 689.100 1496.000 689.380 1500.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.660 1496.000 728.940 1500.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 768.220 1496.000 768.500 1500.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 57.520 1496.000 57.800 1500.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 807.320 1496.000 807.600 1500.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 846.880 1496.000 847.160 1500.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 886.440 1496.000 886.720 1500.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 926.000 1496.000 926.280 1500.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 965.560 1496.000 965.840 1500.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1005.120 1496.000 1005.400 1500.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1044.220 1496.000 1044.500 1500.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1083.780 1496.000 1084.060 1500.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1123.340 1496.000 1123.620 1500.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1162.900 1496.000 1163.180 1500.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 97.080 1496.000 97.360 1500.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1202.460 1496.000 1202.740 1500.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1241.560 1496.000 1241.840 1500.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.120 1496.000 1281.400 1500.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1320.680 1496.000 1320.960 1500.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1360.240 1496.000 1360.520 1500.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1399.800 1496.000 1400.080 1500.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1438.900 1496.000 1439.180 1500.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1478.460 1496.000 1478.740 1500.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 136.640 1496.000 136.920 1500.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 175.740 1496.000 176.020 1500.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 215.300 1496.000 215.580 1500.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 254.860 1496.000 255.140 1500.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 294.420 1496.000 294.700 1500.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 333.980 1496.000 334.260 1500.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 373.080 1496.000 373.360 1500.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 31.300 1496.000 31.580 1500.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 425.980 1496.000 426.260 1500.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 465.540 1496.000 465.820 1500.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 505.100 1496.000 505.380 1500.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 544.200 1496.000 544.480 1500.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 583.760 1496.000 584.040 1500.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 623.320 1496.000 623.600 1500.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 662.880 1496.000 663.160 1500.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 702.440 1496.000 702.720 1500.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 741.540 1496.000 741.820 1500.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 781.100 1496.000 781.380 1500.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.860 1496.000 71.140 1500.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 820.660 1496.000 820.940 1500.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 860.220 1496.000 860.500 1500.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 899.780 1496.000 900.060 1500.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 938.880 1496.000 939.160 1500.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 978.440 1496.000 978.720 1500.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1018.000 1496.000 1018.280 1500.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1057.560 1496.000 1057.840 1500.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1097.120 1496.000 1097.400 1500.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1136.680 1496.000 1136.960 1500.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1175.780 1496.000 1176.060 1500.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.960 1496.000 110.240 1500.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1215.340 1496.000 1215.620 1500.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1254.900 1496.000 1255.180 1500.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1294.460 1496.000 1294.740 1500.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1334.020 1496.000 1334.300 1500.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1373.120 1496.000 1373.400 1500.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1412.680 1496.000 1412.960 1500.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1452.240 1496.000 1452.520 1500.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1491.800 1496.000 1492.080 1500.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.520 1496.000 149.800 1500.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 189.080 1496.000 189.360 1500.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 228.640 1496.000 228.920 1500.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 268.200 1496.000 268.480 1500.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 307.300 1496.000 307.580 1500.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 346.860 1496.000 347.140 1500.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 386.420 1496.000 386.700 1500.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 324.320 0.000 324.600 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1242.480 0.000 1242.760 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1251.680 0.000 1251.960 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1260.880 0.000 1261.160 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1270.080 0.000 1270.360 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1279.280 0.000 1279.560 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1288.480 0.000 1288.760 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1297.680 0.000 1297.960 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1306.880 0.000 1307.160 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1316.080 0.000 1316.360 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1325.280 0.000 1325.560 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 416.320 0.000 416.600 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1334.480 0.000 1334.760 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1343.680 0.000 1343.960 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1352.880 0.000 1353.160 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1362.080 0.000 1362.360 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1371.280 0.000 1371.560 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1380.480 0.000 1380.760 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1389.680 0.000 1389.960 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1398.880 0.000 1399.160 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1408.080 0.000 1408.360 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1417.280 0.000 1417.560 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 425.520 0.000 425.800 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1426.480 0.000 1426.760 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1435.680 0.000 1435.960 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1444.880 0.000 1445.160 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1454.080 0.000 1454.360 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1463.280 0.000 1463.560 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1472.480 0.000 1472.760 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1481.680 0.000 1481.960 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1490.880 0.000 1491.160 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 434.720 0.000 435.000 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.460 0.000 443.740 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 452.660 0.000 452.940 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.860 0.000 462.140 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.060 0.000 471.340 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 480.260 0.000 480.540 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 489.460 0.000 489.740 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 498.660 0.000 498.940 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 333.520 0.000 333.800 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 507.860 0.000 508.140 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 517.060 0.000 517.340 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 526.260 0.000 526.540 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 535.460 0.000 535.740 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 544.660 0.000 544.940 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 553.860 0.000 554.140 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 563.060 0.000 563.340 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 572.260 0.000 572.540 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 581.460 0.000 581.740 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 590.660 0.000 590.940 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 342.720 0.000 343.000 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 599.860 0.000 600.140 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 609.060 0.000 609.340 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 618.260 0.000 618.540 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.460 0.000 627.740 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 636.660 0.000 636.940 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 645.860 0.000 646.140 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 655.060 0.000 655.340 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 664.260 0.000 664.540 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 673.460 0.000 673.740 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 682.660 0.000 682.940 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 351.920 0.000 352.200 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 691.860 0.000 692.140 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 701.060 0.000 701.340 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 709.800 0.000 710.080 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 719.000 0.000 719.280 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 728.200 0.000 728.480 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 737.400 0.000 737.680 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 746.600 0.000 746.880 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 755.800 0.000 756.080 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 765.000 0.000 765.280 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 774.200 0.000 774.480 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 361.120 0.000 361.400 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.400 0.000 783.680 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 792.600 0.000 792.880 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 801.800 0.000 802.080 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.000 0.000 811.280 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 820.200 0.000 820.480 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.400 0.000 829.680 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 838.600 0.000 838.880 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 847.800 0.000 848.080 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 857.000 0.000 857.280 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.200 0.000 866.480 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 370.320 0.000 370.600 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 875.400 0.000 875.680 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 884.600 0.000 884.880 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 893.800 0.000 894.080 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 903.000 0.000 903.280 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 912.200 0.000 912.480 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 921.400 0.000 921.680 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 930.600 0.000 930.880 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 939.800 0.000 940.080 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.000 0.000 949.280 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 958.200 0.000 958.480 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 379.520 0.000 379.800 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 967.400 0.000 967.680 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 976.140 0.000 976.420 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 985.340 0.000 985.620 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 994.540 0.000 994.820 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1003.740 0.000 1004.020 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1012.940 0.000 1013.220 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1022.140 0.000 1022.420 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1031.340 0.000 1031.620 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1040.540 0.000 1040.820 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1049.740 0.000 1050.020 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 388.720 0.000 389.000 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1058.940 0.000 1059.220 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1068.140 0.000 1068.420 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1077.340 0.000 1077.620 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1086.540 0.000 1086.820 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1095.740 0.000 1096.020 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1104.940 0.000 1105.220 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1114.140 0.000 1114.420 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1123.340 0.000 1123.620 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1132.540 0.000 1132.820 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1141.740 0.000 1142.020 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 397.920 0.000 398.200 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1150.940 0.000 1151.220 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1160.140 0.000 1160.420 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1169.340 0.000 1169.620 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1178.540 0.000 1178.820 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1187.740 0.000 1188.020 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1196.940 0.000 1197.220 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1206.140 0.000 1206.420 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.340 0.000 1215.620 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1224.540 0.000 1224.820 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.740 0.000 1234.020 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 407.120 0.000 407.400 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 327.540 0.000 327.820 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1245.700 0.000 1245.980 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1254.900 0.000 1255.180 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1264.100 0.000 1264.380 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1273.300 0.000 1273.580 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1282.500 0.000 1282.780 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1291.700 0.000 1291.980 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1300.900 0.000 1301.180 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1310.100 0.000 1310.380 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1319.300 0.000 1319.580 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1328.500 0.000 1328.780 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 419.080 0.000 419.360 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1337.700 0.000 1337.980 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1346.900 0.000 1347.180 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1356.100 0.000 1356.380 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1365.300 0.000 1365.580 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1374.500 0.000 1374.780 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1383.700 0.000 1383.980 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1392.900 0.000 1393.180 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1402.100 0.000 1402.380 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1411.300 0.000 1411.580 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1420.040 0.000 1420.320 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 428.280 0.000 428.560 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1429.240 0.000 1429.520 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1438.440 0.000 1438.720 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1447.640 0.000 1447.920 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1456.840 0.000 1457.120 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1466.040 0.000 1466.320 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1475.240 0.000 1475.520 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1484.440 0.000 1484.720 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1493.640 0.000 1493.920 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 437.480 0.000 437.760 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 446.680 0.000 446.960 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 455.880 0.000 456.160 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 465.080 0.000 465.360 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 474.280 0.000 474.560 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 483.480 0.000 483.760 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 492.680 0.000 492.960 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 501.880 0.000 502.160 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 336.740 0.000 337.020 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 511.080 0.000 511.360 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 520.280 0.000 520.560 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 529.480 0.000 529.760 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 538.680 0.000 538.960 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 547.880 0.000 548.160 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 557.080 0.000 557.360 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 566.280 0.000 566.560 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 575.480 0.000 575.760 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 584.680 0.000 584.960 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 593.880 0.000 594.160 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 345.940 0.000 346.220 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 603.080 0.000 603.360 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 612.280 0.000 612.560 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 621.020 0.000 621.300 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 630.220 0.000 630.500 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 639.420 0.000 639.700 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 648.620 0.000 648.900 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 657.820 0.000 658.100 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 667.020 0.000 667.300 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 676.220 0.000 676.500 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 685.420 0.000 685.700 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.680 0.000 354.960 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 694.620 0.000 694.900 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 703.820 0.000 704.100 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 713.020 0.000 713.300 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 722.220 0.000 722.500 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 731.420 0.000 731.700 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 740.620 0.000 740.900 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 749.820 0.000 750.100 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 759.020 0.000 759.300 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 768.220 0.000 768.500 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 777.420 0.000 777.700 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 363.880 0.000 364.160 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 786.620 0.000 786.900 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 795.820 0.000 796.100 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 805.020 0.000 805.300 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 814.220 0.000 814.500 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 823.420 0.000 823.700 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 832.620 0.000 832.900 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 841.820 0.000 842.100 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 851.020 0.000 851.300 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 860.220 0.000 860.500 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 869.420 0.000 869.700 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 373.080 0.000 373.360 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 878.620 0.000 878.900 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 887.360 0.000 887.640 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 896.560 0.000 896.840 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 905.760 0.000 906.040 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 914.960 0.000 915.240 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 924.160 0.000 924.440 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 933.360 0.000 933.640 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 942.560 0.000 942.840 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 951.760 0.000 952.040 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 960.960 0.000 961.240 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 382.280 0.000 382.560 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 970.160 0.000 970.440 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 979.360 0.000 979.640 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 988.560 0.000 988.840 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 997.760 0.000 998.040 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1006.960 0.000 1007.240 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1016.160 0.000 1016.440 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1025.360 0.000 1025.640 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1034.560 0.000 1034.840 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1043.760 0.000 1044.040 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1052.960 0.000 1053.240 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 391.480 0.000 391.760 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1062.160 0.000 1062.440 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1071.360 0.000 1071.640 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1080.560 0.000 1080.840 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1089.760 0.000 1090.040 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1098.960 0.000 1099.240 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1108.160 0.000 1108.440 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1117.360 0.000 1117.640 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1126.560 0.000 1126.840 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1135.760 0.000 1136.040 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1144.960 0.000 1145.240 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 400.680 0.000 400.960 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1153.700 0.000 1153.980 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1162.900 0.000 1163.180 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1172.100 0.000 1172.380 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1181.300 0.000 1181.580 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1190.500 0.000 1190.780 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1199.700 0.000 1199.980 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1208.900 0.000 1209.180 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1218.100 0.000 1218.380 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1227.300 0.000 1227.580 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1236.500 0.000 1236.780 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.880 0.000 410.160 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 330.300 0.000 330.580 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1248.920 0.000 1249.200 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1258.120 0.000 1258.400 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1267.320 0.000 1267.600 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1276.520 0.000 1276.800 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1285.720 0.000 1286.000 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1294.920 0.000 1295.200 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1304.120 0.000 1304.400 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1313.320 0.000 1313.600 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1322.520 0.000 1322.800 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1331.260 0.000 1331.540 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 422.300 0.000 422.580 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1340.460 0.000 1340.740 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1349.660 0.000 1349.940 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1358.860 0.000 1359.140 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1368.060 0.000 1368.340 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1377.260 0.000 1377.540 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1386.460 0.000 1386.740 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1395.660 0.000 1395.940 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1404.860 0.000 1405.140 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1414.060 0.000 1414.340 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1423.260 0.000 1423.540 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 431.500 0.000 431.780 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1432.460 0.000 1432.740 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1441.660 0.000 1441.940 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1450.860 0.000 1451.140 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1460.060 0.000 1460.340 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1469.260 0.000 1469.540 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1478.460 0.000 1478.740 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1487.660 0.000 1487.940 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1496.860 0.000 1497.140 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 440.700 0.000 440.980 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 449.900 0.000 450.180 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 459.100 0.000 459.380 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 468.300 0.000 468.580 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.500 0.000 477.780 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 486.700 0.000 486.980 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 495.900 0.000 496.180 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 505.100 0.000 505.380 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 339.500 0.000 339.780 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 514.300 0.000 514.580 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 523.500 0.000 523.780 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 532.240 0.000 532.520 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 541.440 0.000 541.720 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 550.640 0.000 550.920 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 559.840 0.000 560.120 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 569.040 0.000 569.320 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 578.240 0.000 578.520 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.440 0.000 587.720 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 596.640 0.000 596.920 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 348.700 0.000 348.980 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 605.840 0.000 606.120 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 615.040 0.000 615.320 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 624.240 0.000 624.520 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 633.440 0.000 633.720 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 642.640 0.000 642.920 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 651.840 0.000 652.120 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 661.040 0.000 661.320 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 670.240 0.000 670.520 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 679.440 0.000 679.720 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 688.640 0.000 688.920 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.900 0.000 358.180 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 697.840 0.000 698.120 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 707.040 0.000 707.320 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 716.240 0.000 716.520 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 725.440 0.000 725.720 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.640 0.000 734.920 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 743.840 0.000 744.120 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 753.040 0.000 753.320 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 762.240 0.000 762.520 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 771.440 0.000 771.720 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 780.640 0.000 780.920 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 367.100 0.000 367.380 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 789.840 0.000 790.120 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 798.580 0.000 798.860 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 807.780 0.000 808.060 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 816.980 0.000 817.260 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 826.180 0.000 826.460 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 835.380 0.000 835.660 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 844.580 0.000 844.860 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 853.780 0.000 854.060 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 862.980 0.000 863.260 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 872.180 0.000 872.460 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 376.300 0.000 376.580 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 881.380 0.000 881.660 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 890.580 0.000 890.860 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 899.780 0.000 900.060 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 908.980 0.000 909.260 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.180 0.000 918.460 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 927.380 0.000 927.660 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 936.580 0.000 936.860 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 945.780 0.000 946.060 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 954.980 0.000 955.260 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 964.180 0.000 964.460 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 385.500 0.000 385.780 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 973.380 0.000 973.660 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 982.580 0.000 982.860 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 991.780 0.000 992.060 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1000.980 0.000 1001.260 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1010.180 0.000 1010.460 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1019.380 0.000 1019.660 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1028.580 0.000 1028.860 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1037.780 0.000 1038.060 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1046.980 0.000 1047.260 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1056.180 0.000 1056.460 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 394.700 0.000 394.980 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1064.920 0.000 1065.200 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1074.120 0.000 1074.400 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.320 0.000 1083.600 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1092.520 0.000 1092.800 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1101.720 0.000 1102.000 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1110.920 0.000 1111.200 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1120.120 0.000 1120.400 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1129.320 0.000 1129.600 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1138.520 0.000 1138.800 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1147.720 0.000 1148.000 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.900 0.000 404.180 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1156.920 0.000 1157.200 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1166.120 0.000 1166.400 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.320 0.000 1175.600 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1184.520 0.000 1184.800 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1193.720 0.000 1194.000 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1202.920 0.000 1203.200 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1212.120 0.000 1212.400 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1221.320 0.000 1221.600 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1230.520 0.000 1230.800 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1239.720 0.000 1240.000 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 413.100 0.000 413.380 4.000 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.780 0.000 3.060 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 6.000 0.000 6.280 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.960 0.000 18.240 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.380 0.000 122.660 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.580 0.000 131.860 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 140.780 0.000 141.060 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.980 0.000 150.260 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.180 0.000 159.460 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 168.380 0.000 168.660 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 177.120 0.000 177.400 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.320 0.000 186.600 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.520 0.000 195.800 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.720 0.000 205.000 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.380 0.000 30.660 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.920 0.000 214.200 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 223.120 0.000 223.400 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 232.320 0.000 232.600 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 241.520 0.000 241.800 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 250.720 0.000 251.000 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 259.920 0.000 260.200 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.120 0.000 269.400 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 278.320 0.000 278.600 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 287.520 0.000 287.800 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 296.720 0.000 297.000 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.800 0.000 43.080 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 305.920 0.000 306.200 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 315.120 0.000 315.400 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 54.760 0.000 55.040 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.180 0.000 67.460 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 76.380 0.000 76.660 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.580 0.000 85.860 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.780 0.000 95.060 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.980 0.000 104.260 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.180 0.000 113.460 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.760 0.000 9.040 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.180 0.000 21.460 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 125.140 0.000 125.420 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.340 0.000 134.620 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.540 0.000 143.820 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 152.740 0.000 153.020 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 161.940 0.000 162.220 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 171.140 0.000 171.420 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 180.340 0.000 180.620 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 189.540 0.000 189.820 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 198.740 0.000 199.020 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 207.940 0.000 208.220 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.600 0.000 33.880 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.140 0.000 217.420 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 226.340 0.000 226.620 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 235.540 0.000 235.820 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.740 0.000 245.020 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 253.940 0.000 254.220 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.140 0.000 263.420 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 272.340 0.000 272.620 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.540 0.000 281.820 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 290.740 0.000 291.020 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 299.940 0.000 300.220 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.560 0.000 45.840 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 309.140 0.000 309.420 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 318.340 0.000 318.620 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.980 0.000 58.260 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.400 0.000 70.680 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.600 0.000 79.880 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.340 0.000 88.620 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.540 0.000 97.820 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 106.740 0.000 107.020 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.940 0.000 116.220 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.400 0.000 24.680 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.360 0.000 128.640 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.560 0.000 137.840 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.760 0.000 147.040 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.960 0.000 156.240 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 165.160 0.000 165.440 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.360 0.000 174.640 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.560 0.000 183.840 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 192.760 0.000 193.040 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 201.960 0.000 202.240 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 211.160 0.000 211.440 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.360 0.000 36.640 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 220.360 0.000 220.640 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 229.560 0.000 229.840 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 238.760 0.000 239.040 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 247.960 0.000 248.240 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 257.160 0.000 257.440 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 265.900 0.000 266.180 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 275.100 0.000 275.380 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 284.300 0.000 284.580 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 293.500 0.000 293.780 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 302.700 0.000 302.980 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.780 0.000 49.060 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 311.900 0.000 312.180 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 321.100 0.000 321.380 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 61.200 0.000 61.480 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.160 0.000 73.440 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.360 0.000 82.640 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 91.560 0.000 91.840 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.760 0.000 101.040 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.960 0.000 110.240 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.160 0.000 119.440 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 27.160 0.000 27.440 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 39.580 0.000 39.860 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.000 0.000 52.280 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.960 0.000 64.240 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.980 0.000 12.260 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.200 0.000 15.480 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.590 10.640 21.190 1488.080 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.390 10.640 97.990 1488.080 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.070 10.795 1492.630 1487.925 ;
      LAYER met1 ;
        RECT 0.000 4.460 1497.160 1488.080 ;
      LAYER met2 ;
        RECT 0.030 1495.720 4.800 1496.000 ;
        RECT 5.640 1495.720 17.680 1496.000 ;
        RECT 18.520 1495.720 31.020 1496.000 ;
        RECT 31.860 1495.720 43.900 1496.000 ;
        RECT 44.740 1495.720 57.240 1496.000 ;
        RECT 58.080 1495.720 70.580 1496.000 ;
        RECT 71.420 1495.720 83.460 1496.000 ;
        RECT 84.300 1495.720 96.800 1496.000 ;
        RECT 97.640 1495.720 109.680 1496.000 ;
        RECT 110.520 1495.720 123.020 1496.000 ;
        RECT 123.860 1495.720 136.360 1496.000 ;
        RECT 137.200 1495.720 149.240 1496.000 ;
        RECT 150.080 1495.720 162.580 1496.000 ;
        RECT 163.420 1495.720 175.460 1496.000 ;
        RECT 176.300 1495.720 188.800 1496.000 ;
        RECT 189.640 1495.720 202.140 1496.000 ;
        RECT 202.980 1495.720 215.020 1496.000 ;
        RECT 215.860 1495.720 228.360 1496.000 ;
        RECT 229.200 1495.720 241.240 1496.000 ;
        RECT 242.080 1495.720 254.580 1496.000 ;
        RECT 255.420 1495.720 267.920 1496.000 ;
        RECT 268.760 1495.720 280.800 1496.000 ;
        RECT 281.640 1495.720 294.140 1496.000 ;
        RECT 294.980 1495.720 307.020 1496.000 ;
        RECT 307.860 1495.720 320.360 1496.000 ;
        RECT 321.200 1495.720 333.700 1496.000 ;
        RECT 334.540 1495.720 346.580 1496.000 ;
        RECT 347.420 1495.720 359.920 1496.000 ;
        RECT 360.760 1495.720 372.800 1496.000 ;
        RECT 373.640 1495.720 386.140 1496.000 ;
        RECT 386.980 1495.720 399.480 1496.000 ;
        RECT 400.320 1495.720 412.360 1496.000 ;
        RECT 413.200 1495.720 425.700 1496.000 ;
        RECT 426.540 1495.720 438.580 1496.000 ;
        RECT 439.420 1495.720 451.920 1496.000 ;
        RECT 452.760 1495.720 465.260 1496.000 ;
        RECT 466.100 1495.720 478.140 1496.000 ;
        RECT 478.980 1495.720 491.480 1496.000 ;
        RECT 492.320 1495.720 504.820 1496.000 ;
        RECT 505.660 1495.720 517.700 1496.000 ;
        RECT 518.540 1495.720 531.040 1496.000 ;
        RECT 531.880 1495.720 543.920 1496.000 ;
        RECT 544.760 1495.720 557.260 1496.000 ;
        RECT 558.100 1495.720 570.600 1496.000 ;
        RECT 571.440 1495.720 583.480 1496.000 ;
        RECT 584.320 1495.720 596.820 1496.000 ;
        RECT 597.660 1495.720 609.700 1496.000 ;
        RECT 610.540 1495.720 623.040 1496.000 ;
        RECT 623.880 1495.720 636.380 1496.000 ;
        RECT 637.220 1495.720 649.260 1496.000 ;
        RECT 650.100 1495.720 662.600 1496.000 ;
        RECT 663.440 1495.720 675.480 1496.000 ;
        RECT 676.320 1495.720 688.820 1496.000 ;
        RECT 689.660 1495.720 702.160 1496.000 ;
        RECT 703.000 1495.720 715.040 1496.000 ;
        RECT 715.880 1495.720 728.380 1496.000 ;
        RECT 729.220 1495.720 741.260 1496.000 ;
        RECT 742.100 1495.720 754.600 1496.000 ;
        RECT 755.440 1495.720 767.940 1496.000 ;
        RECT 768.780 1495.720 780.820 1496.000 ;
        RECT 781.660 1495.720 794.160 1496.000 ;
        RECT 795.000 1495.720 807.040 1496.000 ;
        RECT 807.880 1495.720 820.380 1496.000 ;
        RECT 821.220 1495.720 833.720 1496.000 ;
        RECT 834.560 1495.720 846.600 1496.000 ;
        RECT 847.440 1495.720 859.940 1496.000 ;
        RECT 860.780 1495.720 872.820 1496.000 ;
        RECT 873.660 1495.720 886.160 1496.000 ;
        RECT 887.000 1495.720 899.500 1496.000 ;
        RECT 900.340 1495.720 912.380 1496.000 ;
        RECT 913.220 1495.720 925.720 1496.000 ;
        RECT 926.560 1495.720 938.600 1496.000 ;
        RECT 939.440 1495.720 951.940 1496.000 ;
        RECT 952.780 1495.720 965.280 1496.000 ;
        RECT 966.120 1495.720 978.160 1496.000 ;
        RECT 979.000 1495.720 991.500 1496.000 ;
        RECT 992.340 1495.720 1004.840 1496.000 ;
        RECT 1005.680 1495.720 1017.720 1496.000 ;
        RECT 1018.560 1495.720 1031.060 1496.000 ;
        RECT 1031.900 1495.720 1043.940 1496.000 ;
        RECT 1044.780 1495.720 1057.280 1496.000 ;
        RECT 1058.120 1495.720 1070.620 1496.000 ;
        RECT 1071.460 1495.720 1083.500 1496.000 ;
        RECT 1084.340 1495.720 1096.840 1496.000 ;
        RECT 1097.680 1495.720 1109.720 1496.000 ;
        RECT 1110.560 1495.720 1123.060 1496.000 ;
        RECT 1123.900 1495.720 1136.400 1496.000 ;
        RECT 1137.240 1495.720 1149.280 1496.000 ;
        RECT 1150.120 1495.720 1162.620 1496.000 ;
        RECT 1163.460 1495.720 1175.500 1496.000 ;
        RECT 1176.340 1495.720 1188.840 1496.000 ;
        RECT 1189.680 1495.720 1202.180 1496.000 ;
        RECT 1203.020 1495.720 1215.060 1496.000 ;
        RECT 1215.900 1495.720 1228.400 1496.000 ;
        RECT 1229.240 1495.720 1241.280 1496.000 ;
        RECT 1242.120 1495.720 1254.620 1496.000 ;
        RECT 1255.460 1495.720 1267.960 1496.000 ;
        RECT 1268.800 1495.720 1280.840 1496.000 ;
        RECT 1281.680 1495.720 1294.180 1496.000 ;
        RECT 1295.020 1495.720 1307.060 1496.000 ;
        RECT 1307.900 1495.720 1320.400 1496.000 ;
        RECT 1321.240 1495.720 1333.740 1496.000 ;
        RECT 1334.580 1495.720 1346.620 1496.000 ;
        RECT 1347.460 1495.720 1359.960 1496.000 ;
        RECT 1360.800 1495.720 1372.840 1496.000 ;
        RECT 1373.680 1495.720 1386.180 1496.000 ;
        RECT 1387.020 1495.720 1399.520 1496.000 ;
        RECT 1400.360 1495.720 1412.400 1496.000 ;
        RECT 1413.240 1495.720 1425.740 1496.000 ;
        RECT 1426.580 1495.720 1438.620 1496.000 ;
        RECT 1439.460 1495.720 1451.960 1496.000 ;
        RECT 1452.800 1495.720 1465.300 1496.000 ;
        RECT 1466.140 1495.720 1478.180 1496.000 ;
        RECT 1479.020 1495.720 1491.520 1496.000 ;
        RECT 1492.360 1495.720 1497.130 1496.000 ;
        RECT 0.030 4.280 1497.130 1495.720 ;
        RECT 0.580 4.000 2.500 4.280 ;
        RECT 3.340 4.000 5.720 4.280 ;
        RECT 6.560 4.000 8.480 4.280 ;
        RECT 9.320 4.000 11.700 4.280 ;
        RECT 12.540 4.000 14.920 4.280 ;
        RECT 15.760 4.000 17.680 4.280 ;
        RECT 18.520 4.000 20.900 4.280 ;
        RECT 21.740 4.000 24.120 4.280 ;
        RECT 24.960 4.000 26.880 4.280 ;
        RECT 27.720 4.000 30.100 4.280 ;
        RECT 30.940 4.000 33.320 4.280 ;
        RECT 34.160 4.000 36.080 4.280 ;
        RECT 36.920 4.000 39.300 4.280 ;
        RECT 40.140 4.000 42.520 4.280 ;
        RECT 43.360 4.000 45.280 4.280 ;
        RECT 46.120 4.000 48.500 4.280 ;
        RECT 49.340 4.000 51.720 4.280 ;
        RECT 52.560 4.000 54.480 4.280 ;
        RECT 55.320 4.000 57.700 4.280 ;
        RECT 58.540 4.000 60.920 4.280 ;
        RECT 61.760 4.000 63.680 4.280 ;
        RECT 64.520 4.000 66.900 4.280 ;
        RECT 67.740 4.000 70.120 4.280 ;
        RECT 70.960 4.000 72.880 4.280 ;
        RECT 73.720 4.000 76.100 4.280 ;
        RECT 76.940 4.000 79.320 4.280 ;
        RECT 80.160 4.000 82.080 4.280 ;
        RECT 82.920 4.000 85.300 4.280 ;
        RECT 86.140 4.000 88.060 4.280 ;
        RECT 88.900 4.000 91.280 4.280 ;
        RECT 92.120 4.000 94.500 4.280 ;
        RECT 95.340 4.000 97.260 4.280 ;
        RECT 98.100 4.000 100.480 4.280 ;
        RECT 101.320 4.000 103.700 4.280 ;
        RECT 104.540 4.000 106.460 4.280 ;
        RECT 107.300 4.000 109.680 4.280 ;
        RECT 110.520 4.000 112.900 4.280 ;
        RECT 113.740 4.000 115.660 4.280 ;
        RECT 116.500 4.000 118.880 4.280 ;
        RECT 119.720 4.000 122.100 4.280 ;
        RECT 122.940 4.000 124.860 4.280 ;
        RECT 125.700 4.000 128.080 4.280 ;
        RECT 128.920 4.000 131.300 4.280 ;
        RECT 132.140 4.000 134.060 4.280 ;
        RECT 134.900 4.000 137.280 4.280 ;
        RECT 138.120 4.000 140.500 4.280 ;
        RECT 141.340 4.000 143.260 4.280 ;
        RECT 144.100 4.000 146.480 4.280 ;
        RECT 147.320 4.000 149.700 4.280 ;
        RECT 150.540 4.000 152.460 4.280 ;
        RECT 153.300 4.000 155.680 4.280 ;
        RECT 156.520 4.000 158.900 4.280 ;
        RECT 159.740 4.000 161.660 4.280 ;
        RECT 162.500 4.000 164.880 4.280 ;
        RECT 165.720 4.000 168.100 4.280 ;
        RECT 168.940 4.000 170.860 4.280 ;
        RECT 171.700 4.000 174.080 4.280 ;
        RECT 174.920 4.000 176.840 4.280 ;
        RECT 177.680 4.000 180.060 4.280 ;
        RECT 180.900 4.000 183.280 4.280 ;
        RECT 184.120 4.000 186.040 4.280 ;
        RECT 186.880 4.000 189.260 4.280 ;
        RECT 190.100 4.000 192.480 4.280 ;
        RECT 193.320 4.000 195.240 4.280 ;
        RECT 196.080 4.000 198.460 4.280 ;
        RECT 199.300 4.000 201.680 4.280 ;
        RECT 202.520 4.000 204.440 4.280 ;
        RECT 205.280 4.000 207.660 4.280 ;
        RECT 208.500 4.000 210.880 4.280 ;
        RECT 211.720 4.000 213.640 4.280 ;
        RECT 214.480 4.000 216.860 4.280 ;
        RECT 217.700 4.000 220.080 4.280 ;
        RECT 220.920 4.000 222.840 4.280 ;
        RECT 223.680 4.000 226.060 4.280 ;
        RECT 226.900 4.000 229.280 4.280 ;
        RECT 230.120 4.000 232.040 4.280 ;
        RECT 232.880 4.000 235.260 4.280 ;
        RECT 236.100 4.000 238.480 4.280 ;
        RECT 239.320 4.000 241.240 4.280 ;
        RECT 242.080 4.000 244.460 4.280 ;
        RECT 245.300 4.000 247.680 4.280 ;
        RECT 248.520 4.000 250.440 4.280 ;
        RECT 251.280 4.000 253.660 4.280 ;
        RECT 254.500 4.000 256.880 4.280 ;
        RECT 257.720 4.000 259.640 4.280 ;
        RECT 260.480 4.000 262.860 4.280 ;
        RECT 263.700 4.000 265.620 4.280 ;
        RECT 266.460 4.000 268.840 4.280 ;
        RECT 269.680 4.000 272.060 4.280 ;
        RECT 272.900 4.000 274.820 4.280 ;
        RECT 275.660 4.000 278.040 4.280 ;
        RECT 278.880 4.000 281.260 4.280 ;
        RECT 282.100 4.000 284.020 4.280 ;
        RECT 284.860 4.000 287.240 4.280 ;
        RECT 288.080 4.000 290.460 4.280 ;
        RECT 291.300 4.000 293.220 4.280 ;
        RECT 294.060 4.000 296.440 4.280 ;
        RECT 297.280 4.000 299.660 4.280 ;
        RECT 300.500 4.000 302.420 4.280 ;
        RECT 303.260 4.000 305.640 4.280 ;
        RECT 306.480 4.000 308.860 4.280 ;
        RECT 309.700 4.000 311.620 4.280 ;
        RECT 312.460 4.000 314.840 4.280 ;
        RECT 315.680 4.000 318.060 4.280 ;
        RECT 318.900 4.000 320.820 4.280 ;
        RECT 321.660 4.000 324.040 4.280 ;
        RECT 324.880 4.000 327.260 4.280 ;
        RECT 328.100 4.000 330.020 4.280 ;
        RECT 330.860 4.000 333.240 4.280 ;
        RECT 334.080 4.000 336.460 4.280 ;
        RECT 337.300 4.000 339.220 4.280 ;
        RECT 340.060 4.000 342.440 4.280 ;
        RECT 343.280 4.000 345.660 4.280 ;
        RECT 346.500 4.000 348.420 4.280 ;
        RECT 349.260 4.000 351.640 4.280 ;
        RECT 352.480 4.000 354.400 4.280 ;
        RECT 355.240 4.000 357.620 4.280 ;
        RECT 358.460 4.000 360.840 4.280 ;
        RECT 361.680 4.000 363.600 4.280 ;
        RECT 364.440 4.000 366.820 4.280 ;
        RECT 367.660 4.000 370.040 4.280 ;
        RECT 370.880 4.000 372.800 4.280 ;
        RECT 373.640 4.000 376.020 4.280 ;
        RECT 376.860 4.000 379.240 4.280 ;
        RECT 380.080 4.000 382.000 4.280 ;
        RECT 382.840 4.000 385.220 4.280 ;
        RECT 386.060 4.000 388.440 4.280 ;
        RECT 389.280 4.000 391.200 4.280 ;
        RECT 392.040 4.000 394.420 4.280 ;
        RECT 395.260 4.000 397.640 4.280 ;
        RECT 398.480 4.000 400.400 4.280 ;
        RECT 401.240 4.000 403.620 4.280 ;
        RECT 404.460 4.000 406.840 4.280 ;
        RECT 407.680 4.000 409.600 4.280 ;
        RECT 410.440 4.000 412.820 4.280 ;
        RECT 413.660 4.000 416.040 4.280 ;
        RECT 416.880 4.000 418.800 4.280 ;
        RECT 419.640 4.000 422.020 4.280 ;
        RECT 422.860 4.000 425.240 4.280 ;
        RECT 426.080 4.000 428.000 4.280 ;
        RECT 428.840 4.000 431.220 4.280 ;
        RECT 432.060 4.000 434.440 4.280 ;
        RECT 435.280 4.000 437.200 4.280 ;
        RECT 438.040 4.000 440.420 4.280 ;
        RECT 441.260 4.000 443.180 4.280 ;
        RECT 444.020 4.000 446.400 4.280 ;
        RECT 447.240 4.000 449.620 4.280 ;
        RECT 450.460 4.000 452.380 4.280 ;
        RECT 453.220 4.000 455.600 4.280 ;
        RECT 456.440 4.000 458.820 4.280 ;
        RECT 459.660 4.000 461.580 4.280 ;
        RECT 462.420 4.000 464.800 4.280 ;
        RECT 465.640 4.000 468.020 4.280 ;
        RECT 468.860 4.000 470.780 4.280 ;
        RECT 471.620 4.000 474.000 4.280 ;
        RECT 474.840 4.000 477.220 4.280 ;
        RECT 478.060 4.000 479.980 4.280 ;
        RECT 480.820 4.000 483.200 4.280 ;
        RECT 484.040 4.000 486.420 4.280 ;
        RECT 487.260 4.000 489.180 4.280 ;
        RECT 490.020 4.000 492.400 4.280 ;
        RECT 493.240 4.000 495.620 4.280 ;
        RECT 496.460 4.000 498.380 4.280 ;
        RECT 499.220 4.000 501.600 4.280 ;
        RECT 502.440 4.000 504.820 4.280 ;
        RECT 505.660 4.000 507.580 4.280 ;
        RECT 508.420 4.000 510.800 4.280 ;
        RECT 511.640 4.000 514.020 4.280 ;
        RECT 514.860 4.000 516.780 4.280 ;
        RECT 517.620 4.000 520.000 4.280 ;
        RECT 520.840 4.000 523.220 4.280 ;
        RECT 524.060 4.000 525.980 4.280 ;
        RECT 526.820 4.000 529.200 4.280 ;
        RECT 530.040 4.000 531.960 4.280 ;
        RECT 532.800 4.000 535.180 4.280 ;
        RECT 536.020 4.000 538.400 4.280 ;
        RECT 539.240 4.000 541.160 4.280 ;
        RECT 542.000 4.000 544.380 4.280 ;
        RECT 545.220 4.000 547.600 4.280 ;
        RECT 548.440 4.000 550.360 4.280 ;
        RECT 551.200 4.000 553.580 4.280 ;
        RECT 554.420 4.000 556.800 4.280 ;
        RECT 557.640 4.000 559.560 4.280 ;
        RECT 560.400 4.000 562.780 4.280 ;
        RECT 563.620 4.000 566.000 4.280 ;
        RECT 566.840 4.000 568.760 4.280 ;
        RECT 569.600 4.000 571.980 4.280 ;
        RECT 572.820 4.000 575.200 4.280 ;
        RECT 576.040 4.000 577.960 4.280 ;
        RECT 578.800 4.000 581.180 4.280 ;
        RECT 582.020 4.000 584.400 4.280 ;
        RECT 585.240 4.000 587.160 4.280 ;
        RECT 588.000 4.000 590.380 4.280 ;
        RECT 591.220 4.000 593.600 4.280 ;
        RECT 594.440 4.000 596.360 4.280 ;
        RECT 597.200 4.000 599.580 4.280 ;
        RECT 600.420 4.000 602.800 4.280 ;
        RECT 603.640 4.000 605.560 4.280 ;
        RECT 606.400 4.000 608.780 4.280 ;
        RECT 609.620 4.000 612.000 4.280 ;
        RECT 612.840 4.000 614.760 4.280 ;
        RECT 615.600 4.000 617.980 4.280 ;
        RECT 618.820 4.000 620.740 4.280 ;
        RECT 621.580 4.000 623.960 4.280 ;
        RECT 624.800 4.000 627.180 4.280 ;
        RECT 628.020 4.000 629.940 4.280 ;
        RECT 630.780 4.000 633.160 4.280 ;
        RECT 634.000 4.000 636.380 4.280 ;
        RECT 637.220 4.000 639.140 4.280 ;
        RECT 639.980 4.000 642.360 4.280 ;
        RECT 643.200 4.000 645.580 4.280 ;
        RECT 646.420 4.000 648.340 4.280 ;
        RECT 649.180 4.000 651.560 4.280 ;
        RECT 652.400 4.000 654.780 4.280 ;
        RECT 655.620 4.000 657.540 4.280 ;
        RECT 658.380 4.000 660.760 4.280 ;
        RECT 661.600 4.000 663.980 4.280 ;
        RECT 664.820 4.000 666.740 4.280 ;
        RECT 667.580 4.000 669.960 4.280 ;
        RECT 670.800 4.000 673.180 4.280 ;
        RECT 674.020 4.000 675.940 4.280 ;
        RECT 676.780 4.000 679.160 4.280 ;
        RECT 680.000 4.000 682.380 4.280 ;
        RECT 683.220 4.000 685.140 4.280 ;
        RECT 685.980 4.000 688.360 4.280 ;
        RECT 689.200 4.000 691.580 4.280 ;
        RECT 692.420 4.000 694.340 4.280 ;
        RECT 695.180 4.000 697.560 4.280 ;
        RECT 698.400 4.000 700.780 4.280 ;
        RECT 701.620 4.000 703.540 4.280 ;
        RECT 704.380 4.000 706.760 4.280 ;
        RECT 707.600 4.000 709.520 4.280 ;
        RECT 710.360 4.000 712.740 4.280 ;
        RECT 713.580 4.000 715.960 4.280 ;
        RECT 716.800 4.000 718.720 4.280 ;
        RECT 719.560 4.000 721.940 4.280 ;
        RECT 722.780 4.000 725.160 4.280 ;
        RECT 726.000 4.000 727.920 4.280 ;
        RECT 728.760 4.000 731.140 4.280 ;
        RECT 731.980 4.000 734.360 4.280 ;
        RECT 735.200 4.000 737.120 4.280 ;
        RECT 737.960 4.000 740.340 4.280 ;
        RECT 741.180 4.000 743.560 4.280 ;
        RECT 744.400 4.000 746.320 4.280 ;
        RECT 747.160 4.000 749.540 4.280 ;
        RECT 750.380 4.000 752.760 4.280 ;
        RECT 753.600 4.000 755.520 4.280 ;
        RECT 756.360 4.000 758.740 4.280 ;
        RECT 759.580 4.000 761.960 4.280 ;
        RECT 762.800 4.000 764.720 4.280 ;
        RECT 765.560 4.000 767.940 4.280 ;
        RECT 768.780 4.000 771.160 4.280 ;
        RECT 772.000 4.000 773.920 4.280 ;
        RECT 774.760 4.000 777.140 4.280 ;
        RECT 777.980 4.000 780.360 4.280 ;
        RECT 781.200 4.000 783.120 4.280 ;
        RECT 783.960 4.000 786.340 4.280 ;
        RECT 787.180 4.000 789.560 4.280 ;
        RECT 790.400 4.000 792.320 4.280 ;
        RECT 793.160 4.000 795.540 4.280 ;
        RECT 796.380 4.000 798.300 4.280 ;
        RECT 799.140 4.000 801.520 4.280 ;
        RECT 802.360 4.000 804.740 4.280 ;
        RECT 805.580 4.000 807.500 4.280 ;
        RECT 808.340 4.000 810.720 4.280 ;
        RECT 811.560 4.000 813.940 4.280 ;
        RECT 814.780 4.000 816.700 4.280 ;
        RECT 817.540 4.000 819.920 4.280 ;
        RECT 820.760 4.000 823.140 4.280 ;
        RECT 823.980 4.000 825.900 4.280 ;
        RECT 826.740 4.000 829.120 4.280 ;
        RECT 829.960 4.000 832.340 4.280 ;
        RECT 833.180 4.000 835.100 4.280 ;
        RECT 835.940 4.000 838.320 4.280 ;
        RECT 839.160 4.000 841.540 4.280 ;
        RECT 842.380 4.000 844.300 4.280 ;
        RECT 845.140 4.000 847.520 4.280 ;
        RECT 848.360 4.000 850.740 4.280 ;
        RECT 851.580 4.000 853.500 4.280 ;
        RECT 854.340 4.000 856.720 4.280 ;
        RECT 857.560 4.000 859.940 4.280 ;
        RECT 860.780 4.000 862.700 4.280 ;
        RECT 863.540 4.000 865.920 4.280 ;
        RECT 866.760 4.000 869.140 4.280 ;
        RECT 869.980 4.000 871.900 4.280 ;
        RECT 872.740 4.000 875.120 4.280 ;
        RECT 875.960 4.000 878.340 4.280 ;
        RECT 879.180 4.000 881.100 4.280 ;
        RECT 881.940 4.000 884.320 4.280 ;
        RECT 885.160 4.000 887.080 4.280 ;
        RECT 887.920 4.000 890.300 4.280 ;
        RECT 891.140 4.000 893.520 4.280 ;
        RECT 894.360 4.000 896.280 4.280 ;
        RECT 897.120 4.000 899.500 4.280 ;
        RECT 900.340 4.000 902.720 4.280 ;
        RECT 903.560 4.000 905.480 4.280 ;
        RECT 906.320 4.000 908.700 4.280 ;
        RECT 909.540 4.000 911.920 4.280 ;
        RECT 912.760 4.000 914.680 4.280 ;
        RECT 915.520 4.000 917.900 4.280 ;
        RECT 918.740 4.000 921.120 4.280 ;
        RECT 921.960 4.000 923.880 4.280 ;
        RECT 924.720 4.000 927.100 4.280 ;
        RECT 927.940 4.000 930.320 4.280 ;
        RECT 931.160 4.000 933.080 4.280 ;
        RECT 933.920 4.000 936.300 4.280 ;
        RECT 937.140 4.000 939.520 4.280 ;
        RECT 940.360 4.000 942.280 4.280 ;
        RECT 943.120 4.000 945.500 4.280 ;
        RECT 946.340 4.000 948.720 4.280 ;
        RECT 949.560 4.000 951.480 4.280 ;
        RECT 952.320 4.000 954.700 4.280 ;
        RECT 955.540 4.000 957.920 4.280 ;
        RECT 958.760 4.000 960.680 4.280 ;
        RECT 961.520 4.000 963.900 4.280 ;
        RECT 964.740 4.000 967.120 4.280 ;
        RECT 967.960 4.000 969.880 4.280 ;
        RECT 970.720 4.000 973.100 4.280 ;
        RECT 973.940 4.000 975.860 4.280 ;
        RECT 976.700 4.000 979.080 4.280 ;
        RECT 979.920 4.000 982.300 4.280 ;
        RECT 983.140 4.000 985.060 4.280 ;
        RECT 985.900 4.000 988.280 4.280 ;
        RECT 989.120 4.000 991.500 4.280 ;
        RECT 992.340 4.000 994.260 4.280 ;
        RECT 995.100 4.000 997.480 4.280 ;
        RECT 998.320 4.000 1000.700 4.280 ;
        RECT 1001.540 4.000 1003.460 4.280 ;
        RECT 1004.300 4.000 1006.680 4.280 ;
        RECT 1007.520 4.000 1009.900 4.280 ;
        RECT 1010.740 4.000 1012.660 4.280 ;
        RECT 1013.500 4.000 1015.880 4.280 ;
        RECT 1016.720 4.000 1019.100 4.280 ;
        RECT 1019.940 4.000 1021.860 4.280 ;
        RECT 1022.700 4.000 1025.080 4.280 ;
        RECT 1025.920 4.000 1028.300 4.280 ;
        RECT 1029.140 4.000 1031.060 4.280 ;
        RECT 1031.900 4.000 1034.280 4.280 ;
        RECT 1035.120 4.000 1037.500 4.280 ;
        RECT 1038.340 4.000 1040.260 4.280 ;
        RECT 1041.100 4.000 1043.480 4.280 ;
        RECT 1044.320 4.000 1046.700 4.280 ;
        RECT 1047.540 4.000 1049.460 4.280 ;
        RECT 1050.300 4.000 1052.680 4.280 ;
        RECT 1053.520 4.000 1055.900 4.280 ;
        RECT 1056.740 4.000 1058.660 4.280 ;
        RECT 1059.500 4.000 1061.880 4.280 ;
        RECT 1062.720 4.000 1064.640 4.280 ;
        RECT 1065.480 4.000 1067.860 4.280 ;
        RECT 1068.700 4.000 1071.080 4.280 ;
        RECT 1071.920 4.000 1073.840 4.280 ;
        RECT 1074.680 4.000 1077.060 4.280 ;
        RECT 1077.900 4.000 1080.280 4.280 ;
        RECT 1081.120 4.000 1083.040 4.280 ;
        RECT 1083.880 4.000 1086.260 4.280 ;
        RECT 1087.100 4.000 1089.480 4.280 ;
        RECT 1090.320 4.000 1092.240 4.280 ;
        RECT 1093.080 4.000 1095.460 4.280 ;
        RECT 1096.300 4.000 1098.680 4.280 ;
        RECT 1099.520 4.000 1101.440 4.280 ;
        RECT 1102.280 4.000 1104.660 4.280 ;
        RECT 1105.500 4.000 1107.880 4.280 ;
        RECT 1108.720 4.000 1110.640 4.280 ;
        RECT 1111.480 4.000 1113.860 4.280 ;
        RECT 1114.700 4.000 1117.080 4.280 ;
        RECT 1117.920 4.000 1119.840 4.280 ;
        RECT 1120.680 4.000 1123.060 4.280 ;
        RECT 1123.900 4.000 1126.280 4.280 ;
        RECT 1127.120 4.000 1129.040 4.280 ;
        RECT 1129.880 4.000 1132.260 4.280 ;
        RECT 1133.100 4.000 1135.480 4.280 ;
        RECT 1136.320 4.000 1138.240 4.280 ;
        RECT 1139.080 4.000 1141.460 4.280 ;
        RECT 1142.300 4.000 1144.680 4.280 ;
        RECT 1145.520 4.000 1147.440 4.280 ;
        RECT 1148.280 4.000 1150.660 4.280 ;
        RECT 1151.500 4.000 1153.420 4.280 ;
        RECT 1154.260 4.000 1156.640 4.280 ;
        RECT 1157.480 4.000 1159.860 4.280 ;
        RECT 1160.700 4.000 1162.620 4.280 ;
        RECT 1163.460 4.000 1165.840 4.280 ;
        RECT 1166.680 4.000 1169.060 4.280 ;
        RECT 1169.900 4.000 1171.820 4.280 ;
        RECT 1172.660 4.000 1175.040 4.280 ;
        RECT 1175.880 4.000 1178.260 4.280 ;
        RECT 1179.100 4.000 1181.020 4.280 ;
        RECT 1181.860 4.000 1184.240 4.280 ;
        RECT 1185.080 4.000 1187.460 4.280 ;
        RECT 1188.300 4.000 1190.220 4.280 ;
        RECT 1191.060 4.000 1193.440 4.280 ;
        RECT 1194.280 4.000 1196.660 4.280 ;
        RECT 1197.500 4.000 1199.420 4.280 ;
        RECT 1200.260 4.000 1202.640 4.280 ;
        RECT 1203.480 4.000 1205.860 4.280 ;
        RECT 1206.700 4.000 1208.620 4.280 ;
        RECT 1209.460 4.000 1211.840 4.280 ;
        RECT 1212.680 4.000 1215.060 4.280 ;
        RECT 1215.900 4.000 1217.820 4.280 ;
        RECT 1218.660 4.000 1221.040 4.280 ;
        RECT 1221.880 4.000 1224.260 4.280 ;
        RECT 1225.100 4.000 1227.020 4.280 ;
        RECT 1227.860 4.000 1230.240 4.280 ;
        RECT 1231.080 4.000 1233.460 4.280 ;
        RECT 1234.300 4.000 1236.220 4.280 ;
        RECT 1237.060 4.000 1239.440 4.280 ;
        RECT 1240.280 4.000 1242.200 4.280 ;
        RECT 1243.040 4.000 1245.420 4.280 ;
        RECT 1246.260 4.000 1248.640 4.280 ;
        RECT 1249.480 4.000 1251.400 4.280 ;
        RECT 1252.240 4.000 1254.620 4.280 ;
        RECT 1255.460 4.000 1257.840 4.280 ;
        RECT 1258.680 4.000 1260.600 4.280 ;
        RECT 1261.440 4.000 1263.820 4.280 ;
        RECT 1264.660 4.000 1267.040 4.280 ;
        RECT 1267.880 4.000 1269.800 4.280 ;
        RECT 1270.640 4.000 1273.020 4.280 ;
        RECT 1273.860 4.000 1276.240 4.280 ;
        RECT 1277.080 4.000 1279.000 4.280 ;
        RECT 1279.840 4.000 1282.220 4.280 ;
        RECT 1283.060 4.000 1285.440 4.280 ;
        RECT 1286.280 4.000 1288.200 4.280 ;
        RECT 1289.040 4.000 1291.420 4.280 ;
        RECT 1292.260 4.000 1294.640 4.280 ;
        RECT 1295.480 4.000 1297.400 4.280 ;
        RECT 1298.240 4.000 1300.620 4.280 ;
        RECT 1301.460 4.000 1303.840 4.280 ;
        RECT 1304.680 4.000 1306.600 4.280 ;
        RECT 1307.440 4.000 1309.820 4.280 ;
        RECT 1310.660 4.000 1313.040 4.280 ;
        RECT 1313.880 4.000 1315.800 4.280 ;
        RECT 1316.640 4.000 1319.020 4.280 ;
        RECT 1319.860 4.000 1322.240 4.280 ;
        RECT 1323.080 4.000 1325.000 4.280 ;
        RECT 1325.840 4.000 1328.220 4.280 ;
        RECT 1329.060 4.000 1330.980 4.280 ;
        RECT 1331.820 4.000 1334.200 4.280 ;
        RECT 1335.040 4.000 1337.420 4.280 ;
        RECT 1338.260 4.000 1340.180 4.280 ;
        RECT 1341.020 4.000 1343.400 4.280 ;
        RECT 1344.240 4.000 1346.620 4.280 ;
        RECT 1347.460 4.000 1349.380 4.280 ;
        RECT 1350.220 4.000 1352.600 4.280 ;
        RECT 1353.440 4.000 1355.820 4.280 ;
        RECT 1356.660 4.000 1358.580 4.280 ;
        RECT 1359.420 4.000 1361.800 4.280 ;
        RECT 1362.640 4.000 1365.020 4.280 ;
        RECT 1365.860 4.000 1367.780 4.280 ;
        RECT 1368.620 4.000 1371.000 4.280 ;
        RECT 1371.840 4.000 1374.220 4.280 ;
        RECT 1375.060 4.000 1376.980 4.280 ;
        RECT 1377.820 4.000 1380.200 4.280 ;
        RECT 1381.040 4.000 1383.420 4.280 ;
        RECT 1384.260 4.000 1386.180 4.280 ;
        RECT 1387.020 4.000 1389.400 4.280 ;
        RECT 1390.240 4.000 1392.620 4.280 ;
        RECT 1393.460 4.000 1395.380 4.280 ;
        RECT 1396.220 4.000 1398.600 4.280 ;
        RECT 1399.440 4.000 1401.820 4.280 ;
        RECT 1402.660 4.000 1404.580 4.280 ;
        RECT 1405.420 4.000 1407.800 4.280 ;
        RECT 1408.640 4.000 1411.020 4.280 ;
        RECT 1411.860 4.000 1413.780 4.280 ;
        RECT 1414.620 4.000 1417.000 4.280 ;
        RECT 1417.840 4.000 1419.760 4.280 ;
        RECT 1420.600 4.000 1422.980 4.280 ;
        RECT 1423.820 4.000 1426.200 4.280 ;
        RECT 1427.040 4.000 1428.960 4.280 ;
        RECT 1429.800 4.000 1432.180 4.280 ;
        RECT 1433.020 4.000 1435.400 4.280 ;
        RECT 1436.240 4.000 1438.160 4.280 ;
        RECT 1439.000 4.000 1441.380 4.280 ;
        RECT 1442.220 4.000 1444.600 4.280 ;
        RECT 1445.440 4.000 1447.360 4.280 ;
        RECT 1448.200 4.000 1450.580 4.280 ;
        RECT 1451.420 4.000 1453.800 4.280 ;
        RECT 1454.640 4.000 1456.560 4.280 ;
        RECT 1457.400 4.000 1459.780 4.280 ;
        RECT 1460.620 4.000 1463.000 4.280 ;
        RECT 1463.840 4.000 1465.760 4.280 ;
        RECT 1466.600 4.000 1468.980 4.280 ;
        RECT 1469.820 4.000 1472.200 4.280 ;
        RECT 1473.040 4.000 1474.960 4.280 ;
        RECT 1475.800 4.000 1478.180 4.280 ;
        RECT 1479.020 4.000 1481.400 4.280 ;
        RECT 1482.240 4.000 1484.160 4.280 ;
        RECT 1485.000 4.000 1487.380 4.280 ;
        RECT 1488.220 4.000 1490.600 4.280 ;
        RECT 1491.440 4.000 1493.360 4.280 ;
        RECT 1494.200 4.000 1496.580 4.280 ;
      LAYER met3 ;
        RECT 2.755 4.255 1485.205 1488.005 ;
      LAYER met4 ;
        RECT 173.190 10.640 1480.390 1488.080 ;
  END
END user_proj_example
END LIBRARY

