VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 1097.880 BY 1100.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.700 1096.000 3.980 1100.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.040 1096.000 293.320 1100.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.020 1096.000 322.300 1100.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 351.000 1096.000 351.280 1100.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 379.520 1096.000 379.800 1100.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.500 1096.000 408.780 1100.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 437.480 1096.000 437.760 1100.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 466.460 1096.000 466.740 1100.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 495.440 1096.000 495.720 1100.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 524.420 1096.000 524.700 1100.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 553.400 1096.000 553.680 1100.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.220 1096.000 32.500 1100.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 582.380 1096.000 582.660 1100.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 611.360 1096.000 611.640 1100.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 640.340 1096.000 640.620 1100.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 669.320 1096.000 669.600 1100.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.300 1096.000 698.580 1100.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 727.280 1096.000 727.560 1100.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 755.800 1096.000 756.080 1100.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 784.780 1096.000 785.060 1100.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 813.760 1096.000 814.040 1100.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 842.740 1096.000 843.020 1100.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.200 1096.000 61.480 1100.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 871.720 1096.000 872.000 1100.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.700 1096.000 900.980 1100.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.680 1096.000 929.960 1100.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 958.660 1096.000 958.940 1100.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 987.640 1096.000 987.920 1100.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1016.620 1096.000 1016.900 1100.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1045.600 1096.000 1045.880 1100.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1074.580 1096.000 1074.860 1100.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.180 1096.000 90.460 1100.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.160 1096.000 119.440 1100.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.140 1096.000 148.420 1100.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 177.120 1096.000 177.400 1100.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.100 1096.000 206.380 1100.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 235.080 1096.000 235.360 1100.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.060 1096.000 264.340 1100.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.900 1096.000 13.180 1100.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 302.700 1096.000 302.980 1100.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 331.680 1096.000 331.960 1100.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 360.660 1096.000 360.940 1100.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 389.180 1096.000 389.460 1100.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 418.160 1096.000 418.440 1100.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 447.140 1096.000 447.420 1100.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 476.120 1096.000 476.400 1100.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 505.100 1096.000 505.380 1100.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 534.080 1096.000 534.360 1100.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 563.060 1096.000 563.340 1100.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.880 1096.000 42.160 1100.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 592.040 1096.000 592.320 1100.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 621.020 1096.000 621.300 1100.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 650.000 1096.000 650.280 1100.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 678.980 1096.000 679.260 1100.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 707.960 1096.000 708.240 1100.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 736.940 1096.000 737.220 1100.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 765.460 1096.000 765.740 1100.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 794.440 1096.000 794.720 1100.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 823.420 1096.000 823.700 1100.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.400 1096.000 852.680 1100.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.860 1096.000 71.140 1100.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 881.380 1096.000 881.660 1100.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 910.360 1096.000 910.640 1100.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 939.340 1096.000 939.620 1100.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 968.320 1096.000 968.600 1100.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 997.300 1096.000 997.580 1100.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1026.280 1096.000 1026.560 1100.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1055.260 1096.000 1055.540 1100.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1084.240 1096.000 1084.520 1100.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.840 1096.000 100.120 1100.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.820 1096.000 129.100 1100.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 157.800 1096.000 158.080 1100.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 186.780 1096.000 187.060 1100.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 215.760 1096.000 216.040 1100.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 244.740 1096.000 245.020 1100.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 273.720 1096.000 274.000 1100.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.560 1096.000 22.840 1100.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 312.360 1096.000 312.640 1100.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.340 1096.000 341.620 1100.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 370.320 1096.000 370.600 1100.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 398.840 1096.000 399.120 1100.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 427.820 1096.000 428.100 1100.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 456.800 1096.000 457.080 1100.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 485.780 1096.000 486.060 1100.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 514.760 1096.000 515.040 1100.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 543.740 1096.000 544.020 1100.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 572.720 1096.000 573.000 1100.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.540 1096.000 51.820 1100.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 601.700 1096.000 601.980 1100.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 630.680 1096.000 630.960 1100.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 659.660 1096.000 659.940 1100.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 688.640 1096.000 688.920 1100.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 717.620 1096.000 717.900 1100.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.140 1096.000 746.420 1100.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 775.120 1096.000 775.400 1100.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 804.100 1096.000 804.380 1100.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 833.080 1096.000 833.360 1100.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 862.060 1096.000 862.340 1100.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.520 1096.000 80.800 1100.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 891.040 1096.000 891.320 1100.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 920.020 1096.000 920.300 1100.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 949.000 1096.000 949.280 1100.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.980 1096.000 978.260 1100.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1006.960 1096.000 1007.240 1100.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1035.940 1096.000 1036.220 1100.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1064.920 1096.000 1065.200 1100.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1093.900 1096.000 1094.180 1100.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.500 1096.000 109.780 1100.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.480 1096.000 138.760 1100.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.460 1096.000 167.740 1100.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.440 1096.000 196.720 1100.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 225.420 1096.000 225.700 1100.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 254.400 1096.000 254.680 1100.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 283.380 1096.000 283.660 1100.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 237.840 0.000 238.120 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 911.280 0.000 911.560 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 917.720 0.000 918.000 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 924.620 0.000 924.900 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 931.520 0.000 931.800 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 937.960 0.000 938.240 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 944.860 0.000 945.140 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 951.300 0.000 951.580 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 958.200 0.000 958.480 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.100 0.000 965.380 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.540 0.000 971.820 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 305.000 0.000 305.280 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 978.440 0.000 978.720 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 985.340 0.000 985.620 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 991.780 0.000 992.060 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 998.680 0.000 998.960 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1005.580 0.000 1005.860 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1012.020 0.000 1012.300 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1018.920 0.000 1019.200 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.360 0.000 1025.640 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.260 0.000 1032.540 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1039.160 0.000 1039.440 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.900 0.000 312.180 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1045.600 0.000 1045.880 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1052.500 0.000 1052.780 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1059.400 0.000 1059.680 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1065.840 0.000 1066.120 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1072.740 0.000 1073.020 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.640 0.000 1079.920 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1086.080 0.000 1086.360 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1092.980 0.000 1093.260 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 318.340 0.000 318.620 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 325.240 0.000 325.520 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 332.140 0.000 332.420 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 338.580 0.000 338.860 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.480 0.000 345.760 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 352.380 0.000 352.660 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 358.820 0.000 359.100 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.720 0.000 366.000 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.280 0.000 244.560 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.620 0.000 372.900 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 379.060 0.000 379.340 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 385.960 0.000 386.240 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.400 0.000 392.680 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 399.300 0.000 399.580 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 406.200 0.000 406.480 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 412.640 0.000 412.920 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.540 0.000 419.820 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.440 0.000 426.720 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.880 0.000 433.160 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 251.180 0.000 251.460 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 439.780 0.000 440.060 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 446.680 0.000 446.960 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 453.120 0.000 453.400 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.020 0.000 460.300 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 466.460 0.000 466.740 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 473.360 0.000 473.640 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 480.260 0.000 480.540 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 486.700 0.000 486.980 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 493.600 0.000 493.880 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 500.500 0.000 500.780 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.080 0.000 258.360 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 506.940 0.000 507.220 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.840 0.000 514.120 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 520.740 0.000 521.020 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.180 0.000 527.460 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 534.080 0.000 534.360 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 540.520 0.000 540.800 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 547.420 0.000 547.700 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 554.320 0.000 554.600 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 560.760 0.000 561.040 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.660 0.000 567.940 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.520 0.000 264.800 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 574.560 0.000 574.840 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 581.000 0.000 581.280 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.900 0.000 588.180 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 594.800 0.000 595.080 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 601.240 0.000 601.520 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 608.140 0.000 608.420 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 615.040 0.000 615.320 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 621.480 0.000 621.760 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 628.380 0.000 628.660 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 634.820 0.000 635.100 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.420 0.000 271.700 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 641.720 0.000 642.000 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 648.620 0.000 648.900 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 655.060 0.000 655.340 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 661.960 0.000 662.240 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.860 0.000 669.140 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 675.300 0.000 675.580 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 682.200 0.000 682.480 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 689.100 0.000 689.380 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 695.540 0.000 695.820 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 702.440 0.000 702.720 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 278.320 0.000 278.600 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 708.880 0.000 709.160 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 715.780 0.000 716.060 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.680 0.000 722.960 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 729.120 0.000 729.400 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 736.020 0.000 736.300 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 742.920 0.000 743.200 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 749.360 0.000 749.640 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 756.260 0.000 756.540 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 763.160 0.000 763.440 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.600 0.000 769.880 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 284.760 0.000 285.040 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 776.500 0.000 776.780 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 782.940 0.000 783.220 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 789.840 0.000 790.120 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 796.740 0.000 797.020 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 803.180 0.000 803.460 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 810.080 0.000 810.360 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 816.980 0.000 817.260 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.420 0.000 823.700 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 830.320 0.000 830.600 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 837.220 0.000 837.500 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 291.660 0.000 291.940 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 843.660 0.000 843.940 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 850.560 0.000 850.840 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 857.460 0.000 857.740 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 863.900 0.000 864.180 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 870.800 0.000 871.080 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 877.240 0.000 877.520 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 884.140 0.000 884.420 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 891.040 0.000 891.320 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 897.480 0.000 897.760 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 904.380 0.000 904.660 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 298.100 0.000 298.380 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 240.140 0.000 240.420 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 913.120 0.000 913.400 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 920.020 0.000 920.300 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 926.920 0.000 927.200 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 933.360 0.000 933.640 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 940.260 0.000 940.540 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 947.160 0.000 947.440 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 953.600 0.000 953.880 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 960.500 0.000 960.780 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 967.400 0.000 967.680 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 973.840 0.000 974.120 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 307.300 0.000 307.580 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 980.740 0.000 981.020 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 987.640 0.000 987.920 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 994.080 0.000 994.360 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1000.980 0.000 1001.260 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1007.420 0.000 1007.700 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1014.320 0.000 1014.600 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1021.220 0.000 1021.500 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1027.660 0.000 1027.940 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1034.560 0.000 1034.840 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1041.460 0.000 1041.740 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 314.200 0.000 314.480 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1047.900 0.000 1048.180 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1054.800 0.000 1055.080 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1061.700 0.000 1061.980 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1068.140 0.000 1068.420 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1075.040 0.000 1075.320 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1081.480 0.000 1081.760 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1088.380 0.000 1088.660 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1095.280 0.000 1095.560 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 320.640 0.000 320.920 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 327.540 0.000 327.820 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 334.440 0.000 334.720 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 340.880 0.000 341.160 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.780 0.000 348.060 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.220 0.000 354.500 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 361.120 0.000 361.400 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.020 0.000 368.300 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 246.580 0.000 246.860 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 374.460 0.000 374.740 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 381.360 0.000 381.640 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.260 0.000 388.540 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 394.700 0.000 394.980 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 401.600 0.000 401.880 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 408.500 0.000 408.780 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 414.940 0.000 415.220 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 421.840 0.000 422.120 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 428.740 0.000 429.020 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 435.180 0.000 435.460 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 253.480 0.000 253.760 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 442.080 0.000 442.360 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.520 0.000 448.800 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 455.420 0.000 455.700 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 462.320 0.000 462.600 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 468.760 0.000 469.040 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 475.660 0.000 475.940 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 482.560 0.000 482.840 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.000 0.000 489.280 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 495.900 0.000 496.180 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.800 0.000 503.080 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 260.380 0.000 260.660 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 509.240 0.000 509.520 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 516.140 0.000 516.420 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 522.580 0.000 522.860 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 529.480 0.000 529.760 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 536.380 0.000 536.660 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 542.820 0.000 543.100 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 549.720 0.000 550.000 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 556.620 0.000 556.900 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 563.060 0.000 563.340 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 569.960 0.000 570.240 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 266.820 0.000 267.100 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 576.860 0.000 577.140 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 583.300 0.000 583.580 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 590.200 0.000 590.480 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 596.640 0.000 596.920 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 603.540 0.000 603.820 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 610.440 0.000 610.720 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 616.880 0.000 617.160 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 623.780 0.000 624.060 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 630.680 0.000 630.960 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 637.120 0.000 637.400 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 273.720 0.000 274.000 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 644.020 0.000 644.300 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 650.920 0.000 651.200 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 657.360 0.000 657.640 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 664.260 0.000 664.540 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 670.700 0.000 670.980 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 677.600 0.000 677.880 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 684.500 0.000 684.780 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 690.940 0.000 691.220 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 697.840 0.000 698.120 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 704.740 0.000 705.020 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 280.160 0.000 280.440 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 711.180 0.000 711.460 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 718.080 0.000 718.360 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 724.980 0.000 725.260 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 731.420 0.000 731.700 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 738.320 0.000 738.600 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 745.220 0.000 745.500 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 751.660 0.000 751.940 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 758.560 0.000 758.840 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 765.000 0.000 765.280 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 771.900 0.000 772.180 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.060 0.000 287.340 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 778.800 0.000 779.080 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 785.240 0.000 785.520 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 792.140 0.000 792.420 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.040 0.000 799.320 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 805.480 0.000 805.760 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 812.380 0.000 812.660 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 819.280 0.000 819.560 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 825.720 0.000 826.000 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 832.620 0.000 832.900 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 839.060 0.000 839.340 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 293.960 0.000 294.240 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 845.960 0.000 846.240 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.860 0.000 853.140 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 859.300 0.000 859.580 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 866.200 0.000 866.480 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 873.100 0.000 873.380 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 879.540 0.000 879.820 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 886.440 0.000 886.720 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 893.340 0.000 893.620 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 899.780 0.000 900.060 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.680 0.000 906.960 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 300.400 0.000 300.680 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 241.980 0.000 242.260 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 915.420 0.000 915.700 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 922.320 0.000 922.600 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.220 0.000 929.500 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 935.660 0.000 935.940 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 942.560 0.000 942.840 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.460 0.000 949.740 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 955.900 0.000 956.180 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 962.800 0.000 963.080 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 969.240 0.000 969.520 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 976.140 0.000 976.420 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 309.600 0.000 309.880 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.040 0.000 983.320 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.480 0.000 989.760 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 996.380 0.000 996.660 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1003.280 0.000 1003.560 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1009.720 0.000 1010.000 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1016.620 0.000 1016.900 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1023.520 0.000 1023.800 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1029.960 0.000 1030.240 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1036.860 0.000 1037.140 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.760 0.000 1044.040 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.500 0.000 316.780 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1050.200 0.000 1050.480 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1057.100 0.000 1057.380 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.540 0.000 1063.820 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1070.440 0.000 1070.720 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1077.340 0.000 1077.620 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.780 0.000 1084.060 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.680 0.000 1090.960 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1097.580 0.000 1097.860 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.940 0.000 323.220 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.840 0.000 330.120 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 336.280 0.000 336.560 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 343.180 0.000 343.460 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 350.080 0.000 350.360 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 356.520 0.000 356.800 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 363.420 0.000 363.700 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 370.320 0.000 370.600 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 248.880 0.000 249.160 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 376.760 0.000 377.040 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.660 0.000 383.940 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.560 0.000 390.840 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 397.000 0.000 397.280 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.900 0.000 404.180 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 410.340 0.000 410.620 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 417.240 0.000 417.520 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.140 0.000 424.420 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 430.580 0.000 430.860 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 437.480 0.000 437.760 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 255.780 0.000 256.060 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 444.380 0.000 444.660 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 450.820 0.000 451.100 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 457.720 0.000 458.000 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 464.620 0.000 464.900 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.060 0.000 471.340 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.960 0.000 478.240 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 484.400 0.000 484.680 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 491.300 0.000 491.580 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 498.200 0.000 498.480 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 504.640 0.000 504.920 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 262.220 0.000 262.500 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 511.540 0.000 511.820 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 518.440 0.000 518.720 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 524.880 0.000 525.160 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.780 0.000 532.060 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 538.680 0.000 538.960 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 545.120 0.000 545.400 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 552.020 0.000 552.300 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 558.920 0.000 559.200 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 565.360 0.000 565.640 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 572.260 0.000 572.540 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.120 0.000 269.400 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 578.700 0.000 578.980 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.600 0.000 585.880 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 592.500 0.000 592.780 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 598.940 0.000 599.220 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 605.840 0.000 606.120 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 612.740 0.000 613.020 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 619.180 0.000 619.460 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 626.080 0.000 626.360 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.980 0.000 633.260 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 639.420 0.000 639.700 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 276.020 0.000 276.300 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 646.320 0.000 646.600 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 652.760 0.000 653.040 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 659.660 0.000 659.940 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 666.560 0.000 666.840 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 673.000 0.000 673.280 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 679.900 0.000 680.180 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.800 0.000 687.080 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 693.240 0.000 693.520 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 700.140 0.000 700.420 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 707.040 0.000 707.320 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.460 0.000 282.740 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 713.480 0.000 713.760 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 720.380 0.000 720.660 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 726.820 0.000 727.100 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 733.720 0.000 734.000 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.620 0.000 740.900 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 747.060 0.000 747.340 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 753.960 0.000 754.240 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 760.860 0.000 761.140 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 767.300 0.000 767.580 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 774.200 0.000 774.480 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 289.360 0.000 289.640 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 781.100 0.000 781.380 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.540 0.000 787.820 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 794.440 0.000 794.720 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 801.340 0.000 801.620 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 807.780 0.000 808.060 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 814.680 0.000 814.960 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 821.120 0.000 821.400 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 828.020 0.000 828.300 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 834.920 0.000 835.200 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 841.360 0.000 841.640 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 296.260 0.000 296.540 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 848.260 0.000 848.540 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 855.160 0.000 855.440 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 861.600 0.000 861.880 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 868.500 0.000 868.780 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 875.400 0.000 875.680 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 881.840 0.000 882.120 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 888.740 0.000 889.020 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 895.180 0.000 895.460 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 902.080 0.000 902.360 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 908.980 0.000 909.260 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.700 0.000 302.980 4.000 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.860 0.000 2.140 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.160 0.000 4.440 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.360 0.000 13.640 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.720 0.000 90.000 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.160 0.000 96.440 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.060 0.000 103.340 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.960 0.000 110.240 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.400 0.000 116.680 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.300 0.000 123.580 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.200 0.000 130.480 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.640 0.000 136.920 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.540 0.000 143.820 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.980 0.000 150.260 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.100 0.000 22.380 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.880 0.000 157.160 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 163.780 0.000 164.060 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.220 0.000 170.500 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 177.120 0.000 177.400 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.020 0.000 184.300 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.460 0.000 190.740 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 197.360 0.000 197.640 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.260 0.000 204.540 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.700 0.000 210.980 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.600 0.000 217.880 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.300 0.000 31.580 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.040 0.000 224.320 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 230.940 0.000 231.220 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.040 0.000 40.320 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.240 0.000 49.520 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.680 0.000 55.960 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.580 0.000 62.860 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.480 0.000 69.760 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.920 0.000 76.200 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.820 0.000 83.100 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.460 0.000 6.740 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.660 0.000 15.940 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.020 0.000 92.300 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.460 0.000 98.740 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.360 0.000 105.640 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.800 0.000 112.080 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.700 0.000 118.980 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 125.600 0.000 125.880 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.040 0.000 132.320 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.940 0.000 139.220 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.840 0.000 146.120 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 152.280 0.000 152.560 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.400 0.000 24.680 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.180 0.000 159.460 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.080 0.000 166.360 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.520 0.000 172.800 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.420 0.000 179.700 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.320 0.000 186.600 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.760 0.000 193.040 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 199.660 0.000 199.940 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.100 0.000 206.380 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.000 0.000 213.280 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 219.900 0.000 220.180 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.600 0.000 33.880 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 226.340 0.000 226.620 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 233.240 0.000 233.520 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.340 0.000 42.620 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.540 0.000 51.820 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.980 0.000 58.260 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.880 0.000 65.160 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.780 0.000 72.060 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.220 0.000 78.500 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.120 0.000 85.400 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.960 0.000 18.240 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.860 0.000 94.140 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.760 0.000 101.040 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.660 0.000 107.940 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.100 0.000 114.380 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.000 0.000 121.280 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.900 0.000 128.180 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.340 0.000 134.620 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 141.240 0.000 141.520 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 148.140 0.000 148.420 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 154.580 0.000 154.860 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.700 0.000 26.980 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 161.480 0.000 161.760 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.920 0.000 168.200 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.820 0.000 175.100 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.720 0.000 182.000 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 188.160 0.000 188.440 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 195.060 0.000 195.340 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 201.960 0.000 202.240 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.400 0.000 208.680 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 215.300 0.000 215.580 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.200 0.000 222.480 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.900 0.000 36.180 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 228.640 0.000 228.920 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 235.540 0.000 235.820 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.640 0.000 44.920 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.840 0.000 54.120 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.280 0.000 60.560 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.180 0.000 67.460 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.080 0.000 74.360 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.520 0.000 80.800 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.420 0.000 87.700 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.800 0.000 20.080 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.000 0.000 29.280 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.740 0.000 38.020 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.940 0.000 47.220 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.760 0.000 9.040 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.060 0.000 11.340 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.050 10.640 21.650 1088.240 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.850 10.640 98.450 1088.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.530 7.225 1093.350 1088.085 ;
      LAYER met1 ;
        RECT 0.000 5.480 1097.880 1095.780 ;
      LAYER met2 ;
        RECT 0.030 1095.720 3.420 1096.000 ;
        RECT 4.260 1095.720 12.620 1096.000 ;
        RECT 13.460 1095.720 22.280 1096.000 ;
        RECT 23.120 1095.720 31.940 1096.000 ;
        RECT 32.780 1095.720 41.600 1096.000 ;
        RECT 42.440 1095.720 51.260 1096.000 ;
        RECT 52.100 1095.720 60.920 1096.000 ;
        RECT 61.760 1095.720 70.580 1096.000 ;
        RECT 71.420 1095.720 80.240 1096.000 ;
        RECT 81.080 1095.720 89.900 1096.000 ;
        RECT 90.740 1095.720 99.560 1096.000 ;
        RECT 100.400 1095.720 109.220 1096.000 ;
        RECT 110.060 1095.720 118.880 1096.000 ;
        RECT 119.720 1095.720 128.540 1096.000 ;
        RECT 129.380 1095.720 138.200 1096.000 ;
        RECT 139.040 1095.720 147.860 1096.000 ;
        RECT 148.700 1095.720 157.520 1096.000 ;
        RECT 158.360 1095.720 167.180 1096.000 ;
        RECT 168.020 1095.720 176.840 1096.000 ;
        RECT 177.680 1095.720 186.500 1096.000 ;
        RECT 187.340 1095.720 196.160 1096.000 ;
        RECT 197.000 1095.720 205.820 1096.000 ;
        RECT 206.660 1095.720 215.480 1096.000 ;
        RECT 216.320 1095.720 225.140 1096.000 ;
        RECT 225.980 1095.720 234.800 1096.000 ;
        RECT 235.640 1095.720 244.460 1096.000 ;
        RECT 245.300 1095.720 254.120 1096.000 ;
        RECT 254.960 1095.720 263.780 1096.000 ;
        RECT 264.620 1095.720 273.440 1096.000 ;
        RECT 274.280 1095.720 283.100 1096.000 ;
        RECT 283.940 1095.720 292.760 1096.000 ;
        RECT 293.600 1095.720 302.420 1096.000 ;
        RECT 303.260 1095.720 312.080 1096.000 ;
        RECT 312.920 1095.720 321.740 1096.000 ;
        RECT 322.580 1095.720 331.400 1096.000 ;
        RECT 332.240 1095.720 341.060 1096.000 ;
        RECT 341.900 1095.720 350.720 1096.000 ;
        RECT 351.560 1095.720 360.380 1096.000 ;
        RECT 361.220 1095.720 370.040 1096.000 ;
        RECT 370.880 1095.720 379.240 1096.000 ;
        RECT 380.080 1095.720 388.900 1096.000 ;
        RECT 389.740 1095.720 398.560 1096.000 ;
        RECT 399.400 1095.720 408.220 1096.000 ;
        RECT 409.060 1095.720 417.880 1096.000 ;
        RECT 418.720 1095.720 427.540 1096.000 ;
        RECT 428.380 1095.720 437.200 1096.000 ;
        RECT 438.040 1095.720 446.860 1096.000 ;
        RECT 447.700 1095.720 456.520 1096.000 ;
        RECT 457.360 1095.720 466.180 1096.000 ;
        RECT 467.020 1095.720 475.840 1096.000 ;
        RECT 476.680 1095.720 485.500 1096.000 ;
        RECT 486.340 1095.720 495.160 1096.000 ;
        RECT 496.000 1095.720 504.820 1096.000 ;
        RECT 505.660 1095.720 514.480 1096.000 ;
        RECT 515.320 1095.720 524.140 1096.000 ;
        RECT 524.980 1095.720 533.800 1096.000 ;
        RECT 534.640 1095.720 543.460 1096.000 ;
        RECT 544.300 1095.720 553.120 1096.000 ;
        RECT 553.960 1095.720 562.780 1096.000 ;
        RECT 563.620 1095.720 572.440 1096.000 ;
        RECT 573.280 1095.720 582.100 1096.000 ;
        RECT 582.940 1095.720 591.760 1096.000 ;
        RECT 592.600 1095.720 601.420 1096.000 ;
        RECT 602.260 1095.720 611.080 1096.000 ;
        RECT 611.920 1095.720 620.740 1096.000 ;
        RECT 621.580 1095.720 630.400 1096.000 ;
        RECT 631.240 1095.720 640.060 1096.000 ;
        RECT 640.900 1095.720 649.720 1096.000 ;
        RECT 650.560 1095.720 659.380 1096.000 ;
        RECT 660.220 1095.720 669.040 1096.000 ;
        RECT 669.880 1095.720 678.700 1096.000 ;
        RECT 679.540 1095.720 688.360 1096.000 ;
        RECT 689.200 1095.720 698.020 1096.000 ;
        RECT 698.860 1095.720 707.680 1096.000 ;
        RECT 708.520 1095.720 717.340 1096.000 ;
        RECT 718.180 1095.720 727.000 1096.000 ;
        RECT 727.840 1095.720 736.660 1096.000 ;
        RECT 737.500 1095.720 745.860 1096.000 ;
        RECT 746.700 1095.720 755.520 1096.000 ;
        RECT 756.360 1095.720 765.180 1096.000 ;
        RECT 766.020 1095.720 774.840 1096.000 ;
        RECT 775.680 1095.720 784.500 1096.000 ;
        RECT 785.340 1095.720 794.160 1096.000 ;
        RECT 795.000 1095.720 803.820 1096.000 ;
        RECT 804.660 1095.720 813.480 1096.000 ;
        RECT 814.320 1095.720 823.140 1096.000 ;
        RECT 823.980 1095.720 832.800 1096.000 ;
        RECT 833.640 1095.720 842.460 1096.000 ;
        RECT 843.300 1095.720 852.120 1096.000 ;
        RECT 852.960 1095.720 861.780 1096.000 ;
        RECT 862.620 1095.720 871.440 1096.000 ;
        RECT 872.280 1095.720 881.100 1096.000 ;
        RECT 881.940 1095.720 890.760 1096.000 ;
        RECT 891.600 1095.720 900.420 1096.000 ;
        RECT 901.260 1095.720 910.080 1096.000 ;
        RECT 910.920 1095.720 919.740 1096.000 ;
        RECT 920.580 1095.720 929.400 1096.000 ;
        RECT 930.240 1095.720 939.060 1096.000 ;
        RECT 939.900 1095.720 948.720 1096.000 ;
        RECT 949.560 1095.720 958.380 1096.000 ;
        RECT 959.220 1095.720 968.040 1096.000 ;
        RECT 968.880 1095.720 977.700 1096.000 ;
        RECT 978.540 1095.720 987.360 1096.000 ;
        RECT 988.200 1095.720 997.020 1096.000 ;
        RECT 997.860 1095.720 1006.680 1096.000 ;
        RECT 1007.520 1095.720 1016.340 1096.000 ;
        RECT 1017.180 1095.720 1026.000 1096.000 ;
        RECT 1026.840 1095.720 1035.660 1096.000 ;
        RECT 1036.500 1095.720 1045.320 1096.000 ;
        RECT 1046.160 1095.720 1054.980 1096.000 ;
        RECT 1055.820 1095.720 1064.640 1096.000 ;
        RECT 1065.480 1095.720 1074.300 1096.000 ;
        RECT 1075.140 1095.720 1083.960 1096.000 ;
        RECT 1084.800 1095.720 1093.620 1096.000 ;
        RECT 1094.460 1095.720 1097.850 1096.000 ;
        RECT 0.030 4.280 1097.850 1095.720 ;
        RECT 0.580 4.000 1.580 4.280 ;
        RECT 2.420 4.000 3.880 4.280 ;
        RECT 4.720 4.000 6.180 4.280 ;
        RECT 7.020 4.000 8.480 4.280 ;
        RECT 9.320 4.000 10.780 4.280 ;
        RECT 11.620 4.000 13.080 4.280 ;
        RECT 13.920 4.000 15.380 4.280 ;
        RECT 16.220 4.000 17.680 4.280 ;
        RECT 18.520 4.000 19.520 4.280 ;
        RECT 20.360 4.000 21.820 4.280 ;
        RECT 22.660 4.000 24.120 4.280 ;
        RECT 24.960 4.000 26.420 4.280 ;
        RECT 27.260 4.000 28.720 4.280 ;
        RECT 29.560 4.000 31.020 4.280 ;
        RECT 31.860 4.000 33.320 4.280 ;
        RECT 34.160 4.000 35.620 4.280 ;
        RECT 36.460 4.000 37.460 4.280 ;
        RECT 38.300 4.000 39.760 4.280 ;
        RECT 40.600 4.000 42.060 4.280 ;
        RECT 42.900 4.000 44.360 4.280 ;
        RECT 45.200 4.000 46.660 4.280 ;
        RECT 47.500 4.000 48.960 4.280 ;
        RECT 49.800 4.000 51.260 4.280 ;
        RECT 52.100 4.000 53.560 4.280 ;
        RECT 54.400 4.000 55.400 4.280 ;
        RECT 56.240 4.000 57.700 4.280 ;
        RECT 58.540 4.000 60.000 4.280 ;
        RECT 60.840 4.000 62.300 4.280 ;
        RECT 63.140 4.000 64.600 4.280 ;
        RECT 65.440 4.000 66.900 4.280 ;
        RECT 67.740 4.000 69.200 4.280 ;
        RECT 70.040 4.000 71.500 4.280 ;
        RECT 72.340 4.000 73.800 4.280 ;
        RECT 74.640 4.000 75.640 4.280 ;
        RECT 76.480 4.000 77.940 4.280 ;
        RECT 78.780 4.000 80.240 4.280 ;
        RECT 81.080 4.000 82.540 4.280 ;
        RECT 83.380 4.000 84.840 4.280 ;
        RECT 85.680 4.000 87.140 4.280 ;
        RECT 87.980 4.000 89.440 4.280 ;
        RECT 90.280 4.000 91.740 4.280 ;
        RECT 92.580 4.000 93.580 4.280 ;
        RECT 94.420 4.000 95.880 4.280 ;
        RECT 96.720 4.000 98.180 4.280 ;
        RECT 99.020 4.000 100.480 4.280 ;
        RECT 101.320 4.000 102.780 4.280 ;
        RECT 103.620 4.000 105.080 4.280 ;
        RECT 105.920 4.000 107.380 4.280 ;
        RECT 108.220 4.000 109.680 4.280 ;
        RECT 110.520 4.000 111.520 4.280 ;
        RECT 112.360 4.000 113.820 4.280 ;
        RECT 114.660 4.000 116.120 4.280 ;
        RECT 116.960 4.000 118.420 4.280 ;
        RECT 119.260 4.000 120.720 4.280 ;
        RECT 121.560 4.000 123.020 4.280 ;
        RECT 123.860 4.000 125.320 4.280 ;
        RECT 126.160 4.000 127.620 4.280 ;
        RECT 128.460 4.000 129.920 4.280 ;
        RECT 130.760 4.000 131.760 4.280 ;
        RECT 132.600 4.000 134.060 4.280 ;
        RECT 134.900 4.000 136.360 4.280 ;
        RECT 137.200 4.000 138.660 4.280 ;
        RECT 139.500 4.000 140.960 4.280 ;
        RECT 141.800 4.000 143.260 4.280 ;
        RECT 144.100 4.000 145.560 4.280 ;
        RECT 146.400 4.000 147.860 4.280 ;
        RECT 148.700 4.000 149.700 4.280 ;
        RECT 150.540 4.000 152.000 4.280 ;
        RECT 152.840 4.000 154.300 4.280 ;
        RECT 155.140 4.000 156.600 4.280 ;
        RECT 157.440 4.000 158.900 4.280 ;
        RECT 159.740 4.000 161.200 4.280 ;
        RECT 162.040 4.000 163.500 4.280 ;
        RECT 164.340 4.000 165.800 4.280 ;
        RECT 166.640 4.000 167.640 4.280 ;
        RECT 168.480 4.000 169.940 4.280 ;
        RECT 170.780 4.000 172.240 4.280 ;
        RECT 173.080 4.000 174.540 4.280 ;
        RECT 175.380 4.000 176.840 4.280 ;
        RECT 177.680 4.000 179.140 4.280 ;
        RECT 179.980 4.000 181.440 4.280 ;
        RECT 182.280 4.000 183.740 4.280 ;
        RECT 184.580 4.000 186.040 4.280 ;
        RECT 186.880 4.000 187.880 4.280 ;
        RECT 188.720 4.000 190.180 4.280 ;
        RECT 191.020 4.000 192.480 4.280 ;
        RECT 193.320 4.000 194.780 4.280 ;
        RECT 195.620 4.000 197.080 4.280 ;
        RECT 197.920 4.000 199.380 4.280 ;
        RECT 200.220 4.000 201.680 4.280 ;
        RECT 202.520 4.000 203.980 4.280 ;
        RECT 204.820 4.000 205.820 4.280 ;
        RECT 206.660 4.000 208.120 4.280 ;
        RECT 208.960 4.000 210.420 4.280 ;
        RECT 211.260 4.000 212.720 4.280 ;
        RECT 213.560 4.000 215.020 4.280 ;
        RECT 215.860 4.000 217.320 4.280 ;
        RECT 218.160 4.000 219.620 4.280 ;
        RECT 220.460 4.000 221.920 4.280 ;
        RECT 222.760 4.000 223.760 4.280 ;
        RECT 224.600 4.000 226.060 4.280 ;
        RECT 226.900 4.000 228.360 4.280 ;
        RECT 229.200 4.000 230.660 4.280 ;
        RECT 231.500 4.000 232.960 4.280 ;
        RECT 233.800 4.000 235.260 4.280 ;
        RECT 236.100 4.000 237.560 4.280 ;
        RECT 238.400 4.000 239.860 4.280 ;
        RECT 240.700 4.000 241.700 4.280 ;
        RECT 242.540 4.000 244.000 4.280 ;
        RECT 244.840 4.000 246.300 4.280 ;
        RECT 247.140 4.000 248.600 4.280 ;
        RECT 249.440 4.000 250.900 4.280 ;
        RECT 251.740 4.000 253.200 4.280 ;
        RECT 254.040 4.000 255.500 4.280 ;
        RECT 256.340 4.000 257.800 4.280 ;
        RECT 258.640 4.000 260.100 4.280 ;
        RECT 260.940 4.000 261.940 4.280 ;
        RECT 262.780 4.000 264.240 4.280 ;
        RECT 265.080 4.000 266.540 4.280 ;
        RECT 267.380 4.000 268.840 4.280 ;
        RECT 269.680 4.000 271.140 4.280 ;
        RECT 271.980 4.000 273.440 4.280 ;
        RECT 274.280 4.000 275.740 4.280 ;
        RECT 276.580 4.000 278.040 4.280 ;
        RECT 278.880 4.000 279.880 4.280 ;
        RECT 280.720 4.000 282.180 4.280 ;
        RECT 283.020 4.000 284.480 4.280 ;
        RECT 285.320 4.000 286.780 4.280 ;
        RECT 287.620 4.000 289.080 4.280 ;
        RECT 289.920 4.000 291.380 4.280 ;
        RECT 292.220 4.000 293.680 4.280 ;
        RECT 294.520 4.000 295.980 4.280 ;
        RECT 296.820 4.000 297.820 4.280 ;
        RECT 298.660 4.000 300.120 4.280 ;
        RECT 300.960 4.000 302.420 4.280 ;
        RECT 303.260 4.000 304.720 4.280 ;
        RECT 305.560 4.000 307.020 4.280 ;
        RECT 307.860 4.000 309.320 4.280 ;
        RECT 310.160 4.000 311.620 4.280 ;
        RECT 312.460 4.000 313.920 4.280 ;
        RECT 314.760 4.000 316.220 4.280 ;
        RECT 317.060 4.000 318.060 4.280 ;
        RECT 318.900 4.000 320.360 4.280 ;
        RECT 321.200 4.000 322.660 4.280 ;
        RECT 323.500 4.000 324.960 4.280 ;
        RECT 325.800 4.000 327.260 4.280 ;
        RECT 328.100 4.000 329.560 4.280 ;
        RECT 330.400 4.000 331.860 4.280 ;
        RECT 332.700 4.000 334.160 4.280 ;
        RECT 335.000 4.000 336.000 4.280 ;
        RECT 336.840 4.000 338.300 4.280 ;
        RECT 339.140 4.000 340.600 4.280 ;
        RECT 341.440 4.000 342.900 4.280 ;
        RECT 343.740 4.000 345.200 4.280 ;
        RECT 346.040 4.000 347.500 4.280 ;
        RECT 348.340 4.000 349.800 4.280 ;
        RECT 350.640 4.000 352.100 4.280 ;
        RECT 352.940 4.000 353.940 4.280 ;
        RECT 354.780 4.000 356.240 4.280 ;
        RECT 357.080 4.000 358.540 4.280 ;
        RECT 359.380 4.000 360.840 4.280 ;
        RECT 361.680 4.000 363.140 4.280 ;
        RECT 363.980 4.000 365.440 4.280 ;
        RECT 366.280 4.000 367.740 4.280 ;
        RECT 368.580 4.000 370.040 4.280 ;
        RECT 370.880 4.000 372.340 4.280 ;
        RECT 373.180 4.000 374.180 4.280 ;
        RECT 375.020 4.000 376.480 4.280 ;
        RECT 377.320 4.000 378.780 4.280 ;
        RECT 379.620 4.000 381.080 4.280 ;
        RECT 381.920 4.000 383.380 4.280 ;
        RECT 384.220 4.000 385.680 4.280 ;
        RECT 386.520 4.000 387.980 4.280 ;
        RECT 388.820 4.000 390.280 4.280 ;
        RECT 391.120 4.000 392.120 4.280 ;
        RECT 392.960 4.000 394.420 4.280 ;
        RECT 395.260 4.000 396.720 4.280 ;
        RECT 397.560 4.000 399.020 4.280 ;
        RECT 399.860 4.000 401.320 4.280 ;
        RECT 402.160 4.000 403.620 4.280 ;
        RECT 404.460 4.000 405.920 4.280 ;
        RECT 406.760 4.000 408.220 4.280 ;
        RECT 409.060 4.000 410.060 4.280 ;
        RECT 410.900 4.000 412.360 4.280 ;
        RECT 413.200 4.000 414.660 4.280 ;
        RECT 415.500 4.000 416.960 4.280 ;
        RECT 417.800 4.000 419.260 4.280 ;
        RECT 420.100 4.000 421.560 4.280 ;
        RECT 422.400 4.000 423.860 4.280 ;
        RECT 424.700 4.000 426.160 4.280 ;
        RECT 427.000 4.000 428.460 4.280 ;
        RECT 429.300 4.000 430.300 4.280 ;
        RECT 431.140 4.000 432.600 4.280 ;
        RECT 433.440 4.000 434.900 4.280 ;
        RECT 435.740 4.000 437.200 4.280 ;
        RECT 438.040 4.000 439.500 4.280 ;
        RECT 440.340 4.000 441.800 4.280 ;
        RECT 442.640 4.000 444.100 4.280 ;
        RECT 444.940 4.000 446.400 4.280 ;
        RECT 447.240 4.000 448.240 4.280 ;
        RECT 449.080 4.000 450.540 4.280 ;
        RECT 451.380 4.000 452.840 4.280 ;
        RECT 453.680 4.000 455.140 4.280 ;
        RECT 455.980 4.000 457.440 4.280 ;
        RECT 458.280 4.000 459.740 4.280 ;
        RECT 460.580 4.000 462.040 4.280 ;
        RECT 462.880 4.000 464.340 4.280 ;
        RECT 465.180 4.000 466.180 4.280 ;
        RECT 467.020 4.000 468.480 4.280 ;
        RECT 469.320 4.000 470.780 4.280 ;
        RECT 471.620 4.000 473.080 4.280 ;
        RECT 473.920 4.000 475.380 4.280 ;
        RECT 476.220 4.000 477.680 4.280 ;
        RECT 478.520 4.000 479.980 4.280 ;
        RECT 480.820 4.000 482.280 4.280 ;
        RECT 483.120 4.000 484.120 4.280 ;
        RECT 484.960 4.000 486.420 4.280 ;
        RECT 487.260 4.000 488.720 4.280 ;
        RECT 489.560 4.000 491.020 4.280 ;
        RECT 491.860 4.000 493.320 4.280 ;
        RECT 494.160 4.000 495.620 4.280 ;
        RECT 496.460 4.000 497.920 4.280 ;
        RECT 498.760 4.000 500.220 4.280 ;
        RECT 501.060 4.000 502.520 4.280 ;
        RECT 503.360 4.000 504.360 4.280 ;
        RECT 505.200 4.000 506.660 4.280 ;
        RECT 507.500 4.000 508.960 4.280 ;
        RECT 509.800 4.000 511.260 4.280 ;
        RECT 512.100 4.000 513.560 4.280 ;
        RECT 514.400 4.000 515.860 4.280 ;
        RECT 516.700 4.000 518.160 4.280 ;
        RECT 519.000 4.000 520.460 4.280 ;
        RECT 521.300 4.000 522.300 4.280 ;
        RECT 523.140 4.000 524.600 4.280 ;
        RECT 525.440 4.000 526.900 4.280 ;
        RECT 527.740 4.000 529.200 4.280 ;
        RECT 530.040 4.000 531.500 4.280 ;
        RECT 532.340 4.000 533.800 4.280 ;
        RECT 534.640 4.000 536.100 4.280 ;
        RECT 536.940 4.000 538.400 4.280 ;
        RECT 539.240 4.000 540.240 4.280 ;
        RECT 541.080 4.000 542.540 4.280 ;
        RECT 543.380 4.000 544.840 4.280 ;
        RECT 545.680 4.000 547.140 4.280 ;
        RECT 547.980 4.000 549.440 4.280 ;
        RECT 550.280 4.000 551.740 4.280 ;
        RECT 552.580 4.000 554.040 4.280 ;
        RECT 554.880 4.000 556.340 4.280 ;
        RECT 557.180 4.000 558.640 4.280 ;
        RECT 559.480 4.000 560.480 4.280 ;
        RECT 561.320 4.000 562.780 4.280 ;
        RECT 563.620 4.000 565.080 4.280 ;
        RECT 565.920 4.000 567.380 4.280 ;
        RECT 568.220 4.000 569.680 4.280 ;
        RECT 570.520 4.000 571.980 4.280 ;
        RECT 572.820 4.000 574.280 4.280 ;
        RECT 575.120 4.000 576.580 4.280 ;
        RECT 577.420 4.000 578.420 4.280 ;
        RECT 579.260 4.000 580.720 4.280 ;
        RECT 581.560 4.000 583.020 4.280 ;
        RECT 583.860 4.000 585.320 4.280 ;
        RECT 586.160 4.000 587.620 4.280 ;
        RECT 588.460 4.000 589.920 4.280 ;
        RECT 590.760 4.000 592.220 4.280 ;
        RECT 593.060 4.000 594.520 4.280 ;
        RECT 595.360 4.000 596.360 4.280 ;
        RECT 597.200 4.000 598.660 4.280 ;
        RECT 599.500 4.000 600.960 4.280 ;
        RECT 601.800 4.000 603.260 4.280 ;
        RECT 604.100 4.000 605.560 4.280 ;
        RECT 606.400 4.000 607.860 4.280 ;
        RECT 608.700 4.000 610.160 4.280 ;
        RECT 611.000 4.000 612.460 4.280 ;
        RECT 613.300 4.000 614.760 4.280 ;
        RECT 615.600 4.000 616.600 4.280 ;
        RECT 617.440 4.000 618.900 4.280 ;
        RECT 619.740 4.000 621.200 4.280 ;
        RECT 622.040 4.000 623.500 4.280 ;
        RECT 624.340 4.000 625.800 4.280 ;
        RECT 626.640 4.000 628.100 4.280 ;
        RECT 628.940 4.000 630.400 4.280 ;
        RECT 631.240 4.000 632.700 4.280 ;
        RECT 633.540 4.000 634.540 4.280 ;
        RECT 635.380 4.000 636.840 4.280 ;
        RECT 637.680 4.000 639.140 4.280 ;
        RECT 639.980 4.000 641.440 4.280 ;
        RECT 642.280 4.000 643.740 4.280 ;
        RECT 644.580 4.000 646.040 4.280 ;
        RECT 646.880 4.000 648.340 4.280 ;
        RECT 649.180 4.000 650.640 4.280 ;
        RECT 651.480 4.000 652.480 4.280 ;
        RECT 653.320 4.000 654.780 4.280 ;
        RECT 655.620 4.000 657.080 4.280 ;
        RECT 657.920 4.000 659.380 4.280 ;
        RECT 660.220 4.000 661.680 4.280 ;
        RECT 662.520 4.000 663.980 4.280 ;
        RECT 664.820 4.000 666.280 4.280 ;
        RECT 667.120 4.000 668.580 4.280 ;
        RECT 669.420 4.000 670.420 4.280 ;
        RECT 671.260 4.000 672.720 4.280 ;
        RECT 673.560 4.000 675.020 4.280 ;
        RECT 675.860 4.000 677.320 4.280 ;
        RECT 678.160 4.000 679.620 4.280 ;
        RECT 680.460 4.000 681.920 4.280 ;
        RECT 682.760 4.000 684.220 4.280 ;
        RECT 685.060 4.000 686.520 4.280 ;
        RECT 687.360 4.000 688.820 4.280 ;
        RECT 689.660 4.000 690.660 4.280 ;
        RECT 691.500 4.000 692.960 4.280 ;
        RECT 693.800 4.000 695.260 4.280 ;
        RECT 696.100 4.000 697.560 4.280 ;
        RECT 698.400 4.000 699.860 4.280 ;
        RECT 700.700 4.000 702.160 4.280 ;
        RECT 703.000 4.000 704.460 4.280 ;
        RECT 705.300 4.000 706.760 4.280 ;
        RECT 707.600 4.000 708.600 4.280 ;
        RECT 709.440 4.000 710.900 4.280 ;
        RECT 711.740 4.000 713.200 4.280 ;
        RECT 714.040 4.000 715.500 4.280 ;
        RECT 716.340 4.000 717.800 4.280 ;
        RECT 718.640 4.000 720.100 4.280 ;
        RECT 720.940 4.000 722.400 4.280 ;
        RECT 723.240 4.000 724.700 4.280 ;
        RECT 725.540 4.000 726.540 4.280 ;
        RECT 727.380 4.000 728.840 4.280 ;
        RECT 729.680 4.000 731.140 4.280 ;
        RECT 731.980 4.000 733.440 4.280 ;
        RECT 734.280 4.000 735.740 4.280 ;
        RECT 736.580 4.000 738.040 4.280 ;
        RECT 738.880 4.000 740.340 4.280 ;
        RECT 741.180 4.000 742.640 4.280 ;
        RECT 743.480 4.000 744.940 4.280 ;
        RECT 745.780 4.000 746.780 4.280 ;
        RECT 747.620 4.000 749.080 4.280 ;
        RECT 749.920 4.000 751.380 4.280 ;
        RECT 752.220 4.000 753.680 4.280 ;
        RECT 754.520 4.000 755.980 4.280 ;
        RECT 756.820 4.000 758.280 4.280 ;
        RECT 759.120 4.000 760.580 4.280 ;
        RECT 761.420 4.000 762.880 4.280 ;
        RECT 763.720 4.000 764.720 4.280 ;
        RECT 765.560 4.000 767.020 4.280 ;
        RECT 767.860 4.000 769.320 4.280 ;
        RECT 770.160 4.000 771.620 4.280 ;
        RECT 772.460 4.000 773.920 4.280 ;
        RECT 774.760 4.000 776.220 4.280 ;
        RECT 777.060 4.000 778.520 4.280 ;
        RECT 779.360 4.000 780.820 4.280 ;
        RECT 781.660 4.000 782.660 4.280 ;
        RECT 783.500 4.000 784.960 4.280 ;
        RECT 785.800 4.000 787.260 4.280 ;
        RECT 788.100 4.000 789.560 4.280 ;
        RECT 790.400 4.000 791.860 4.280 ;
        RECT 792.700 4.000 794.160 4.280 ;
        RECT 795.000 4.000 796.460 4.280 ;
        RECT 797.300 4.000 798.760 4.280 ;
        RECT 799.600 4.000 801.060 4.280 ;
        RECT 801.900 4.000 802.900 4.280 ;
        RECT 803.740 4.000 805.200 4.280 ;
        RECT 806.040 4.000 807.500 4.280 ;
        RECT 808.340 4.000 809.800 4.280 ;
        RECT 810.640 4.000 812.100 4.280 ;
        RECT 812.940 4.000 814.400 4.280 ;
        RECT 815.240 4.000 816.700 4.280 ;
        RECT 817.540 4.000 819.000 4.280 ;
        RECT 819.840 4.000 820.840 4.280 ;
        RECT 821.680 4.000 823.140 4.280 ;
        RECT 823.980 4.000 825.440 4.280 ;
        RECT 826.280 4.000 827.740 4.280 ;
        RECT 828.580 4.000 830.040 4.280 ;
        RECT 830.880 4.000 832.340 4.280 ;
        RECT 833.180 4.000 834.640 4.280 ;
        RECT 835.480 4.000 836.940 4.280 ;
        RECT 837.780 4.000 838.780 4.280 ;
        RECT 839.620 4.000 841.080 4.280 ;
        RECT 841.920 4.000 843.380 4.280 ;
        RECT 844.220 4.000 845.680 4.280 ;
        RECT 846.520 4.000 847.980 4.280 ;
        RECT 848.820 4.000 850.280 4.280 ;
        RECT 851.120 4.000 852.580 4.280 ;
        RECT 853.420 4.000 854.880 4.280 ;
        RECT 855.720 4.000 857.180 4.280 ;
        RECT 858.020 4.000 859.020 4.280 ;
        RECT 859.860 4.000 861.320 4.280 ;
        RECT 862.160 4.000 863.620 4.280 ;
        RECT 864.460 4.000 865.920 4.280 ;
        RECT 866.760 4.000 868.220 4.280 ;
        RECT 869.060 4.000 870.520 4.280 ;
        RECT 871.360 4.000 872.820 4.280 ;
        RECT 873.660 4.000 875.120 4.280 ;
        RECT 875.960 4.000 876.960 4.280 ;
        RECT 877.800 4.000 879.260 4.280 ;
        RECT 880.100 4.000 881.560 4.280 ;
        RECT 882.400 4.000 883.860 4.280 ;
        RECT 884.700 4.000 886.160 4.280 ;
        RECT 887.000 4.000 888.460 4.280 ;
        RECT 889.300 4.000 890.760 4.280 ;
        RECT 891.600 4.000 893.060 4.280 ;
        RECT 893.900 4.000 894.900 4.280 ;
        RECT 895.740 4.000 897.200 4.280 ;
        RECT 898.040 4.000 899.500 4.280 ;
        RECT 900.340 4.000 901.800 4.280 ;
        RECT 902.640 4.000 904.100 4.280 ;
        RECT 904.940 4.000 906.400 4.280 ;
        RECT 907.240 4.000 908.700 4.280 ;
        RECT 909.540 4.000 911.000 4.280 ;
        RECT 911.840 4.000 912.840 4.280 ;
        RECT 913.680 4.000 915.140 4.280 ;
        RECT 915.980 4.000 917.440 4.280 ;
        RECT 918.280 4.000 919.740 4.280 ;
        RECT 920.580 4.000 922.040 4.280 ;
        RECT 922.880 4.000 924.340 4.280 ;
        RECT 925.180 4.000 926.640 4.280 ;
        RECT 927.480 4.000 928.940 4.280 ;
        RECT 929.780 4.000 931.240 4.280 ;
        RECT 932.080 4.000 933.080 4.280 ;
        RECT 933.920 4.000 935.380 4.280 ;
        RECT 936.220 4.000 937.680 4.280 ;
        RECT 938.520 4.000 939.980 4.280 ;
        RECT 940.820 4.000 942.280 4.280 ;
        RECT 943.120 4.000 944.580 4.280 ;
        RECT 945.420 4.000 946.880 4.280 ;
        RECT 947.720 4.000 949.180 4.280 ;
        RECT 950.020 4.000 951.020 4.280 ;
        RECT 951.860 4.000 953.320 4.280 ;
        RECT 954.160 4.000 955.620 4.280 ;
        RECT 956.460 4.000 957.920 4.280 ;
        RECT 958.760 4.000 960.220 4.280 ;
        RECT 961.060 4.000 962.520 4.280 ;
        RECT 963.360 4.000 964.820 4.280 ;
        RECT 965.660 4.000 967.120 4.280 ;
        RECT 967.960 4.000 968.960 4.280 ;
        RECT 969.800 4.000 971.260 4.280 ;
        RECT 972.100 4.000 973.560 4.280 ;
        RECT 974.400 4.000 975.860 4.280 ;
        RECT 976.700 4.000 978.160 4.280 ;
        RECT 979.000 4.000 980.460 4.280 ;
        RECT 981.300 4.000 982.760 4.280 ;
        RECT 983.600 4.000 985.060 4.280 ;
        RECT 985.900 4.000 987.360 4.280 ;
        RECT 988.200 4.000 989.200 4.280 ;
        RECT 990.040 4.000 991.500 4.280 ;
        RECT 992.340 4.000 993.800 4.280 ;
        RECT 994.640 4.000 996.100 4.280 ;
        RECT 996.940 4.000 998.400 4.280 ;
        RECT 999.240 4.000 1000.700 4.280 ;
        RECT 1001.540 4.000 1003.000 4.280 ;
        RECT 1003.840 4.000 1005.300 4.280 ;
        RECT 1006.140 4.000 1007.140 4.280 ;
        RECT 1007.980 4.000 1009.440 4.280 ;
        RECT 1010.280 4.000 1011.740 4.280 ;
        RECT 1012.580 4.000 1014.040 4.280 ;
        RECT 1014.880 4.000 1016.340 4.280 ;
        RECT 1017.180 4.000 1018.640 4.280 ;
        RECT 1019.480 4.000 1020.940 4.280 ;
        RECT 1021.780 4.000 1023.240 4.280 ;
        RECT 1024.080 4.000 1025.080 4.280 ;
        RECT 1025.920 4.000 1027.380 4.280 ;
        RECT 1028.220 4.000 1029.680 4.280 ;
        RECT 1030.520 4.000 1031.980 4.280 ;
        RECT 1032.820 4.000 1034.280 4.280 ;
        RECT 1035.120 4.000 1036.580 4.280 ;
        RECT 1037.420 4.000 1038.880 4.280 ;
        RECT 1039.720 4.000 1041.180 4.280 ;
        RECT 1042.020 4.000 1043.480 4.280 ;
        RECT 1044.320 4.000 1045.320 4.280 ;
        RECT 1046.160 4.000 1047.620 4.280 ;
        RECT 1048.460 4.000 1049.920 4.280 ;
        RECT 1050.760 4.000 1052.220 4.280 ;
        RECT 1053.060 4.000 1054.520 4.280 ;
        RECT 1055.360 4.000 1056.820 4.280 ;
        RECT 1057.660 4.000 1059.120 4.280 ;
        RECT 1059.960 4.000 1061.420 4.280 ;
        RECT 1062.260 4.000 1063.260 4.280 ;
        RECT 1064.100 4.000 1065.560 4.280 ;
        RECT 1066.400 4.000 1067.860 4.280 ;
        RECT 1068.700 4.000 1070.160 4.280 ;
        RECT 1071.000 4.000 1072.460 4.280 ;
        RECT 1073.300 4.000 1074.760 4.280 ;
        RECT 1075.600 4.000 1077.060 4.280 ;
        RECT 1077.900 4.000 1079.360 4.280 ;
        RECT 1080.200 4.000 1081.200 4.280 ;
        RECT 1082.040 4.000 1083.500 4.280 ;
        RECT 1084.340 4.000 1085.800 4.280 ;
        RECT 1086.640 4.000 1088.100 4.280 ;
        RECT 1088.940 4.000 1090.400 4.280 ;
        RECT 1091.240 4.000 1092.700 4.280 ;
        RECT 1093.540 4.000 1095.000 4.280 ;
        RECT 1095.840 4.000 1097.300 4.280 ;
      LAYER met3 ;
        RECT 1.835 10.715 1085.925 1088.165 ;
      LAYER met4 ;
        RECT 65.545 10.640 96.450 1088.240 ;
        RECT 98.850 10.640 1082.475 1088.240 ;
  END
END user_proj_example
END LIBRARY

