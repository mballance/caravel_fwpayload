VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN -0.005 0.000 ;
  SIZE 1197.705 BY 1200.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.170 1196.000 4.450 1200.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.730 1196.000 320.010 1200.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 351.470 1196.000 351.750 1200.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 382.750 1196.000 383.030 1200.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.490 1196.000 414.770 1200.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 446.230 1196.000 446.510 1200.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.510 1196.000 477.790 1200.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 509.250 1196.000 509.530 1200.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 540.990 1196.000 541.270 1200.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 572.270 1196.000 572.550 1200.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 604.010 1196.000 604.290 1200.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.450 1196.000 35.730 1200.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 635.750 1196.000 636.030 1200.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 667.030 1196.000 667.310 1200.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.770 1196.000 699.050 1200.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 730.510 1196.000 730.790 1200.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 761.790 1196.000 762.070 1200.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.530 1196.000 793.810 1200.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 825.270 1196.000 825.550 1200.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 856.550 1196.000 856.830 1200.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 888.290 1196.000 888.570 1200.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 920.030 1196.000 920.310 1200.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 67.190 1196.000 67.470 1200.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 951.310 1196.000 951.590 1200.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.050 1196.000 983.330 1200.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1014.790 1196.000 1015.070 1200.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1046.070 1196.000 1046.350 1200.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1077.810 1196.000 1078.090 1200.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1109.550 1196.000 1109.830 1200.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1140.830 1196.000 1141.110 1200.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1172.570 1196.000 1172.850 1200.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.470 1196.000 98.750 1200.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.210 1196.000 130.490 1200.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 161.950 1196.000 162.230 1200.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.230 1196.000 193.510 1200.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.970 1196.000 225.250 1200.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.710 1196.000 256.990 1200.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 287.990 1196.000 288.270 1200.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 14.290 1196.000 14.570 1200.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 330.310 1196.000 330.590 1200.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 362.050 1196.000 362.330 1200.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 393.330 1196.000 393.610 1200.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 425.070 1196.000 425.350 1200.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 456.810 1196.000 457.090 1200.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 488.090 1196.000 488.370 1200.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 519.830 1196.000 520.110 1200.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 551.570 1196.000 551.850 1200.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 582.850 1196.000 583.130 1200.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 614.590 1196.000 614.870 1200.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.030 1196.000 46.310 1200.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 646.330 1196.000 646.610 1200.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 677.610 1196.000 677.890 1200.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 709.350 1196.000 709.630 1200.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 741.090 1196.000 741.370 1200.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 772.370 1196.000 772.650 1200.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 804.110 1196.000 804.390 1200.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 835.390 1196.000 835.670 1200.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 867.130 1196.000 867.410 1200.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 898.870 1196.000 899.150 1200.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 930.150 1196.000 930.430 1200.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 77.770 1196.000 78.050 1200.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 961.890 1196.000 962.170 1200.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 993.630 1196.000 993.910 1200.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1024.910 1196.000 1025.190 1200.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1056.650 1196.000 1056.930 1200.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1088.390 1196.000 1088.670 1200.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1119.670 1196.000 1119.950 1200.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1151.410 1196.000 1151.690 1200.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1183.150 1196.000 1183.430 1200.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.050 1196.000 109.330 1200.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 140.790 1196.000 141.070 1200.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.530 1196.000 172.810 1200.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 203.810 1196.000 204.090 1200.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 235.550 1196.000 235.830 1200.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 267.290 1196.000 267.570 1200.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 298.570 1196.000 298.850 1200.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.870 1196.000 25.150 1200.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 340.890 1196.000 341.170 1200.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 372.630 1196.000 372.910 1200.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 403.910 1196.000 404.190 1200.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 435.650 1196.000 435.930 1200.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.930 1196.000 467.210 1200.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 498.670 1196.000 498.950 1200.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 530.410 1196.000 530.690 1200.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 561.690 1196.000 561.970 1200.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 593.430 1196.000 593.710 1200.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 625.170 1196.000 625.450 1200.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 56.610 1196.000 56.890 1200.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 656.450 1196.000 656.730 1200.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 688.190 1196.000 688.470 1200.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 719.930 1196.000 720.210 1200.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 751.210 1196.000 751.490 1200.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 782.950 1196.000 783.230 1200.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 814.690 1196.000 814.970 1200.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 845.970 1196.000 846.250 1200.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 877.710 1196.000 877.990 1200.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 909.450 1196.000 909.730 1200.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 940.730 1196.000 941.010 1200.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.350 1196.000 88.630 1200.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 972.470 1196.000 972.750 1200.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1004.210 1196.000 1004.490 1200.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1035.490 1196.000 1035.770 1200.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1067.230 1196.000 1067.510 1200.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1098.970 1196.000 1099.250 1200.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1130.250 1196.000 1130.530 1200.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1161.990 1196.000 1162.270 1200.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1193.730 1196.000 1194.010 1200.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.630 1196.000 119.910 1200.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 151.370 1196.000 151.650 1200.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.110 1196.000 183.390 1200.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 214.390 1196.000 214.670 1200.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 246.130 1196.000 246.410 1200.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 277.870 1196.000 278.150 1200.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 309.150 1196.000 309.430 1200.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 259.470 0.000 259.750 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 994.090 0.000 994.370 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.450 0.000 1001.730 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1008.810 0.000 1009.090 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1016.170 0.000 1016.450 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1023.530 0.000 1023.810 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1030.890 0.000 1031.170 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1038.250 0.000 1038.530 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1045.610 0.000 1045.890 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1052.970 0.000 1053.250 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1060.330 0.000 1060.610 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 333.070 0.000 333.350 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1067.690 0.000 1067.970 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1075.050 0.000 1075.330 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1082.410 0.000 1082.690 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1089.770 0.000 1090.050 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1097.130 0.000 1097.410 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1104.490 0.000 1104.770 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1111.850 0.000 1112.130 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1119.210 0.000 1119.490 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1126.570 0.000 1126.850 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1133.930 0.000 1134.210 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 340.430 0.000 340.710 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1141.290 0.000 1141.570 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1148.650 0.000 1148.930 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1156.010 0.000 1156.290 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1163.370 0.000 1163.650 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1170.730 0.000 1171.010 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1178.090 0.000 1178.370 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.450 0.000 1185.730 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1192.810 0.000 1193.090 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 347.790 0.000 348.070 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 355.150 0.000 355.430 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 362.510 0.000 362.790 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 369.410 0.000 369.690 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 376.770 0.000 377.050 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 384.130 0.000 384.410 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 391.490 0.000 391.770 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 398.850 0.000 399.130 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 266.830 0.000 267.110 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 406.210 0.000 406.490 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 413.570 0.000 413.850 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 420.930 0.000 421.210 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 428.290 0.000 428.570 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 435.650 0.000 435.930 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 443.010 0.000 443.290 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 450.370 0.000 450.650 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 457.730 0.000 458.010 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 465.090 0.000 465.370 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.450 0.000 472.730 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 274.190 0.000 274.470 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 479.810 0.000 480.090 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 487.170 0.000 487.450 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 494.530 0.000 494.810 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 501.890 0.000 502.170 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 509.250 0.000 509.530 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 516.610 0.000 516.890 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 523.970 0.000 524.250 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.330 0.000 531.610 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 538.690 0.000 538.970 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 546.050 0.000 546.330 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.550 0.000 281.830 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 553.410 0.000 553.690 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 560.770 0.000 561.050 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 568.130 0.000 568.410 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 575.490 0.000 575.770 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 582.850 0.000 583.130 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 590.210 0.000 590.490 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 597.570 0.000 597.850 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 604.930 0.000 605.210 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 612.290 0.000 612.570 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 619.650 0.000 619.930 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.910 0.000 289.190 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.010 0.000 627.290 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 634.370 0.000 634.650 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 641.730 0.000 642.010 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 648.630 0.000 648.910 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 655.990 0.000 656.270 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 663.350 0.000 663.630 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 670.710 0.000 670.990 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 678.070 0.000 678.350 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 685.430 0.000 685.710 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 692.790 0.000 693.070 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 296.270 0.000 296.550 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 700.150 0.000 700.430 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 707.510 0.000 707.790 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.870 0.000 715.150 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.230 0.000 722.510 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 729.590 0.000 729.870 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 736.950 0.000 737.230 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 744.310 0.000 744.590 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 751.670 0.000 751.950 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 759.030 0.000 759.310 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 766.390 0.000 766.670 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 303.630 0.000 303.910 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 773.750 0.000 774.030 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 781.110 0.000 781.390 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 788.470 0.000 788.750 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 795.830 0.000 796.110 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 803.190 0.000 803.470 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 810.550 0.000 810.830 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 817.910 0.000 818.190 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 825.270 0.000 825.550 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 832.630 0.000 832.910 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 839.990 0.000 840.270 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 310.990 0.000 311.270 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 847.350 0.000 847.630 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 854.710 0.000 854.990 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 862.070 0.000 862.350 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 869.430 0.000 869.710 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.790 0.000 877.070 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 884.150 0.000 884.430 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 891.510 0.000 891.790 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 898.870 0.000 899.150 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 906.230 0.000 906.510 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 913.590 0.000 913.870 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 318.350 0.000 318.630 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 920.950 0.000 921.230 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 927.850 0.000 928.130 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 935.210 0.000 935.490 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 942.570 0.000 942.850 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.930 0.000 950.210 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 957.290 0.000 957.570 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 964.650 0.000 964.930 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 972.010 0.000 972.290 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 979.370 0.000 979.650 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 986.730 0.000 987.010 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 325.710 0.000 325.990 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 261.770 0.000 262.050 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 996.850 0.000 997.130 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1004.210 0.000 1004.490 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1011.570 0.000 1011.850 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1018.470 0.000 1018.750 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1025.830 0.000 1026.110 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1033.190 0.000 1033.470 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1040.550 0.000 1040.830 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1047.910 0.000 1048.190 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1055.270 0.000 1055.550 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1062.630 0.000 1062.910 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 335.370 0.000 335.650 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1069.990 0.000 1070.270 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1077.350 0.000 1077.630 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1084.710 0.000 1084.990 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1092.070 0.000 1092.350 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1099.430 0.000 1099.710 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1106.790 0.000 1107.070 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1114.150 0.000 1114.430 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1121.510 0.000 1121.790 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1128.870 0.000 1129.150 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1136.230 0.000 1136.510 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 342.730 0.000 343.010 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1143.590 0.000 1143.870 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1150.950 0.000 1151.230 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1158.310 0.000 1158.590 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1165.670 0.000 1165.950 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.030 0.000 1173.310 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1180.390 0.000 1180.670 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1187.750 0.000 1188.030 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1195.110 0.000 1195.390 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 350.090 0.000 350.370 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 357.450 0.000 357.730 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.810 0.000 365.090 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 372.170 0.000 372.450 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 379.530 0.000 379.810 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 386.890 0.000 387.170 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 394.250 0.000 394.530 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 401.610 0.000 401.890 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 269.130 0.000 269.410 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 408.970 0.000 409.250 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 416.330 0.000 416.610 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 423.690 0.000 423.970 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 431.050 0.000 431.330 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.410 0.000 438.690 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 445.770 0.000 446.050 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 453.130 0.000 453.410 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 460.490 0.000 460.770 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 467.390 0.000 467.670 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 474.750 0.000 475.030 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 276.490 0.000 276.770 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 482.110 0.000 482.390 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.470 0.000 489.750 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 496.830 0.000 497.110 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 504.190 0.000 504.470 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 511.550 0.000 511.830 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 518.910 0.000 519.190 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 526.270 0.000 526.550 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 533.630 0.000 533.910 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 540.990 0.000 541.270 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 548.350 0.000 548.630 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 283.850 0.000 284.130 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.710 0.000 555.990 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 563.070 0.000 563.350 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 570.430 0.000 570.710 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 577.790 0.000 578.070 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 585.150 0.000 585.430 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 592.510 0.000 592.790 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 599.870 0.000 600.150 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 607.230 0.000 607.510 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 614.590 0.000 614.870 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 621.950 0.000 622.230 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 291.210 0.000 291.490 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 629.310 0.000 629.590 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 636.670 0.000 636.950 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 644.030 0.000 644.310 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 651.390 0.000 651.670 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 658.750 0.000 659.030 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 666.110 0.000 666.390 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 673.470 0.000 673.750 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 680.830 0.000 681.110 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 688.190 0.000 688.470 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 695.550 0.000 695.830 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 298.570 0.000 298.850 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 702.910 0.000 703.190 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 710.270 0.000 710.550 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 717.630 0.000 717.910 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 724.990 0.000 725.270 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 732.350 0.000 732.630 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 739.250 0.000 739.530 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.610 0.000 746.890 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 753.970 0.000 754.250 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 761.330 0.000 761.610 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 768.690 0.000 768.970 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.930 0.000 306.210 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 776.050 0.000 776.330 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 783.410 0.000 783.690 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 790.770 0.000 791.050 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 798.130 0.000 798.410 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 805.490 0.000 805.770 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 812.850 0.000 813.130 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 820.210 0.000 820.490 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 827.570 0.000 827.850 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 834.930 0.000 835.210 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 842.290 0.000 842.570 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 313.290 0.000 313.570 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 849.650 0.000 849.930 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 857.010 0.000 857.290 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 864.370 0.000 864.650 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 871.730 0.000 872.010 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 879.090 0.000 879.370 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 886.450 0.000 886.730 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 893.810 0.000 894.090 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 901.170 0.000 901.450 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 908.530 0.000 908.810 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 915.890 0.000 916.170 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 320.650 0.000 320.930 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 923.250 0.000 923.530 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 930.610 0.000 930.890 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 937.970 0.000 938.250 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 945.330 0.000 945.610 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 952.690 0.000 952.970 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 960.050 0.000 960.330 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 967.410 0.000 967.690 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 974.770 0.000 975.050 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 982.130 0.000 982.410 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 989.490 0.000 989.770 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 328.010 0.000 328.290 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.530 0.000 264.810 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 999.150 0.000 999.430 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1006.510 0.000 1006.790 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1013.870 0.000 1014.150 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1021.230 0.000 1021.510 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1028.590 0.000 1028.870 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1035.950 0.000 1036.230 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.310 0.000 1043.590 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1050.670 0.000 1050.950 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1058.030 0.000 1058.310 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1065.390 0.000 1065.670 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.670 0.000 337.950 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1072.750 0.000 1073.030 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1080.110 0.000 1080.390 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1087.470 0.000 1087.750 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1094.830 0.000 1095.110 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1102.190 0.000 1102.470 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1109.090 0.000 1109.370 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1116.450 0.000 1116.730 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1123.810 0.000 1124.090 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1131.170 0.000 1131.450 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1138.530 0.000 1138.810 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.030 0.000 345.310 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1145.890 0.000 1146.170 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1153.250 0.000 1153.530 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1160.610 0.000 1160.890 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1167.970 0.000 1168.250 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1175.330 0.000 1175.610 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1182.690 0.000 1182.970 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1190.050 0.000 1190.330 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1197.410 0.000 1197.690 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 352.390 0.000 352.670 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 359.750 0.000 360.030 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 367.110 0.000 367.390 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 374.470 0.000 374.750 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.830 0.000 382.110 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 389.190 0.000 389.470 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 396.550 0.000 396.830 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.910 0.000 404.190 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.890 0.000 272.170 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 411.270 0.000 411.550 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 418.630 0.000 418.910 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 425.990 0.000 426.270 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 433.350 0.000 433.630 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 440.710 0.000 440.990 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 448.070 0.000 448.350 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.430 0.000 455.710 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.790 0.000 463.070 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 470.150 0.000 470.430 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.510 0.000 477.790 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 278.790 0.000 279.070 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 484.870 0.000 485.150 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 492.230 0.000 492.510 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 499.590 0.000 499.870 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 506.950 0.000 507.230 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 514.310 0.000 514.590 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 521.670 0.000 521.950 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 529.030 0.000 529.310 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 536.390 0.000 536.670 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 543.750 0.000 544.030 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 551.110 0.000 551.390 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 286.150 0.000 286.430 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 558.010 0.000 558.290 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 565.370 0.000 565.650 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 572.730 0.000 573.010 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 580.090 0.000 580.370 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.450 0.000 587.730 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 594.810 0.000 595.090 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 602.170 0.000 602.450 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 609.530 0.000 609.810 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 616.890 0.000 617.170 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 624.250 0.000 624.530 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.510 0.000 293.790 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 631.610 0.000 631.890 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 638.970 0.000 639.250 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 646.330 0.000 646.610 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 653.690 0.000 653.970 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 661.050 0.000 661.330 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.410 0.000 668.690 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 675.770 0.000 676.050 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 683.130 0.000 683.410 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 690.490 0.000 690.770 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 697.850 0.000 698.130 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.870 0.000 301.150 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 705.210 0.000 705.490 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 712.570 0.000 712.850 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 719.930 0.000 720.210 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 727.290 0.000 727.570 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.650 0.000 734.930 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 742.010 0.000 742.290 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 749.370 0.000 749.650 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 756.730 0.000 757.010 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 764.090 0.000 764.370 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 771.450 0.000 771.730 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 308.230 0.000 308.510 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 778.810 0.000 779.090 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 786.170 0.000 786.450 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 793.530 0.000 793.810 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 800.890 0.000 801.170 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 808.250 0.000 808.530 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 815.610 0.000 815.890 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 822.970 0.000 823.250 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 830.330 0.000 830.610 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 837.230 0.000 837.510 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 844.590 0.000 844.870 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 315.590 0.000 315.870 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 851.950 0.000 852.230 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 859.310 0.000 859.590 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 866.670 0.000 866.950 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 874.030 0.000 874.310 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 881.390 0.000 881.670 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 888.750 0.000 889.030 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.110 0.000 896.390 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 903.470 0.000 903.750 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 910.830 0.000 911.110 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.190 0.000 918.470 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.950 0.000 323.230 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 925.550 0.000 925.830 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 932.910 0.000 933.190 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 940.270 0.000 940.550 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 947.630 0.000 947.910 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 954.990 0.000 955.270 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 962.350 0.000 962.630 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 969.710 0.000 969.990 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 977.070 0.000 977.350 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.430 0.000 984.710 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 991.790 0.000 992.070 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 330.310 0.000 330.590 4.000 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.030 0.000 0.310 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.330 0.000 2.610 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.630 0.000 4.910 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 14.290 0.000 14.570 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 97.550 0.000 97.830 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.910 0.000 105.190 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.270 0.000 112.550 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.630 0.000 119.910 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.990 0.000 127.270 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 134.350 0.000 134.630 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 141.710 0.000 141.990 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.070 0.000 149.350 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.430 0.000 156.710 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 163.790 0.000 164.070 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.410 0.000 24.690 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 171.150 0.000 171.430 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.510 0.000 178.790 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.870 0.000 186.150 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 193.230 0.000 193.510 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.590 0.000 200.870 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 207.950 0.000 208.230 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.310 0.000 215.590 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 222.670 0.000 222.950 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 230.030 0.000 230.310 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 237.390 0.000 237.670 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.070 0.000 34.350 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.750 0.000 245.030 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 252.110 0.000 252.390 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.730 0.000 44.010 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.850 0.000 54.130 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.210 0.000 61.490 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.570 0.000 68.850 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.930 0.000 76.210 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.290 0.000 83.570 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.650 0.000 90.930 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.930 0.000 7.210 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 17.050 0.000 17.330 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.310 0.000 100.590 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 107.670 0.000 107.950 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 115.030 0.000 115.310 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.390 0.000 122.670 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 129.750 0.000 130.030 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.110 0.000 137.390 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.470 0.000 144.750 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.830 0.000 152.110 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.190 0.000 159.470 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.550 0.000 166.830 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.710 0.000 26.990 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.910 0.000 174.190 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 181.270 0.000 181.550 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 188.170 0.000 188.450 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 195.530 0.000 195.810 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.890 0.000 203.170 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.250 0.000 210.530 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.610 0.000 217.890 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.970 0.000 225.250 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 232.330 0.000 232.610 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 239.690 0.000 239.970 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 36.370 0.000 36.650 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.050 0.000 247.330 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.410 0.000 254.690 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.490 0.000 46.770 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.150 0.000 56.430 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 63.510 0.000 63.790 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.870 0.000 71.150 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.230 0.000 78.510 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.590 0.000 85.870 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.950 0.000 93.230 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 19.350 0.000 19.630 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.610 0.000 102.890 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.970 0.000 110.250 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.330 0.000 117.610 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.690 0.000 124.970 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.050 0.000 132.330 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.410 0.000 139.690 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.770 0.000 147.050 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 154.130 0.000 154.410 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 161.490 0.000 161.770 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 168.850 0.000 169.130 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.010 0.000 29.290 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.210 0.000 176.490 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.570 0.000 183.850 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 190.930 0.000 191.210 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 198.290 0.000 198.570 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 205.650 0.000 205.930 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.010 0.000 213.290 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 220.370 0.000 220.650 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 227.730 0.000 228.010 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 235.090 0.000 235.370 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 242.450 0.000 242.730 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.130 0.000 39.410 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 249.810 0.000 250.090 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 257.170 0.000 257.450 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 48.790 0.000 49.070 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 58.450 0.000 58.730 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 65.810 0.000 66.090 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.170 0.000 73.450 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.530 0.000 80.810 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.890 0.000 88.170 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 95.250 0.000 95.530 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 21.650 0.000 21.930 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.770 0.000 32.050 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.430 0.000 41.710 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.090 0.000 51.370 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.690 0.000 9.970 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.990 0.000 12.270 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.060 10.640 21.660 1188.880 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.860 10.640 98.460 1188.880 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.540 10.795 1193.180 1188.725 ;
      LAYER met1 ;
        RECT 4.540 5.480 1197.710 1188.880 ;
      LAYER met2 ;
        RECT 0.030 1195.720 3.890 1196.000 ;
        RECT 4.730 1195.720 14.010 1196.000 ;
        RECT 14.850 1195.720 24.590 1196.000 ;
        RECT 25.430 1195.720 35.170 1196.000 ;
        RECT 36.010 1195.720 45.750 1196.000 ;
        RECT 46.590 1195.720 56.330 1196.000 ;
        RECT 57.170 1195.720 66.910 1196.000 ;
        RECT 67.750 1195.720 77.490 1196.000 ;
        RECT 78.330 1195.720 88.070 1196.000 ;
        RECT 88.910 1195.720 98.190 1196.000 ;
        RECT 99.030 1195.720 108.770 1196.000 ;
        RECT 109.610 1195.720 119.350 1196.000 ;
        RECT 120.190 1195.720 129.930 1196.000 ;
        RECT 130.770 1195.720 140.510 1196.000 ;
        RECT 141.350 1195.720 151.090 1196.000 ;
        RECT 151.930 1195.720 161.670 1196.000 ;
        RECT 162.510 1195.720 172.250 1196.000 ;
        RECT 173.090 1195.720 182.830 1196.000 ;
        RECT 183.670 1195.720 192.950 1196.000 ;
        RECT 193.790 1195.720 203.530 1196.000 ;
        RECT 204.370 1195.720 214.110 1196.000 ;
        RECT 214.950 1195.720 224.690 1196.000 ;
        RECT 225.530 1195.720 235.270 1196.000 ;
        RECT 236.110 1195.720 245.850 1196.000 ;
        RECT 246.690 1195.720 256.430 1196.000 ;
        RECT 257.270 1195.720 267.010 1196.000 ;
        RECT 267.850 1195.720 277.590 1196.000 ;
        RECT 278.430 1195.720 287.710 1196.000 ;
        RECT 288.550 1195.720 298.290 1196.000 ;
        RECT 299.130 1195.720 308.870 1196.000 ;
        RECT 309.710 1195.720 319.450 1196.000 ;
        RECT 320.290 1195.720 330.030 1196.000 ;
        RECT 330.870 1195.720 340.610 1196.000 ;
        RECT 341.450 1195.720 351.190 1196.000 ;
        RECT 352.030 1195.720 361.770 1196.000 ;
        RECT 362.610 1195.720 372.350 1196.000 ;
        RECT 373.190 1195.720 382.470 1196.000 ;
        RECT 383.310 1195.720 393.050 1196.000 ;
        RECT 393.890 1195.720 403.630 1196.000 ;
        RECT 404.470 1195.720 414.210 1196.000 ;
        RECT 415.050 1195.720 424.790 1196.000 ;
        RECT 425.630 1195.720 435.370 1196.000 ;
        RECT 436.210 1195.720 445.950 1196.000 ;
        RECT 446.790 1195.720 456.530 1196.000 ;
        RECT 457.370 1195.720 466.650 1196.000 ;
        RECT 467.490 1195.720 477.230 1196.000 ;
        RECT 478.070 1195.720 487.810 1196.000 ;
        RECT 488.650 1195.720 498.390 1196.000 ;
        RECT 499.230 1195.720 508.970 1196.000 ;
        RECT 509.810 1195.720 519.550 1196.000 ;
        RECT 520.390 1195.720 530.130 1196.000 ;
        RECT 530.970 1195.720 540.710 1196.000 ;
        RECT 541.550 1195.720 551.290 1196.000 ;
        RECT 552.130 1195.720 561.410 1196.000 ;
        RECT 562.250 1195.720 571.990 1196.000 ;
        RECT 572.830 1195.720 582.570 1196.000 ;
        RECT 583.410 1195.720 593.150 1196.000 ;
        RECT 593.990 1195.720 603.730 1196.000 ;
        RECT 604.570 1195.720 614.310 1196.000 ;
        RECT 615.150 1195.720 624.890 1196.000 ;
        RECT 625.730 1195.720 635.470 1196.000 ;
        RECT 636.310 1195.720 646.050 1196.000 ;
        RECT 646.890 1195.720 656.170 1196.000 ;
        RECT 657.010 1195.720 666.750 1196.000 ;
        RECT 667.590 1195.720 677.330 1196.000 ;
        RECT 678.170 1195.720 687.910 1196.000 ;
        RECT 688.750 1195.720 698.490 1196.000 ;
        RECT 699.330 1195.720 709.070 1196.000 ;
        RECT 709.910 1195.720 719.650 1196.000 ;
        RECT 720.490 1195.720 730.230 1196.000 ;
        RECT 731.070 1195.720 740.810 1196.000 ;
        RECT 741.650 1195.720 750.930 1196.000 ;
        RECT 751.770 1195.720 761.510 1196.000 ;
        RECT 762.350 1195.720 772.090 1196.000 ;
        RECT 772.930 1195.720 782.670 1196.000 ;
        RECT 783.510 1195.720 793.250 1196.000 ;
        RECT 794.090 1195.720 803.830 1196.000 ;
        RECT 804.670 1195.720 814.410 1196.000 ;
        RECT 815.250 1195.720 824.990 1196.000 ;
        RECT 825.830 1195.720 835.110 1196.000 ;
        RECT 835.950 1195.720 845.690 1196.000 ;
        RECT 846.530 1195.720 856.270 1196.000 ;
        RECT 857.110 1195.720 866.850 1196.000 ;
        RECT 867.690 1195.720 877.430 1196.000 ;
        RECT 878.270 1195.720 888.010 1196.000 ;
        RECT 888.850 1195.720 898.590 1196.000 ;
        RECT 899.430 1195.720 909.170 1196.000 ;
        RECT 910.010 1195.720 919.750 1196.000 ;
        RECT 920.590 1195.720 929.870 1196.000 ;
        RECT 930.710 1195.720 940.450 1196.000 ;
        RECT 941.290 1195.720 951.030 1196.000 ;
        RECT 951.870 1195.720 961.610 1196.000 ;
        RECT 962.450 1195.720 972.190 1196.000 ;
        RECT 973.030 1195.720 982.770 1196.000 ;
        RECT 983.610 1195.720 993.350 1196.000 ;
        RECT 994.190 1195.720 1003.930 1196.000 ;
        RECT 1004.770 1195.720 1014.510 1196.000 ;
        RECT 1015.350 1195.720 1024.630 1196.000 ;
        RECT 1025.470 1195.720 1035.210 1196.000 ;
        RECT 1036.050 1195.720 1045.790 1196.000 ;
        RECT 1046.630 1195.720 1056.370 1196.000 ;
        RECT 1057.210 1195.720 1066.950 1196.000 ;
        RECT 1067.790 1195.720 1077.530 1196.000 ;
        RECT 1078.370 1195.720 1088.110 1196.000 ;
        RECT 1088.950 1195.720 1098.690 1196.000 ;
        RECT 1099.530 1195.720 1109.270 1196.000 ;
        RECT 1110.110 1195.720 1119.390 1196.000 ;
        RECT 1120.230 1195.720 1129.970 1196.000 ;
        RECT 1130.810 1195.720 1140.550 1196.000 ;
        RECT 1141.390 1195.720 1151.130 1196.000 ;
        RECT 1151.970 1195.720 1161.710 1196.000 ;
        RECT 1162.550 1195.720 1172.290 1196.000 ;
        RECT 1173.130 1195.720 1182.870 1196.000 ;
        RECT 1183.710 1195.720 1193.450 1196.000 ;
        RECT 1194.290 1195.720 1197.680 1196.000 ;
        RECT 0.030 4.280 1197.680 1195.720 ;
        RECT 0.590 4.000 2.050 4.280 ;
        RECT 2.890 4.000 4.350 4.280 ;
        RECT 5.190 4.000 6.650 4.280 ;
        RECT 7.490 4.000 9.410 4.280 ;
        RECT 10.250 4.000 11.710 4.280 ;
        RECT 12.550 4.000 14.010 4.280 ;
        RECT 14.850 4.000 16.770 4.280 ;
        RECT 17.610 4.000 19.070 4.280 ;
        RECT 19.910 4.000 21.370 4.280 ;
        RECT 22.210 4.000 24.130 4.280 ;
        RECT 24.970 4.000 26.430 4.280 ;
        RECT 27.270 4.000 28.730 4.280 ;
        RECT 29.570 4.000 31.490 4.280 ;
        RECT 32.330 4.000 33.790 4.280 ;
        RECT 34.630 4.000 36.090 4.280 ;
        RECT 36.930 4.000 38.850 4.280 ;
        RECT 39.690 4.000 41.150 4.280 ;
        RECT 41.990 4.000 43.450 4.280 ;
        RECT 44.290 4.000 46.210 4.280 ;
        RECT 47.050 4.000 48.510 4.280 ;
        RECT 49.350 4.000 50.810 4.280 ;
        RECT 51.650 4.000 53.570 4.280 ;
        RECT 54.410 4.000 55.870 4.280 ;
        RECT 56.710 4.000 58.170 4.280 ;
        RECT 59.010 4.000 60.930 4.280 ;
        RECT 61.770 4.000 63.230 4.280 ;
        RECT 64.070 4.000 65.530 4.280 ;
        RECT 66.370 4.000 68.290 4.280 ;
        RECT 69.130 4.000 70.590 4.280 ;
        RECT 71.430 4.000 72.890 4.280 ;
        RECT 73.730 4.000 75.650 4.280 ;
        RECT 76.490 4.000 77.950 4.280 ;
        RECT 78.790 4.000 80.250 4.280 ;
        RECT 81.090 4.000 83.010 4.280 ;
        RECT 83.850 4.000 85.310 4.280 ;
        RECT 86.150 4.000 87.610 4.280 ;
        RECT 88.450 4.000 90.370 4.280 ;
        RECT 91.210 4.000 92.670 4.280 ;
        RECT 93.510 4.000 94.970 4.280 ;
        RECT 95.810 4.000 97.270 4.280 ;
        RECT 98.110 4.000 100.030 4.280 ;
        RECT 100.870 4.000 102.330 4.280 ;
        RECT 103.170 4.000 104.630 4.280 ;
        RECT 105.470 4.000 107.390 4.280 ;
        RECT 108.230 4.000 109.690 4.280 ;
        RECT 110.530 4.000 111.990 4.280 ;
        RECT 112.830 4.000 114.750 4.280 ;
        RECT 115.590 4.000 117.050 4.280 ;
        RECT 117.890 4.000 119.350 4.280 ;
        RECT 120.190 4.000 122.110 4.280 ;
        RECT 122.950 4.000 124.410 4.280 ;
        RECT 125.250 4.000 126.710 4.280 ;
        RECT 127.550 4.000 129.470 4.280 ;
        RECT 130.310 4.000 131.770 4.280 ;
        RECT 132.610 4.000 134.070 4.280 ;
        RECT 134.910 4.000 136.830 4.280 ;
        RECT 137.670 4.000 139.130 4.280 ;
        RECT 139.970 4.000 141.430 4.280 ;
        RECT 142.270 4.000 144.190 4.280 ;
        RECT 145.030 4.000 146.490 4.280 ;
        RECT 147.330 4.000 148.790 4.280 ;
        RECT 149.630 4.000 151.550 4.280 ;
        RECT 152.390 4.000 153.850 4.280 ;
        RECT 154.690 4.000 156.150 4.280 ;
        RECT 156.990 4.000 158.910 4.280 ;
        RECT 159.750 4.000 161.210 4.280 ;
        RECT 162.050 4.000 163.510 4.280 ;
        RECT 164.350 4.000 166.270 4.280 ;
        RECT 167.110 4.000 168.570 4.280 ;
        RECT 169.410 4.000 170.870 4.280 ;
        RECT 171.710 4.000 173.630 4.280 ;
        RECT 174.470 4.000 175.930 4.280 ;
        RECT 176.770 4.000 178.230 4.280 ;
        RECT 179.070 4.000 180.990 4.280 ;
        RECT 181.830 4.000 183.290 4.280 ;
        RECT 184.130 4.000 185.590 4.280 ;
        RECT 186.430 4.000 187.890 4.280 ;
        RECT 188.730 4.000 190.650 4.280 ;
        RECT 191.490 4.000 192.950 4.280 ;
        RECT 193.790 4.000 195.250 4.280 ;
        RECT 196.090 4.000 198.010 4.280 ;
        RECT 198.850 4.000 200.310 4.280 ;
        RECT 201.150 4.000 202.610 4.280 ;
        RECT 203.450 4.000 205.370 4.280 ;
        RECT 206.210 4.000 207.670 4.280 ;
        RECT 208.510 4.000 209.970 4.280 ;
        RECT 210.810 4.000 212.730 4.280 ;
        RECT 213.570 4.000 215.030 4.280 ;
        RECT 215.870 4.000 217.330 4.280 ;
        RECT 218.170 4.000 220.090 4.280 ;
        RECT 220.930 4.000 222.390 4.280 ;
        RECT 223.230 4.000 224.690 4.280 ;
        RECT 225.530 4.000 227.450 4.280 ;
        RECT 228.290 4.000 229.750 4.280 ;
        RECT 230.590 4.000 232.050 4.280 ;
        RECT 232.890 4.000 234.810 4.280 ;
        RECT 235.650 4.000 237.110 4.280 ;
        RECT 237.950 4.000 239.410 4.280 ;
        RECT 240.250 4.000 242.170 4.280 ;
        RECT 243.010 4.000 244.470 4.280 ;
        RECT 245.310 4.000 246.770 4.280 ;
        RECT 247.610 4.000 249.530 4.280 ;
        RECT 250.370 4.000 251.830 4.280 ;
        RECT 252.670 4.000 254.130 4.280 ;
        RECT 254.970 4.000 256.890 4.280 ;
        RECT 257.730 4.000 259.190 4.280 ;
        RECT 260.030 4.000 261.490 4.280 ;
        RECT 262.330 4.000 264.250 4.280 ;
        RECT 265.090 4.000 266.550 4.280 ;
        RECT 267.390 4.000 268.850 4.280 ;
        RECT 269.690 4.000 271.610 4.280 ;
        RECT 272.450 4.000 273.910 4.280 ;
        RECT 274.750 4.000 276.210 4.280 ;
        RECT 277.050 4.000 278.510 4.280 ;
        RECT 279.350 4.000 281.270 4.280 ;
        RECT 282.110 4.000 283.570 4.280 ;
        RECT 284.410 4.000 285.870 4.280 ;
        RECT 286.710 4.000 288.630 4.280 ;
        RECT 289.470 4.000 290.930 4.280 ;
        RECT 291.770 4.000 293.230 4.280 ;
        RECT 294.070 4.000 295.990 4.280 ;
        RECT 296.830 4.000 298.290 4.280 ;
        RECT 299.130 4.000 300.590 4.280 ;
        RECT 301.430 4.000 303.350 4.280 ;
        RECT 304.190 4.000 305.650 4.280 ;
        RECT 306.490 4.000 307.950 4.280 ;
        RECT 308.790 4.000 310.710 4.280 ;
        RECT 311.550 4.000 313.010 4.280 ;
        RECT 313.850 4.000 315.310 4.280 ;
        RECT 316.150 4.000 318.070 4.280 ;
        RECT 318.910 4.000 320.370 4.280 ;
        RECT 321.210 4.000 322.670 4.280 ;
        RECT 323.510 4.000 325.430 4.280 ;
        RECT 326.270 4.000 327.730 4.280 ;
        RECT 328.570 4.000 330.030 4.280 ;
        RECT 330.870 4.000 332.790 4.280 ;
        RECT 333.630 4.000 335.090 4.280 ;
        RECT 335.930 4.000 337.390 4.280 ;
        RECT 338.230 4.000 340.150 4.280 ;
        RECT 340.990 4.000 342.450 4.280 ;
        RECT 343.290 4.000 344.750 4.280 ;
        RECT 345.590 4.000 347.510 4.280 ;
        RECT 348.350 4.000 349.810 4.280 ;
        RECT 350.650 4.000 352.110 4.280 ;
        RECT 352.950 4.000 354.870 4.280 ;
        RECT 355.710 4.000 357.170 4.280 ;
        RECT 358.010 4.000 359.470 4.280 ;
        RECT 360.310 4.000 362.230 4.280 ;
        RECT 363.070 4.000 364.530 4.280 ;
        RECT 365.370 4.000 366.830 4.280 ;
        RECT 367.670 4.000 369.130 4.280 ;
        RECT 369.970 4.000 371.890 4.280 ;
        RECT 372.730 4.000 374.190 4.280 ;
        RECT 375.030 4.000 376.490 4.280 ;
        RECT 377.330 4.000 379.250 4.280 ;
        RECT 380.090 4.000 381.550 4.280 ;
        RECT 382.390 4.000 383.850 4.280 ;
        RECT 384.690 4.000 386.610 4.280 ;
        RECT 387.450 4.000 388.910 4.280 ;
        RECT 389.750 4.000 391.210 4.280 ;
        RECT 392.050 4.000 393.970 4.280 ;
        RECT 394.810 4.000 396.270 4.280 ;
        RECT 397.110 4.000 398.570 4.280 ;
        RECT 399.410 4.000 401.330 4.280 ;
        RECT 402.170 4.000 403.630 4.280 ;
        RECT 404.470 4.000 405.930 4.280 ;
        RECT 406.770 4.000 408.690 4.280 ;
        RECT 409.530 4.000 410.990 4.280 ;
        RECT 411.830 4.000 413.290 4.280 ;
        RECT 414.130 4.000 416.050 4.280 ;
        RECT 416.890 4.000 418.350 4.280 ;
        RECT 419.190 4.000 420.650 4.280 ;
        RECT 421.490 4.000 423.410 4.280 ;
        RECT 424.250 4.000 425.710 4.280 ;
        RECT 426.550 4.000 428.010 4.280 ;
        RECT 428.850 4.000 430.770 4.280 ;
        RECT 431.610 4.000 433.070 4.280 ;
        RECT 433.910 4.000 435.370 4.280 ;
        RECT 436.210 4.000 438.130 4.280 ;
        RECT 438.970 4.000 440.430 4.280 ;
        RECT 441.270 4.000 442.730 4.280 ;
        RECT 443.570 4.000 445.490 4.280 ;
        RECT 446.330 4.000 447.790 4.280 ;
        RECT 448.630 4.000 450.090 4.280 ;
        RECT 450.930 4.000 452.850 4.280 ;
        RECT 453.690 4.000 455.150 4.280 ;
        RECT 455.990 4.000 457.450 4.280 ;
        RECT 458.290 4.000 460.210 4.280 ;
        RECT 461.050 4.000 462.510 4.280 ;
        RECT 463.350 4.000 464.810 4.280 ;
        RECT 465.650 4.000 467.110 4.280 ;
        RECT 467.950 4.000 469.870 4.280 ;
        RECT 470.710 4.000 472.170 4.280 ;
        RECT 473.010 4.000 474.470 4.280 ;
        RECT 475.310 4.000 477.230 4.280 ;
        RECT 478.070 4.000 479.530 4.280 ;
        RECT 480.370 4.000 481.830 4.280 ;
        RECT 482.670 4.000 484.590 4.280 ;
        RECT 485.430 4.000 486.890 4.280 ;
        RECT 487.730 4.000 489.190 4.280 ;
        RECT 490.030 4.000 491.950 4.280 ;
        RECT 492.790 4.000 494.250 4.280 ;
        RECT 495.090 4.000 496.550 4.280 ;
        RECT 497.390 4.000 499.310 4.280 ;
        RECT 500.150 4.000 501.610 4.280 ;
        RECT 502.450 4.000 503.910 4.280 ;
        RECT 504.750 4.000 506.670 4.280 ;
        RECT 507.510 4.000 508.970 4.280 ;
        RECT 509.810 4.000 511.270 4.280 ;
        RECT 512.110 4.000 514.030 4.280 ;
        RECT 514.870 4.000 516.330 4.280 ;
        RECT 517.170 4.000 518.630 4.280 ;
        RECT 519.470 4.000 521.390 4.280 ;
        RECT 522.230 4.000 523.690 4.280 ;
        RECT 524.530 4.000 525.990 4.280 ;
        RECT 526.830 4.000 528.750 4.280 ;
        RECT 529.590 4.000 531.050 4.280 ;
        RECT 531.890 4.000 533.350 4.280 ;
        RECT 534.190 4.000 536.110 4.280 ;
        RECT 536.950 4.000 538.410 4.280 ;
        RECT 539.250 4.000 540.710 4.280 ;
        RECT 541.550 4.000 543.470 4.280 ;
        RECT 544.310 4.000 545.770 4.280 ;
        RECT 546.610 4.000 548.070 4.280 ;
        RECT 548.910 4.000 550.830 4.280 ;
        RECT 551.670 4.000 553.130 4.280 ;
        RECT 553.970 4.000 555.430 4.280 ;
        RECT 556.270 4.000 557.730 4.280 ;
        RECT 558.570 4.000 560.490 4.280 ;
        RECT 561.330 4.000 562.790 4.280 ;
        RECT 563.630 4.000 565.090 4.280 ;
        RECT 565.930 4.000 567.850 4.280 ;
        RECT 568.690 4.000 570.150 4.280 ;
        RECT 570.990 4.000 572.450 4.280 ;
        RECT 573.290 4.000 575.210 4.280 ;
        RECT 576.050 4.000 577.510 4.280 ;
        RECT 578.350 4.000 579.810 4.280 ;
        RECT 580.650 4.000 582.570 4.280 ;
        RECT 583.410 4.000 584.870 4.280 ;
        RECT 585.710 4.000 587.170 4.280 ;
        RECT 588.010 4.000 589.930 4.280 ;
        RECT 590.770 4.000 592.230 4.280 ;
        RECT 593.070 4.000 594.530 4.280 ;
        RECT 595.370 4.000 597.290 4.280 ;
        RECT 598.130 4.000 599.590 4.280 ;
        RECT 600.430 4.000 601.890 4.280 ;
        RECT 602.730 4.000 604.650 4.280 ;
        RECT 605.490 4.000 606.950 4.280 ;
        RECT 607.790 4.000 609.250 4.280 ;
        RECT 610.090 4.000 612.010 4.280 ;
        RECT 612.850 4.000 614.310 4.280 ;
        RECT 615.150 4.000 616.610 4.280 ;
        RECT 617.450 4.000 619.370 4.280 ;
        RECT 620.210 4.000 621.670 4.280 ;
        RECT 622.510 4.000 623.970 4.280 ;
        RECT 624.810 4.000 626.730 4.280 ;
        RECT 627.570 4.000 629.030 4.280 ;
        RECT 629.870 4.000 631.330 4.280 ;
        RECT 632.170 4.000 634.090 4.280 ;
        RECT 634.930 4.000 636.390 4.280 ;
        RECT 637.230 4.000 638.690 4.280 ;
        RECT 639.530 4.000 641.450 4.280 ;
        RECT 642.290 4.000 643.750 4.280 ;
        RECT 644.590 4.000 646.050 4.280 ;
        RECT 646.890 4.000 648.350 4.280 ;
        RECT 649.190 4.000 651.110 4.280 ;
        RECT 651.950 4.000 653.410 4.280 ;
        RECT 654.250 4.000 655.710 4.280 ;
        RECT 656.550 4.000 658.470 4.280 ;
        RECT 659.310 4.000 660.770 4.280 ;
        RECT 661.610 4.000 663.070 4.280 ;
        RECT 663.910 4.000 665.830 4.280 ;
        RECT 666.670 4.000 668.130 4.280 ;
        RECT 668.970 4.000 670.430 4.280 ;
        RECT 671.270 4.000 673.190 4.280 ;
        RECT 674.030 4.000 675.490 4.280 ;
        RECT 676.330 4.000 677.790 4.280 ;
        RECT 678.630 4.000 680.550 4.280 ;
        RECT 681.390 4.000 682.850 4.280 ;
        RECT 683.690 4.000 685.150 4.280 ;
        RECT 685.990 4.000 687.910 4.280 ;
        RECT 688.750 4.000 690.210 4.280 ;
        RECT 691.050 4.000 692.510 4.280 ;
        RECT 693.350 4.000 695.270 4.280 ;
        RECT 696.110 4.000 697.570 4.280 ;
        RECT 698.410 4.000 699.870 4.280 ;
        RECT 700.710 4.000 702.630 4.280 ;
        RECT 703.470 4.000 704.930 4.280 ;
        RECT 705.770 4.000 707.230 4.280 ;
        RECT 708.070 4.000 709.990 4.280 ;
        RECT 710.830 4.000 712.290 4.280 ;
        RECT 713.130 4.000 714.590 4.280 ;
        RECT 715.430 4.000 717.350 4.280 ;
        RECT 718.190 4.000 719.650 4.280 ;
        RECT 720.490 4.000 721.950 4.280 ;
        RECT 722.790 4.000 724.710 4.280 ;
        RECT 725.550 4.000 727.010 4.280 ;
        RECT 727.850 4.000 729.310 4.280 ;
        RECT 730.150 4.000 732.070 4.280 ;
        RECT 732.910 4.000 734.370 4.280 ;
        RECT 735.210 4.000 736.670 4.280 ;
        RECT 737.510 4.000 738.970 4.280 ;
        RECT 739.810 4.000 741.730 4.280 ;
        RECT 742.570 4.000 744.030 4.280 ;
        RECT 744.870 4.000 746.330 4.280 ;
        RECT 747.170 4.000 749.090 4.280 ;
        RECT 749.930 4.000 751.390 4.280 ;
        RECT 752.230 4.000 753.690 4.280 ;
        RECT 754.530 4.000 756.450 4.280 ;
        RECT 757.290 4.000 758.750 4.280 ;
        RECT 759.590 4.000 761.050 4.280 ;
        RECT 761.890 4.000 763.810 4.280 ;
        RECT 764.650 4.000 766.110 4.280 ;
        RECT 766.950 4.000 768.410 4.280 ;
        RECT 769.250 4.000 771.170 4.280 ;
        RECT 772.010 4.000 773.470 4.280 ;
        RECT 774.310 4.000 775.770 4.280 ;
        RECT 776.610 4.000 778.530 4.280 ;
        RECT 779.370 4.000 780.830 4.280 ;
        RECT 781.670 4.000 783.130 4.280 ;
        RECT 783.970 4.000 785.890 4.280 ;
        RECT 786.730 4.000 788.190 4.280 ;
        RECT 789.030 4.000 790.490 4.280 ;
        RECT 791.330 4.000 793.250 4.280 ;
        RECT 794.090 4.000 795.550 4.280 ;
        RECT 796.390 4.000 797.850 4.280 ;
        RECT 798.690 4.000 800.610 4.280 ;
        RECT 801.450 4.000 802.910 4.280 ;
        RECT 803.750 4.000 805.210 4.280 ;
        RECT 806.050 4.000 807.970 4.280 ;
        RECT 808.810 4.000 810.270 4.280 ;
        RECT 811.110 4.000 812.570 4.280 ;
        RECT 813.410 4.000 815.330 4.280 ;
        RECT 816.170 4.000 817.630 4.280 ;
        RECT 818.470 4.000 819.930 4.280 ;
        RECT 820.770 4.000 822.690 4.280 ;
        RECT 823.530 4.000 824.990 4.280 ;
        RECT 825.830 4.000 827.290 4.280 ;
        RECT 828.130 4.000 830.050 4.280 ;
        RECT 830.890 4.000 832.350 4.280 ;
        RECT 833.190 4.000 834.650 4.280 ;
        RECT 835.490 4.000 836.950 4.280 ;
        RECT 837.790 4.000 839.710 4.280 ;
        RECT 840.550 4.000 842.010 4.280 ;
        RECT 842.850 4.000 844.310 4.280 ;
        RECT 845.150 4.000 847.070 4.280 ;
        RECT 847.910 4.000 849.370 4.280 ;
        RECT 850.210 4.000 851.670 4.280 ;
        RECT 852.510 4.000 854.430 4.280 ;
        RECT 855.270 4.000 856.730 4.280 ;
        RECT 857.570 4.000 859.030 4.280 ;
        RECT 859.870 4.000 861.790 4.280 ;
        RECT 862.630 4.000 864.090 4.280 ;
        RECT 864.930 4.000 866.390 4.280 ;
        RECT 867.230 4.000 869.150 4.280 ;
        RECT 869.990 4.000 871.450 4.280 ;
        RECT 872.290 4.000 873.750 4.280 ;
        RECT 874.590 4.000 876.510 4.280 ;
        RECT 877.350 4.000 878.810 4.280 ;
        RECT 879.650 4.000 881.110 4.280 ;
        RECT 881.950 4.000 883.870 4.280 ;
        RECT 884.710 4.000 886.170 4.280 ;
        RECT 887.010 4.000 888.470 4.280 ;
        RECT 889.310 4.000 891.230 4.280 ;
        RECT 892.070 4.000 893.530 4.280 ;
        RECT 894.370 4.000 895.830 4.280 ;
        RECT 896.670 4.000 898.590 4.280 ;
        RECT 899.430 4.000 900.890 4.280 ;
        RECT 901.730 4.000 903.190 4.280 ;
        RECT 904.030 4.000 905.950 4.280 ;
        RECT 906.790 4.000 908.250 4.280 ;
        RECT 909.090 4.000 910.550 4.280 ;
        RECT 911.390 4.000 913.310 4.280 ;
        RECT 914.150 4.000 915.610 4.280 ;
        RECT 916.450 4.000 917.910 4.280 ;
        RECT 918.750 4.000 920.670 4.280 ;
        RECT 921.510 4.000 922.970 4.280 ;
        RECT 923.810 4.000 925.270 4.280 ;
        RECT 926.110 4.000 927.570 4.280 ;
        RECT 928.410 4.000 930.330 4.280 ;
        RECT 931.170 4.000 932.630 4.280 ;
        RECT 933.470 4.000 934.930 4.280 ;
        RECT 935.770 4.000 937.690 4.280 ;
        RECT 938.530 4.000 939.990 4.280 ;
        RECT 940.830 4.000 942.290 4.280 ;
        RECT 943.130 4.000 945.050 4.280 ;
        RECT 945.890 4.000 947.350 4.280 ;
        RECT 948.190 4.000 949.650 4.280 ;
        RECT 950.490 4.000 952.410 4.280 ;
        RECT 953.250 4.000 954.710 4.280 ;
        RECT 955.550 4.000 957.010 4.280 ;
        RECT 957.850 4.000 959.770 4.280 ;
        RECT 960.610 4.000 962.070 4.280 ;
        RECT 962.910 4.000 964.370 4.280 ;
        RECT 965.210 4.000 967.130 4.280 ;
        RECT 967.970 4.000 969.430 4.280 ;
        RECT 970.270 4.000 971.730 4.280 ;
        RECT 972.570 4.000 974.490 4.280 ;
        RECT 975.330 4.000 976.790 4.280 ;
        RECT 977.630 4.000 979.090 4.280 ;
        RECT 979.930 4.000 981.850 4.280 ;
        RECT 982.690 4.000 984.150 4.280 ;
        RECT 984.990 4.000 986.450 4.280 ;
        RECT 987.290 4.000 989.210 4.280 ;
        RECT 990.050 4.000 991.510 4.280 ;
        RECT 992.350 4.000 993.810 4.280 ;
        RECT 994.650 4.000 996.570 4.280 ;
        RECT 997.410 4.000 998.870 4.280 ;
        RECT 999.710 4.000 1001.170 4.280 ;
        RECT 1002.010 4.000 1003.930 4.280 ;
        RECT 1004.770 4.000 1006.230 4.280 ;
        RECT 1007.070 4.000 1008.530 4.280 ;
        RECT 1009.370 4.000 1011.290 4.280 ;
        RECT 1012.130 4.000 1013.590 4.280 ;
        RECT 1014.430 4.000 1015.890 4.280 ;
        RECT 1016.730 4.000 1018.190 4.280 ;
        RECT 1019.030 4.000 1020.950 4.280 ;
        RECT 1021.790 4.000 1023.250 4.280 ;
        RECT 1024.090 4.000 1025.550 4.280 ;
        RECT 1026.390 4.000 1028.310 4.280 ;
        RECT 1029.150 4.000 1030.610 4.280 ;
        RECT 1031.450 4.000 1032.910 4.280 ;
        RECT 1033.750 4.000 1035.670 4.280 ;
        RECT 1036.510 4.000 1037.970 4.280 ;
        RECT 1038.810 4.000 1040.270 4.280 ;
        RECT 1041.110 4.000 1043.030 4.280 ;
        RECT 1043.870 4.000 1045.330 4.280 ;
        RECT 1046.170 4.000 1047.630 4.280 ;
        RECT 1048.470 4.000 1050.390 4.280 ;
        RECT 1051.230 4.000 1052.690 4.280 ;
        RECT 1053.530 4.000 1054.990 4.280 ;
        RECT 1055.830 4.000 1057.750 4.280 ;
        RECT 1058.590 4.000 1060.050 4.280 ;
        RECT 1060.890 4.000 1062.350 4.280 ;
        RECT 1063.190 4.000 1065.110 4.280 ;
        RECT 1065.950 4.000 1067.410 4.280 ;
        RECT 1068.250 4.000 1069.710 4.280 ;
        RECT 1070.550 4.000 1072.470 4.280 ;
        RECT 1073.310 4.000 1074.770 4.280 ;
        RECT 1075.610 4.000 1077.070 4.280 ;
        RECT 1077.910 4.000 1079.830 4.280 ;
        RECT 1080.670 4.000 1082.130 4.280 ;
        RECT 1082.970 4.000 1084.430 4.280 ;
        RECT 1085.270 4.000 1087.190 4.280 ;
        RECT 1088.030 4.000 1089.490 4.280 ;
        RECT 1090.330 4.000 1091.790 4.280 ;
        RECT 1092.630 4.000 1094.550 4.280 ;
        RECT 1095.390 4.000 1096.850 4.280 ;
        RECT 1097.690 4.000 1099.150 4.280 ;
        RECT 1099.990 4.000 1101.910 4.280 ;
        RECT 1102.750 4.000 1104.210 4.280 ;
        RECT 1105.050 4.000 1106.510 4.280 ;
        RECT 1107.350 4.000 1108.810 4.280 ;
        RECT 1109.650 4.000 1111.570 4.280 ;
        RECT 1112.410 4.000 1113.870 4.280 ;
        RECT 1114.710 4.000 1116.170 4.280 ;
        RECT 1117.010 4.000 1118.930 4.280 ;
        RECT 1119.770 4.000 1121.230 4.280 ;
        RECT 1122.070 4.000 1123.530 4.280 ;
        RECT 1124.370 4.000 1126.290 4.280 ;
        RECT 1127.130 4.000 1128.590 4.280 ;
        RECT 1129.430 4.000 1130.890 4.280 ;
        RECT 1131.730 4.000 1133.650 4.280 ;
        RECT 1134.490 4.000 1135.950 4.280 ;
        RECT 1136.790 4.000 1138.250 4.280 ;
        RECT 1139.090 4.000 1141.010 4.280 ;
        RECT 1141.850 4.000 1143.310 4.280 ;
        RECT 1144.150 4.000 1145.610 4.280 ;
        RECT 1146.450 4.000 1148.370 4.280 ;
        RECT 1149.210 4.000 1150.670 4.280 ;
        RECT 1151.510 4.000 1152.970 4.280 ;
        RECT 1153.810 4.000 1155.730 4.280 ;
        RECT 1156.570 4.000 1158.030 4.280 ;
        RECT 1158.870 4.000 1160.330 4.280 ;
        RECT 1161.170 4.000 1163.090 4.280 ;
        RECT 1163.930 4.000 1165.390 4.280 ;
        RECT 1166.230 4.000 1167.690 4.280 ;
        RECT 1168.530 4.000 1170.450 4.280 ;
        RECT 1171.290 4.000 1172.750 4.280 ;
        RECT 1173.590 4.000 1175.050 4.280 ;
        RECT 1175.890 4.000 1177.810 4.280 ;
        RECT 1178.650 4.000 1180.110 4.280 ;
        RECT 1180.950 4.000 1182.410 4.280 ;
        RECT 1183.250 4.000 1185.170 4.280 ;
        RECT 1186.010 4.000 1187.470 4.280 ;
        RECT 1188.310 4.000 1189.770 4.280 ;
        RECT 1190.610 4.000 1192.530 4.280 ;
        RECT 1193.370 4.000 1194.830 4.280 ;
        RECT 1195.670 4.000 1197.130 4.280 ;
      LAYER met3 ;
        RECT 0.005 4.255 1177.935 1188.805 ;
      LAYER met4 ;
        RECT 95.915 10.640 96.460 1188.880 ;
        RECT 98.860 10.640 1173.660 1188.880 ;
  END
END user_proj_example
END LIBRARY

