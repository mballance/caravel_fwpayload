magic
tech sky130A
magscale 1 2
timestamp 1608227625
<< obsli1 >>
rect 906 2159 238634 237745
<< obsm1 >>
rect 0 960 239540 237776
<< metal2 >>
rect 832 239200 888 240000
rect 2856 239200 2912 240000
rect 4972 239200 5028 240000
rect 7088 239200 7144 240000
rect 9204 239200 9260 240000
rect 11320 239200 11376 240000
rect 13436 239200 13492 240000
rect 15552 239200 15608 240000
rect 17668 239200 17724 240000
rect 19692 239200 19748 240000
rect 21808 239200 21864 240000
rect 23924 239200 23980 240000
rect 26040 239200 26096 240000
rect 28156 239200 28212 240000
rect 30272 239200 30328 240000
rect 32388 239200 32444 240000
rect 34504 239200 34560 240000
rect 36620 239200 36676 240000
rect 38644 239200 38700 240000
rect 40760 239200 40816 240000
rect 42876 239200 42932 240000
rect 44992 239200 45048 240000
rect 47108 239200 47164 240000
rect 49224 239200 49280 240000
rect 51340 239200 51396 240000
rect 53456 239200 53512 240000
rect 55572 239200 55628 240000
rect 57596 239200 57652 240000
rect 59712 239200 59768 240000
rect 61828 239200 61884 240000
rect 63944 239200 64000 240000
rect 66060 239200 66116 240000
rect 68176 239200 68232 240000
rect 70292 239200 70348 240000
rect 72408 239200 72464 240000
rect 74524 239200 74580 240000
rect 76548 239200 76604 240000
rect 78664 239200 78720 240000
rect 80780 239200 80836 240000
rect 82896 239200 82952 240000
rect 85012 239200 85068 240000
rect 87128 239200 87184 240000
rect 89244 239200 89300 240000
rect 91360 239200 91416 240000
rect 93384 239200 93440 240000
rect 95500 239200 95556 240000
rect 97616 239200 97672 240000
rect 99732 239200 99788 240000
rect 101848 239200 101904 240000
rect 103964 239200 104020 240000
rect 106080 239200 106136 240000
rect 108196 239200 108252 240000
rect 110312 239200 110368 240000
rect 112336 239200 112392 240000
rect 114452 239200 114508 240000
rect 116568 239200 116624 240000
rect 118684 239200 118740 240000
rect 120800 239200 120856 240000
rect 122916 239200 122972 240000
rect 125032 239200 125088 240000
rect 127148 239200 127204 240000
rect 129264 239200 129320 240000
rect 131288 239200 131344 240000
rect 133404 239200 133460 240000
rect 135520 239200 135576 240000
rect 137636 239200 137692 240000
rect 139752 239200 139808 240000
rect 141868 239200 141924 240000
rect 143984 239200 144040 240000
rect 146100 239200 146156 240000
rect 148216 239200 148272 240000
rect 150240 239200 150296 240000
rect 152356 239200 152412 240000
rect 154472 239200 154528 240000
rect 156588 239200 156644 240000
rect 158704 239200 158760 240000
rect 160820 239200 160876 240000
rect 162936 239200 162992 240000
rect 165052 239200 165108 240000
rect 167076 239200 167132 240000
rect 169192 239200 169248 240000
rect 171308 239200 171364 240000
rect 173424 239200 173480 240000
rect 175540 239200 175596 240000
rect 177656 239200 177712 240000
rect 179772 239200 179828 240000
rect 181888 239200 181944 240000
rect 184004 239200 184060 240000
rect 186028 239200 186084 240000
rect 188144 239200 188200 240000
rect 190260 239200 190316 240000
rect 192376 239200 192432 240000
rect 194492 239200 194548 240000
rect 196608 239200 196664 240000
rect 198724 239200 198780 240000
rect 200840 239200 200896 240000
rect 202956 239200 203012 240000
rect 204980 239200 205036 240000
rect 207096 239200 207152 240000
rect 209212 239200 209268 240000
rect 211328 239200 211384 240000
rect 213444 239200 213500 240000
rect 215560 239200 215616 240000
rect 217676 239200 217732 240000
rect 219792 239200 219848 240000
rect 221908 239200 221964 240000
rect 223932 239200 223988 240000
rect 226048 239200 226104 240000
rect 228164 239200 228220 240000
rect 230280 239200 230336 240000
rect 232396 239200 232452 240000
rect 234512 239200 234568 240000
rect 236628 239200 236684 240000
rect 238744 239200 238800 240000
rect 4 0 60 800
rect 464 0 520 800
rect 924 0 980 800
rect 1384 0 1440 800
rect 1936 0 1992 800
rect 2396 0 2452 800
rect 2856 0 2912 800
rect 3408 0 3464 800
rect 3868 0 3924 800
rect 4328 0 4384 800
rect 4880 0 4936 800
rect 5340 0 5396 800
rect 5800 0 5856 800
rect 6352 0 6408 800
rect 6812 0 6868 800
rect 7272 0 7328 800
rect 7824 0 7880 800
rect 8284 0 8340 800
rect 8744 0 8800 800
rect 9296 0 9352 800
rect 9756 0 9812 800
rect 10216 0 10272 800
rect 10768 0 10824 800
rect 11228 0 11284 800
rect 11688 0 11744 800
rect 12240 0 12296 800
rect 12700 0 12756 800
rect 13160 0 13216 800
rect 13712 0 13768 800
rect 14172 0 14228 800
rect 14632 0 14688 800
rect 15184 0 15240 800
rect 15644 0 15700 800
rect 16104 0 16160 800
rect 16656 0 16712 800
rect 17116 0 17172 800
rect 17576 0 17632 800
rect 18128 0 18184 800
rect 18588 0 18644 800
rect 19048 0 19104 800
rect 19508 0 19564 800
rect 20060 0 20116 800
rect 20520 0 20576 800
rect 20980 0 21036 800
rect 21532 0 21588 800
rect 21992 0 22048 800
rect 22452 0 22508 800
rect 23004 0 23060 800
rect 23464 0 23520 800
rect 23924 0 23980 800
rect 24476 0 24532 800
rect 24936 0 24992 800
rect 25396 0 25452 800
rect 25948 0 26004 800
rect 26408 0 26464 800
rect 26868 0 26924 800
rect 27420 0 27476 800
rect 27880 0 27936 800
rect 28340 0 28396 800
rect 28892 0 28948 800
rect 29352 0 29408 800
rect 29812 0 29868 800
rect 30364 0 30420 800
rect 30824 0 30880 800
rect 31284 0 31340 800
rect 31836 0 31892 800
rect 32296 0 32352 800
rect 32756 0 32812 800
rect 33308 0 33364 800
rect 33768 0 33824 800
rect 34228 0 34284 800
rect 34780 0 34836 800
rect 35240 0 35296 800
rect 35700 0 35756 800
rect 36252 0 36308 800
rect 36712 0 36768 800
rect 37172 0 37228 800
rect 37632 0 37688 800
rect 38184 0 38240 800
rect 38644 0 38700 800
rect 39104 0 39160 800
rect 39656 0 39712 800
rect 40116 0 40172 800
rect 40576 0 40632 800
rect 41128 0 41184 800
rect 41588 0 41644 800
rect 42048 0 42104 800
rect 42600 0 42656 800
rect 43060 0 43116 800
rect 43520 0 43576 800
rect 44072 0 44128 800
rect 44532 0 44588 800
rect 44992 0 45048 800
rect 45544 0 45600 800
rect 46004 0 46060 800
rect 46464 0 46520 800
rect 47016 0 47072 800
rect 47476 0 47532 800
rect 47936 0 47992 800
rect 48488 0 48544 800
rect 48948 0 49004 800
rect 49408 0 49464 800
rect 49960 0 50016 800
rect 50420 0 50476 800
rect 50880 0 50936 800
rect 51432 0 51488 800
rect 51892 0 51948 800
rect 52352 0 52408 800
rect 52904 0 52960 800
rect 53364 0 53420 800
rect 53824 0 53880 800
rect 54376 0 54432 800
rect 54836 0 54892 800
rect 55296 0 55352 800
rect 55756 0 55812 800
rect 56308 0 56364 800
rect 56768 0 56824 800
rect 57228 0 57284 800
rect 57780 0 57836 800
rect 58240 0 58296 800
rect 58700 0 58756 800
rect 59252 0 59308 800
rect 59712 0 59768 800
rect 60172 0 60228 800
rect 60724 0 60780 800
rect 61184 0 61240 800
rect 61644 0 61700 800
rect 62196 0 62252 800
rect 62656 0 62712 800
rect 63116 0 63172 800
rect 63668 0 63724 800
rect 64128 0 64184 800
rect 64588 0 64644 800
rect 65140 0 65196 800
rect 65600 0 65656 800
rect 66060 0 66116 800
rect 66612 0 66668 800
rect 67072 0 67128 800
rect 67532 0 67588 800
rect 68084 0 68140 800
rect 68544 0 68600 800
rect 69004 0 69060 800
rect 69556 0 69612 800
rect 70016 0 70072 800
rect 70476 0 70532 800
rect 71028 0 71084 800
rect 71488 0 71544 800
rect 71948 0 72004 800
rect 72500 0 72556 800
rect 72960 0 73016 800
rect 73420 0 73476 800
rect 73880 0 73936 800
rect 74432 0 74488 800
rect 74892 0 74948 800
rect 75352 0 75408 800
rect 75904 0 75960 800
rect 76364 0 76420 800
rect 76824 0 76880 800
rect 77376 0 77432 800
rect 77836 0 77892 800
rect 78296 0 78352 800
rect 78848 0 78904 800
rect 79308 0 79364 800
rect 79768 0 79824 800
rect 80320 0 80376 800
rect 80780 0 80836 800
rect 81240 0 81296 800
rect 81792 0 81848 800
rect 82252 0 82308 800
rect 82712 0 82768 800
rect 83264 0 83320 800
rect 83724 0 83780 800
rect 84184 0 84240 800
rect 84736 0 84792 800
rect 85196 0 85252 800
rect 85656 0 85712 800
rect 86208 0 86264 800
rect 86668 0 86724 800
rect 87128 0 87184 800
rect 87680 0 87736 800
rect 88140 0 88196 800
rect 88600 0 88656 800
rect 89152 0 89208 800
rect 89612 0 89668 800
rect 90072 0 90128 800
rect 90624 0 90680 800
rect 91084 0 91140 800
rect 91544 0 91600 800
rect 92096 0 92152 800
rect 92556 0 92612 800
rect 93016 0 93072 800
rect 93476 0 93532 800
rect 94028 0 94084 800
rect 94488 0 94544 800
rect 94948 0 95004 800
rect 95500 0 95556 800
rect 95960 0 96016 800
rect 96420 0 96476 800
rect 96972 0 97028 800
rect 97432 0 97488 800
rect 97892 0 97948 800
rect 98444 0 98500 800
rect 98904 0 98960 800
rect 99364 0 99420 800
rect 99916 0 99972 800
rect 100376 0 100432 800
rect 100836 0 100892 800
rect 101388 0 101444 800
rect 101848 0 101904 800
rect 102308 0 102364 800
rect 102860 0 102916 800
rect 103320 0 103376 800
rect 103780 0 103836 800
rect 104332 0 104388 800
rect 104792 0 104848 800
rect 105252 0 105308 800
rect 105804 0 105860 800
rect 106264 0 106320 800
rect 106724 0 106780 800
rect 107276 0 107332 800
rect 107736 0 107792 800
rect 108196 0 108252 800
rect 108748 0 108804 800
rect 109208 0 109264 800
rect 109668 0 109724 800
rect 110220 0 110276 800
rect 110680 0 110736 800
rect 111140 0 111196 800
rect 111600 0 111656 800
rect 112152 0 112208 800
rect 112612 0 112668 800
rect 113072 0 113128 800
rect 113624 0 113680 800
rect 114084 0 114140 800
rect 114544 0 114600 800
rect 115096 0 115152 800
rect 115556 0 115612 800
rect 116016 0 116072 800
rect 116568 0 116624 800
rect 117028 0 117084 800
rect 117488 0 117544 800
rect 118040 0 118096 800
rect 118500 0 118556 800
rect 118960 0 119016 800
rect 119512 0 119568 800
rect 119972 0 120028 800
rect 120432 0 120488 800
rect 120984 0 121040 800
rect 121444 0 121500 800
rect 121904 0 121960 800
rect 122456 0 122512 800
rect 122916 0 122972 800
rect 123376 0 123432 800
rect 123928 0 123984 800
rect 124388 0 124444 800
rect 124848 0 124904 800
rect 125400 0 125456 800
rect 125860 0 125916 800
rect 126320 0 126376 800
rect 126872 0 126928 800
rect 127332 0 127388 800
rect 127792 0 127848 800
rect 128344 0 128400 800
rect 128804 0 128860 800
rect 129264 0 129320 800
rect 129724 0 129780 800
rect 130276 0 130332 800
rect 130736 0 130792 800
rect 131196 0 131252 800
rect 131748 0 131804 800
rect 132208 0 132264 800
rect 132668 0 132724 800
rect 133220 0 133276 800
rect 133680 0 133736 800
rect 134140 0 134196 800
rect 134692 0 134748 800
rect 135152 0 135208 800
rect 135612 0 135668 800
rect 136164 0 136220 800
rect 136624 0 136680 800
rect 137084 0 137140 800
rect 137636 0 137692 800
rect 138096 0 138152 800
rect 138556 0 138612 800
rect 139108 0 139164 800
rect 139568 0 139624 800
rect 140028 0 140084 800
rect 140580 0 140636 800
rect 141040 0 141096 800
rect 141500 0 141556 800
rect 142052 0 142108 800
rect 142512 0 142568 800
rect 142972 0 143028 800
rect 143524 0 143580 800
rect 143984 0 144040 800
rect 144444 0 144500 800
rect 144996 0 145052 800
rect 145456 0 145512 800
rect 145916 0 145972 800
rect 146468 0 146524 800
rect 146928 0 146984 800
rect 147388 0 147444 800
rect 147848 0 147904 800
rect 148400 0 148456 800
rect 148860 0 148916 800
rect 149320 0 149376 800
rect 149872 0 149928 800
rect 150332 0 150388 800
rect 150792 0 150848 800
rect 151344 0 151400 800
rect 151804 0 151860 800
rect 152264 0 152320 800
rect 152816 0 152872 800
rect 153276 0 153332 800
rect 153736 0 153792 800
rect 154288 0 154344 800
rect 154748 0 154804 800
rect 155208 0 155264 800
rect 155760 0 155816 800
rect 156220 0 156276 800
rect 156680 0 156736 800
rect 157232 0 157288 800
rect 157692 0 157748 800
rect 158152 0 158208 800
rect 158704 0 158760 800
rect 159164 0 159220 800
rect 159624 0 159680 800
rect 160176 0 160232 800
rect 160636 0 160692 800
rect 161096 0 161152 800
rect 161648 0 161704 800
rect 162108 0 162164 800
rect 162568 0 162624 800
rect 163120 0 163176 800
rect 163580 0 163636 800
rect 164040 0 164096 800
rect 164592 0 164648 800
rect 165052 0 165108 800
rect 165512 0 165568 800
rect 166064 0 166120 800
rect 166524 0 166580 800
rect 166984 0 167040 800
rect 167444 0 167500 800
rect 167996 0 168052 800
rect 168456 0 168512 800
rect 168916 0 168972 800
rect 169468 0 169524 800
rect 169928 0 169984 800
rect 170388 0 170444 800
rect 170940 0 170996 800
rect 171400 0 171456 800
rect 171860 0 171916 800
rect 172412 0 172468 800
rect 172872 0 172928 800
rect 173332 0 173388 800
rect 173884 0 173940 800
rect 174344 0 174400 800
rect 174804 0 174860 800
rect 175356 0 175412 800
rect 175816 0 175872 800
rect 176276 0 176332 800
rect 176828 0 176884 800
rect 177288 0 177344 800
rect 177748 0 177804 800
rect 178300 0 178356 800
rect 178760 0 178816 800
rect 179220 0 179276 800
rect 179772 0 179828 800
rect 180232 0 180288 800
rect 180692 0 180748 800
rect 181244 0 181300 800
rect 181704 0 181760 800
rect 182164 0 182220 800
rect 182716 0 182772 800
rect 183176 0 183232 800
rect 183636 0 183692 800
rect 184188 0 184244 800
rect 184648 0 184704 800
rect 185108 0 185164 800
rect 185568 0 185624 800
rect 186120 0 186176 800
rect 186580 0 186636 800
rect 187040 0 187096 800
rect 187592 0 187648 800
rect 188052 0 188108 800
rect 188512 0 188568 800
rect 189064 0 189120 800
rect 189524 0 189580 800
rect 189984 0 190040 800
rect 190536 0 190592 800
rect 190996 0 191052 800
rect 191456 0 191512 800
rect 192008 0 192064 800
rect 192468 0 192524 800
rect 192928 0 192984 800
rect 193480 0 193536 800
rect 193940 0 193996 800
rect 194400 0 194456 800
rect 194952 0 195008 800
rect 195412 0 195468 800
rect 195872 0 195928 800
rect 196424 0 196480 800
rect 196884 0 196940 800
rect 197344 0 197400 800
rect 197896 0 197952 800
rect 198356 0 198412 800
rect 198816 0 198872 800
rect 199368 0 199424 800
rect 199828 0 199884 800
rect 200288 0 200344 800
rect 200840 0 200896 800
rect 201300 0 201356 800
rect 201760 0 201816 800
rect 202312 0 202368 800
rect 202772 0 202828 800
rect 203232 0 203288 800
rect 203692 0 203748 800
rect 204244 0 204300 800
rect 204704 0 204760 800
rect 205164 0 205220 800
rect 205716 0 205772 800
rect 206176 0 206232 800
rect 206636 0 206692 800
rect 207188 0 207244 800
rect 207648 0 207704 800
rect 208108 0 208164 800
rect 208660 0 208716 800
rect 209120 0 209176 800
rect 209580 0 209636 800
rect 210132 0 210188 800
rect 210592 0 210648 800
rect 211052 0 211108 800
rect 211604 0 211660 800
rect 212064 0 212120 800
rect 212524 0 212580 800
rect 213076 0 213132 800
rect 213536 0 213592 800
rect 213996 0 214052 800
rect 214548 0 214604 800
rect 215008 0 215064 800
rect 215468 0 215524 800
rect 216020 0 216076 800
rect 216480 0 216536 800
rect 216940 0 216996 800
rect 217492 0 217548 800
rect 217952 0 218008 800
rect 218412 0 218468 800
rect 218964 0 219020 800
rect 219424 0 219480 800
rect 219884 0 219940 800
rect 220436 0 220492 800
rect 220896 0 220952 800
rect 221356 0 221412 800
rect 221816 0 221872 800
rect 222368 0 222424 800
rect 222828 0 222884 800
rect 223288 0 223344 800
rect 223840 0 223896 800
rect 224300 0 224356 800
rect 224760 0 224816 800
rect 225312 0 225368 800
rect 225772 0 225828 800
rect 226232 0 226288 800
rect 226784 0 226840 800
rect 227244 0 227300 800
rect 227704 0 227760 800
rect 228256 0 228312 800
rect 228716 0 228772 800
rect 229176 0 229232 800
rect 229728 0 229784 800
rect 230188 0 230244 800
rect 230648 0 230704 800
rect 231200 0 231256 800
rect 231660 0 231716 800
rect 232120 0 232176 800
rect 232672 0 232728 800
rect 233132 0 233188 800
rect 233592 0 233648 800
rect 234144 0 234200 800
rect 234604 0 234660 800
rect 235064 0 235120 800
rect 235616 0 235672 800
rect 236076 0 236132 800
rect 236536 0 236592 800
rect 237088 0 237144 800
rect 237548 0 237604 800
rect 238008 0 238064 800
rect 238560 0 238616 800
rect 239020 0 239076 800
rect 239480 0 239536 800
<< obsm2 >>
rect 6 239144 776 239200
rect 944 239144 2800 239200
rect 2968 239144 4916 239200
rect 5084 239144 7032 239200
rect 7200 239144 9148 239200
rect 9316 239144 11264 239200
rect 11432 239144 13380 239200
rect 13548 239144 15496 239200
rect 15664 239144 17612 239200
rect 17780 239144 19636 239200
rect 19804 239144 21752 239200
rect 21920 239144 23868 239200
rect 24036 239144 25984 239200
rect 26152 239144 28100 239200
rect 28268 239144 30216 239200
rect 30384 239144 32332 239200
rect 32500 239144 34448 239200
rect 34616 239144 36564 239200
rect 36732 239144 38588 239200
rect 38756 239144 40704 239200
rect 40872 239144 42820 239200
rect 42988 239144 44936 239200
rect 45104 239144 47052 239200
rect 47220 239144 49168 239200
rect 49336 239144 51284 239200
rect 51452 239144 53400 239200
rect 53568 239144 55516 239200
rect 55684 239144 57540 239200
rect 57708 239144 59656 239200
rect 59824 239144 61772 239200
rect 61940 239144 63888 239200
rect 64056 239144 66004 239200
rect 66172 239144 68120 239200
rect 68288 239144 70236 239200
rect 70404 239144 72352 239200
rect 72520 239144 74468 239200
rect 74636 239144 76492 239200
rect 76660 239144 78608 239200
rect 78776 239144 80724 239200
rect 80892 239144 82840 239200
rect 83008 239144 84956 239200
rect 85124 239144 87072 239200
rect 87240 239144 89188 239200
rect 89356 239144 91304 239200
rect 91472 239144 93328 239200
rect 93496 239144 95444 239200
rect 95612 239144 97560 239200
rect 97728 239144 99676 239200
rect 99844 239144 101792 239200
rect 101960 239144 103908 239200
rect 104076 239144 106024 239200
rect 106192 239144 108140 239200
rect 108308 239144 110256 239200
rect 110424 239144 112280 239200
rect 112448 239144 114396 239200
rect 114564 239144 116512 239200
rect 116680 239144 118628 239200
rect 118796 239144 120744 239200
rect 120912 239144 122860 239200
rect 123028 239144 124976 239200
rect 125144 239144 127092 239200
rect 127260 239144 129208 239200
rect 129376 239144 131232 239200
rect 131400 239144 133348 239200
rect 133516 239144 135464 239200
rect 135632 239144 137580 239200
rect 137748 239144 139696 239200
rect 139864 239144 141812 239200
rect 141980 239144 143928 239200
rect 144096 239144 146044 239200
rect 146212 239144 148160 239200
rect 148328 239144 150184 239200
rect 150352 239144 152300 239200
rect 152468 239144 154416 239200
rect 154584 239144 156532 239200
rect 156700 239144 158648 239200
rect 158816 239144 160764 239200
rect 160932 239144 162880 239200
rect 163048 239144 164996 239200
rect 165164 239144 167020 239200
rect 167188 239144 169136 239200
rect 169304 239144 171252 239200
rect 171420 239144 173368 239200
rect 173536 239144 175484 239200
rect 175652 239144 177600 239200
rect 177768 239144 179716 239200
rect 179884 239144 181832 239200
rect 182000 239144 183948 239200
rect 184116 239144 185972 239200
rect 186140 239144 188088 239200
rect 188256 239144 190204 239200
rect 190372 239144 192320 239200
rect 192488 239144 194436 239200
rect 194604 239144 196552 239200
rect 196720 239144 198668 239200
rect 198836 239144 200784 239200
rect 200952 239144 202900 239200
rect 203068 239144 204924 239200
rect 205092 239144 207040 239200
rect 207208 239144 209156 239200
rect 209324 239144 211272 239200
rect 211440 239144 213388 239200
rect 213556 239144 215504 239200
rect 215672 239144 217620 239200
rect 217788 239144 219736 239200
rect 219904 239144 221852 239200
rect 222020 239144 223876 239200
rect 224044 239144 225992 239200
rect 226160 239144 228108 239200
rect 228276 239144 230224 239200
rect 230392 239144 232340 239200
rect 232508 239144 234456 239200
rect 234624 239144 236572 239200
rect 236740 239144 238688 239200
rect 238856 239144 239534 239200
rect 6 856 239534 239144
rect 116 800 408 856
rect 576 800 868 856
rect 1036 800 1328 856
rect 1496 800 1880 856
rect 2048 800 2340 856
rect 2508 800 2800 856
rect 2968 800 3352 856
rect 3520 800 3812 856
rect 3980 800 4272 856
rect 4440 800 4824 856
rect 4992 800 5284 856
rect 5452 800 5744 856
rect 5912 800 6296 856
rect 6464 800 6756 856
rect 6924 800 7216 856
rect 7384 800 7768 856
rect 7936 800 8228 856
rect 8396 800 8688 856
rect 8856 800 9240 856
rect 9408 800 9700 856
rect 9868 800 10160 856
rect 10328 800 10712 856
rect 10880 800 11172 856
rect 11340 800 11632 856
rect 11800 800 12184 856
rect 12352 800 12644 856
rect 12812 800 13104 856
rect 13272 800 13656 856
rect 13824 800 14116 856
rect 14284 800 14576 856
rect 14744 800 15128 856
rect 15296 800 15588 856
rect 15756 800 16048 856
rect 16216 800 16600 856
rect 16768 800 17060 856
rect 17228 800 17520 856
rect 17688 800 18072 856
rect 18240 800 18532 856
rect 18700 800 18992 856
rect 19160 800 19452 856
rect 19620 800 20004 856
rect 20172 800 20464 856
rect 20632 800 20924 856
rect 21092 800 21476 856
rect 21644 800 21936 856
rect 22104 800 22396 856
rect 22564 800 22948 856
rect 23116 800 23408 856
rect 23576 800 23868 856
rect 24036 800 24420 856
rect 24588 800 24880 856
rect 25048 800 25340 856
rect 25508 800 25892 856
rect 26060 800 26352 856
rect 26520 800 26812 856
rect 26980 800 27364 856
rect 27532 800 27824 856
rect 27992 800 28284 856
rect 28452 800 28836 856
rect 29004 800 29296 856
rect 29464 800 29756 856
rect 29924 800 30308 856
rect 30476 800 30768 856
rect 30936 800 31228 856
rect 31396 800 31780 856
rect 31948 800 32240 856
rect 32408 800 32700 856
rect 32868 800 33252 856
rect 33420 800 33712 856
rect 33880 800 34172 856
rect 34340 800 34724 856
rect 34892 800 35184 856
rect 35352 800 35644 856
rect 35812 800 36196 856
rect 36364 800 36656 856
rect 36824 800 37116 856
rect 37284 800 37576 856
rect 37744 800 38128 856
rect 38296 800 38588 856
rect 38756 800 39048 856
rect 39216 800 39600 856
rect 39768 800 40060 856
rect 40228 800 40520 856
rect 40688 800 41072 856
rect 41240 800 41532 856
rect 41700 800 41992 856
rect 42160 800 42544 856
rect 42712 800 43004 856
rect 43172 800 43464 856
rect 43632 800 44016 856
rect 44184 800 44476 856
rect 44644 800 44936 856
rect 45104 800 45488 856
rect 45656 800 45948 856
rect 46116 800 46408 856
rect 46576 800 46960 856
rect 47128 800 47420 856
rect 47588 800 47880 856
rect 48048 800 48432 856
rect 48600 800 48892 856
rect 49060 800 49352 856
rect 49520 800 49904 856
rect 50072 800 50364 856
rect 50532 800 50824 856
rect 50992 800 51376 856
rect 51544 800 51836 856
rect 52004 800 52296 856
rect 52464 800 52848 856
rect 53016 800 53308 856
rect 53476 800 53768 856
rect 53936 800 54320 856
rect 54488 800 54780 856
rect 54948 800 55240 856
rect 55408 800 55700 856
rect 55868 800 56252 856
rect 56420 800 56712 856
rect 56880 800 57172 856
rect 57340 800 57724 856
rect 57892 800 58184 856
rect 58352 800 58644 856
rect 58812 800 59196 856
rect 59364 800 59656 856
rect 59824 800 60116 856
rect 60284 800 60668 856
rect 60836 800 61128 856
rect 61296 800 61588 856
rect 61756 800 62140 856
rect 62308 800 62600 856
rect 62768 800 63060 856
rect 63228 800 63612 856
rect 63780 800 64072 856
rect 64240 800 64532 856
rect 64700 800 65084 856
rect 65252 800 65544 856
rect 65712 800 66004 856
rect 66172 800 66556 856
rect 66724 800 67016 856
rect 67184 800 67476 856
rect 67644 800 68028 856
rect 68196 800 68488 856
rect 68656 800 68948 856
rect 69116 800 69500 856
rect 69668 800 69960 856
rect 70128 800 70420 856
rect 70588 800 70972 856
rect 71140 800 71432 856
rect 71600 800 71892 856
rect 72060 800 72444 856
rect 72612 800 72904 856
rect 73072 800 73364 856
rect 73532 800 73824 856
rect 73992 800 74376 856
rect 74544 800 74836 856
rect 75004 800 75296 856
rect 75464 800 75848 856
rect 76016 800 76308 856
rect 76476 800 76768 856
rect 76936 800 77320 856
rect 77488 800 77780 856
rect 77948 800 78240 856
rect 78408 800 78792 856
rect 78960 800 79252 856
rect 79420 800 79712 856
rect 79880 800 80264 856
rect 80432 800 80724 856
rect 80892 800 81184 856
rect 81352 800 81736 856
rect 81904 800 82196 856
rect 82364 800 82656 856
rect 82824 800 83208 856
rect 83376 800 83668 856
rect 83836 800 84128 856
rect 84296 800 84680 856
rect 84848 800 85140 856
rect 85308 800 85600 856
rect 85768 800 86152 856
rect 86320 800 86612 856
rect 86780 800 87072 856
rect 87240 800 87624 856
rect 87792 800 88084 856
rect 88252 800 88544 856
rect 88712 800 89096 856
rect 89264 800 89556 856
rect 89724 800 90016 856
rect 90184 800 90568 856
rect 90736 800 91028 856
rect 91196 800 91488 856
rect 91656 800 92040 856
rect 92208 800 92500 856
rect 92668 800 92960 856
rect 93128 800 93420 856
rect 93588 800 93972 856
rect 94140 800 94432 856
rect 94600 800 94892 856
rect 95060 800 95444 856
rect 95612 800 95904 856
rect 96072 800 96364 856
rect 96532 800 96916 856
rect 97084 800 97376 856
rect 97544 800 97836 856
rect 98004 800 98388 856
rect 98556 800 98848 856
rect 99016 800 99308 856
rect 99476 800 99860 856
rect 100028 800 100320 856
rect 100488 800 100780 856
rect 100948 800 101332 856
rect 101500 800 101792 856
rect 101960 800 102252 856
rect 102420 800 102804 856
rect 102972 800 103264 856
rect 103432 800 103724 856
rect 103892 800 104276 856
rect 104444 800 104736 856
rect 104904 800 105196 856
rect 105364 800 105748 856
rect 105916 800 106208 856
rect 106376 800 106668 856
rect 106836 800 107220 856
rect 107388 800 107680 856
rect 107848 800 108140 856
rect 108308 800 108692 856
rect 108860 800 109152 856
rect 109320 800 109612 856
rect 109780 800 110164 856
rect 110332 800 110624 856
rect 110792 800 111084 856
rect 111252 800 111544 856
rect 111712 800 112096 856
rect 112264 800 112556 856
rect 112724 800 113016 856
rect 113184 800 113568 856
rect 113736 800 114028 856
rect 114196 800 114488 856
rect 114656 800 115040 856
rect 115208 800 115500 856
rect 115668 800 115960 856
rect 116128 800 116512 856
rect 116680 800 116972 856
rect 117140 800 117432 856
rect 117600 800 117984 856
rect 118152 800 118444 856
rect 118612 800 118904 856
rect 119072 800 119456 856
rect 119624 800 119916 856
rect 120084 800 120376 856
rect 120544 800 120928 856
rect 121096 800 121388 856
rect 121556 800 121848 856
rect 122016 800 122400 856
rect 122568 800 122860 856
rect 123028 800 123320 856
rect 123488 800 123872 856
rect 124040 800 124332 856
rect 124500 800 124792 856
rect 124960 800 125344 856
rect 125512 800 125804 856
rect 125972 800 126264 856
rect 126432 800 126816 856
rect 126984 800 127276 856
rect 127444 800 127736 856
rect 127904 800 128288 856
rect 128456 800 128748 856
rect 128916 800 129208 856
rect 129376 800 129668 856
rect 129836 800 130220 856
rect 130388 800 130680 856
rect 130848 800 131140 856
rect 131308 800 131692 856
rect 131860 800 132152 856
rect 132320 800 132612 856
rect 132780 800 133164 856
rect 133332 800 133624 856
rect 133792 800 134084 856
rect 134252 800 134636 856
rect 134804 800 135096 856
rect 135264 800 135556 856
rect 135724 800 136108 856
rect 136276 800 136568 856
rect 136736 800 137028 856
rect 137196 800 137580 856
rect 137748 800 138040 856
rect 138208 800 138500 856
rect 138668 800 139052 856
rect 139220 800 139512 856
rect 139680 800 139972 856
rect 140140 800 140524 856
rect 140692 800 140984 856
rect 141152 800 141444 856
rect 141612 800 141996 856
rect 142164 800 142456 856
rect 142624 800 142916 856
rect 143084 800 143468 856
rect 143636 800 143928 856
rect 144096 800 144388 856
rect 144556 800 144940 856
rect 145108 800 145400 856
rect 145568 800 145860 856
rect 146028 800 146412 856
rect 146580 800 146872 856
rect 147040 800 147332 856
rect 147500 800 147792 856
rect 147960 800 148344 856
rect 148512 800 148804 856
rect 148972 800 149264 856
rect 149432 800 149816 856
rect 149984 800 150276 856
rect 150444 800 150736 856
rect 150904 800 151288 856
rect 151456 800 151748 856
rect 151916 800 152208 856
rect 152376 800 152760 856
rect 152928 800 153220 856
rect 153388 800 153680 856
rect 153848 800 154232 856
rect 154400 800 154692 856
rect 154860 800 155152 856
rect 155320 800 155704 856
rect 155872 800 156164 856
rect 156332 800 156624 856
rect 156792 800 157176 856
rect 157344 800 157636 856
rect 157804 800 158096 856
rect 158264 800 158648 856
rect 158816 800 159108 856
rect 159276 800 159568 856
rect 159736 800 160120 856
rect 160288 800 160580 856
rect 160748 800 161040 856
rect 161208 800 161592 856
rect 161760 800 162052 856
rect 162220 800 162512 856
rect 162680 800 163064 856
rect 163232 800 163524 856
rect 163692 800 163984 856
rect 164152 800 164536 856
rect 164704 800 164996 856
rect 165164 800 165456 856
rect 165624 800 166008 856
rect 166176 800 166468 856
rect 166636 800 166928 856
rect 167096 800 167388 856
rect 167556 800 167940 856
rect 168108 800 168400 856
rect 168568 800 168860 856
rect 169028 800 169412 856
rect 169580 800 169872 856
rect 170040 800 170332 856
rect 170500 800 170884 856
rect 171052 800 171344 856
rect 171512 800 171804 856
rect 171972 800 172356 856
rect 172524 800 172816 856
rect 172984 800 173276 856
rect 173444 800 173828 856
rect 173996 800 174288 856
rect 174456 800 174748 856
rect 174916 800 175300 856
rect 175468 800 175760 856
rect 175928 800 176220 856
rect 176388 800 176772 856
rect 176940 800 177232 856
rect 177400 800 177692 856
rect 177860 800 178244 856
rect 178412 800 178704 856
rect 178872 800 179164 856
rect 179332 800 179716 856
rect 179884 800 180176 856
rect 180344 800 180636 856
rect 180804 800 181188 856
rect 181356 800 181648 856
rect 181816 800 182108 856
rect 182276 800 182660 856
rect 182828 800 183120 856
rect 183288 800 183580 856
rect 183748 800 184132 856
rect 184300 800 184592 856
rect 184760 800 185052 856
rect 185220 800 185512 856
rect 185680 800 186064 856
rect 186232 800 186524 856
rect 186692 800 186984 856
rect 187152 800 187536 856
rect 187704 800 187996 856
rect 188164 800 188456 856
rect 188624 800 189008 856
rect 189176 800 189468 856
rect 189636 800 189928 856
rect 190096 800 190480 856
rect 190648 800 190940 856
rect 191108 800 191400 856
rect 191568 800 191952 856
rect 192120 800 192412 856
rect 192580 800 192872 856
rect 193040 800 193424 856
rect 193592 800 193884 856
rect 194052 800 194344 856
rect 194512 800 194896 856
rect 195064 800 195356 856
rect 195524 800 195816 856
rect 195984 800 196368 856
rect 196536 800 196828 856
rect 196996 800 197288 856
rect 197456 800 197840 856
rect 198008 800 198300 856
rect 198468 800 198760 856
rect 198928 800 199312 856
rect 199480 800 199772 856
rect 199940 800 200232 856
rect 200400 800 200784 856
rect 200952 800 201244 856
rect 201412 800 201704 856
rect 201872 800 202256 856
rect 202424 800 202716 856
rect 202884 800 203176 856
rect 203344 800 203636 856
rect 203804 800 204188 856
rect 204356 800 204648 856
rect 204816 800 205108 856
rect 205276 800 205660 856
rect 205828 800 206120 856
rect 206288 800 206580 856
rect 206748 800 207132 856
rect 207300 800 207592 856
rect 207760 800 208052 856
rect 208220 800 208604 856
rect 208772 800 209064 856
rect 209232 800 209524 856
rect 209692 800 210076 856
rect 210244 800 210536 856
rect 210704 800 210996 856
rect 211164 800 211548 856
rect 211716 800 212008 856
rect 212176 800 212468 856
rect 212636 800 213020 856
rect 213188 800 213480 856
rect 213648 800 213940 856
rect 214108 800 214492 856
rect 214660 800 214952 856
rect 215120 800 215412 856
rect 215580 800 215964 856
rect 216132 800 216424 856
rect 216592 800 216884 856
rect 217052 800 217436 856
rect 217604 800 217896 856
rect 218064 800 218356 856
rect 218524 800 218908 856
rect 219076 800 219368 856
rect 219536 800 219828 856
rect 219996 800 220380 856
rect 220548 800 220840 856
rect 221008 800 221300 856
rect 221468 800 221760 856
rect 221928 800 222312 856
rect 222480 800 222772 856
rect 222940 800 223232 856
rect 223400 800 223784 856
rect 223952 800 224244 856
rect 224412 800 224704 856
rect 224872 800 225256 856
rect 225424 800 225716 856
rect 225884 800 226176 856
rect 226344 800 226728 856
rect 226896 800 227188 856
rect 227356 800 227648 856
rect 227816 800 228200 856
rect 228368 800 228660 856
rect 228828 800 229120 856
rect 229288 800 229672 856
rect 229840 800 230132 856
rect 230300 800 230592 856
rect 230760 800 231144 856
rect 231312 800 231604 856
rect 231772 800 232064 856
rect 232232 800 232616 856
rect 232784 800 233076 856
rect 233244 800 233536 856
rect 233704 800 234088 856
rect 234256 800 234548 856
rect 234716 800 235008 856
rect 235176 800 235560 856
rect 235728 800 236020 856
rect 236188 800 236480 856
rect 236648 800 237032 856
rect 237200 800 237492 856
rect 237660 800 237952 856
rect 238120 800 238504 856
rect 238672 800 238964 856
rect 239132 800 239424 856
<< obsm3 >>
rect 459 851 236781 237761
<< metal4 >>
rect 4010 2128 4330 237776
rect 19370 2128 19690 237776
rect 34730 2128 35050 237776
rect 50090 2128 50410 237776
rect 65450 2128 65770 237776
rect 80810 2128 81130 237776
rect 96170 2128 96490 237776
rect 111530 2128 111850 237776
rect 126890 2128 127210 237776
rect 142250 2128 142570 237776
rect 157610 2128 157930 237776
rect 172970 2128 173290 237776
rect 188330 2128 188650 237776
rect 203690 2128 204010 237776
rect 219050 2128 219370 237776
rect 234410 2128 234730 237776
<< obsm4 >>
rect 13477 12139 19290 232933
rect 19770 12139 34650 232933
rect 35130 12139 50010 232933
rect 50490 12139 65370 232933
rect 65850 12139 80730 232933
rect 81210 12139 96090 232933
rect 96570 12139 111450 232933
rect 111930 12139 126810 232933
rect 127290 12139 142170 232933
rect 142650 12139 157530 232933
rect 158010 12139 172890 232933
rect 173370 12139 188250 232933
rect 188730 12139 203610 232933
rect 204090 12139 218970 232933
rect 219450 12139 233975 232933
<< labels >>
rlabel metal2 s 832 239200 888 240000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 63944 239200 64000 240000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 70292 239200 70348 240000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 76548 239200 76604 240000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 82896 239200 82952 240000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 89244 239200 89300 240000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 95500 239200 95556 240000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 101848 239200 101904 240000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 108196 239200 108252 240000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 114452 239200 114508 240000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 120800 239200 120856 240000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 7088 239200 7144 240000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 127148 239200 127204 240000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 133404 239200 133460 240000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 139752 239200 139808 240000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 146100 239200 146156 240000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 152356 239200 152412 240000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 158704 239200 158760 240000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 165052 239200 165108 240000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 171308 239200 171364 240000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 177656 239200 177712 240000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 184004 239200 184060 240000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 13436 239200 13492 240000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 190260 239200 190316 240000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 196608 239200 196664 240000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 202956 239200 203012 240000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 209212 239200 209268 240000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 215560 239200 215616 240000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 221908 239200 221964 240000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 228164 239200 228220 240000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 234512 239200 234568 240000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 19692 239200 19748 240000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 26040 239200 26096 240000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 32388 239200 32444 240000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 38644 239200 38700 240000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 44992 239200 45048 240000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 51340 239200 51396 240000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 57596 239200 57652 240000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2856 239200 2912 240000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 66060 239200 66116 240000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 72408 239200 72464 240000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 78664 239200 78720 240000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 85012 239200 85068 240000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 91360 239200 91416 240000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 97616 239200 97672 240000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 103964 239200 104020 240000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 110312 239200 110368 240000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 116568 239200 116624 240000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 122916 239200 122972 240000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 9204 239200 9260 240000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 129264 239200 129320 240000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 135520 239200 135576 240000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 141868 239200 141924 240000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 148216 239200 148272 240000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 154472 239200 154528 240000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 160820 239200 160876 240000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 167076 239200 167132 240000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 173424 239200 173480 240000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 179772 239200 179828 240000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 186028 239200 186084 240000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 15552 239200 15608 240000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 192376 239200 192432 240000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 198724 239200 198780 240000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 204980 239200 205036 240000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 211328 239200 211384 240000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 217676 239200 217732 240000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 223932 239200 223988 240000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 230280 239200 230336 240000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 236628 239200 236684 240000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 21808 239200 21864 240000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 28156 239200 28212 240000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 34504 239200 34560 240000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 40760 239200 40816 240000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 47108 239200 47164 240000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 53456 239200 53512 240000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 59712 239200 59768 240000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 4972 239200 5028 240000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 68176 239200 68232 240000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 74524 239200 74580 240000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 80780 239200 80836 240000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 87128 239200 87184 240000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 93384 239200 93440 240000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 99732 239200 99788 240000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 106080 239200 106136 240000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 112336 239200 112392 240000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 118684 239200 118740 240000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 125032 239200 125088 240000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 11320 239200 11376 240000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 131288 239200 131344 240000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 137636 239200 137692 240000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 143984 239200 144040 240000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 150240 239200 150296 240000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 156588 239200 156644 240000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 162936 239200 162992 240000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 169192 239200 169248 240000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 175540 239200 175596 240000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 181888 239200 181944 240000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 188144 239200 188200 240000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 17668 239200 17724 240000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 194492 239200 194548 240000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 200840 239200 200896 240000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 207096 239200 207152 240000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 213444 239200 213500 240000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 219792 239200 219848 240000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 226048 239200 226104 240000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 232396 239200 232452 240000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 238744 239200 238800 240000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 23924 239200 23980 240000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 30272 239200 30328 240000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 36620 239200 36676 240000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 42876 239200 42932 240000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 49224 239200 49280 240000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 55572 239200 55628 240000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 61828 239200 61884 240000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 51892 0 51948 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 198816 0 198872 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 200288 0 200344 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 201760 0 201816 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 203232 0 203288 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 204704 0 204760 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 206176 0 206232 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 207648 0 207704 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 209120 0 209176 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 210592 0 210648 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 212064 0 212120 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 66612 0 66668 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 213536 0 213592 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 215008 0 215064 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 216480 0 216536 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 217952 0 218008 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 219424 0 219480 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 220896 0 220952 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 222368 0 222424 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 223840 0 223896 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 225312 0 225368 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 226784 0 226840 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 68084 0 68140 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 228256 0 228312 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 229728 0 229784 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 231200 0 231256 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 232672 0 232728 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 234144 0 234200 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 235616 0 235672 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 237088 0 237144 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 238560 0 238616 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 69556 0 69612 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 71028 0 71084 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 72500 0 72556 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 73880 0 73936 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 75352 0 75408 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 76824 0 76880 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 78296 0 78352 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 79768 0 79824 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 53364 0 53420 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 81240 0 81296 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 82712 0 82768 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 84184 0 84240 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 85656 0 85712 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 87128 0 87184 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 88600 0 88656 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 90072 0 90128 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 91544 0 91600 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 93016 0 93072 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 94488 0 94544 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 54836 0 54892 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 95960 0 96016 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 97432 0 97488 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 98904 0 98960 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 100376 0 100432 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 101848 0 101904 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 103320 0 103376 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 104792 0 104848 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 106264 0 106320 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 107736 0 107792 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 109208 0 109264 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 56308 0 56364 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 110680 0 110736 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 112152 0 112208 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 113624 0 113680 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 115096 0 115152 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 116568 0 116624 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 118040 0 118096 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 119512 0 119568 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 120984 0 121040 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 122456 0 122512 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 123928 0 123984 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 57780 0 57836 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 125400 0 125456 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 126872 0 126928 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 128344 0 128400 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 129724 0 129780 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 131196 0 131252 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 132668 0 132724 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 134140 0 134196 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 135612 0 135668 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 137084 0 137140 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 138556 0 138612 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 59252 0 59308 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 140028 0 140084 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 141500 0 141556 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 142972 0 143028 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 144444 0 144500 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 145916 0 145972 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 147388 0 147444 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 148860 0 148916 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 150332 0 150388 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 151804 0 151860 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 153276 0 153332 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 60724 0 60780 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 154748 0 154804 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 156220 0 156276 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 157692 0 157748 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 159164 0 159220 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 160636 0 160692 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 162108 0 162164 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 163580 0 163636 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 165052 0 165108 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 166524 0 166580 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 167996 0 168052 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 62196 0 62252 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 169468 0 169524 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 170940 0 170996 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 172412 0 172468 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 173884 0 173940 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 175356 0 175412 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 176828 0 176884 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 178300 0 178356 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 179772 0 179828 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 181244 0 181300 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 182716 0 182772 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 63668 0 63724 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 184188 0 184244 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 185568 0 185624 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 187040 0 187096 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 188512 0 188568 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 189984 0 190040 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 191456 0 191512 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 192928 0 192984 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 194400 0 194456 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 195872 0 195928 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 197344 0 197400 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 65140 0 65196 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 52352 0 52408 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 199368 0 199424 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 200840 0 200896 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 202312 0 202368 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 203692 0 203748 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 205164 0 205220 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 206636 0 206692 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 208108 0 208164 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 209580 0 209636 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 211052 0 211108 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 212524 0 212580 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 67072 0 67128 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 213996 0 214052 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 215468 0 215524 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 216940 0 216996 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 218412 0 218468 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 219884 0 219940 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 221356 0 221412 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 222828 0 222884 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 224300 0 224356 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 225772 0 225828 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 227244 0 227300 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 68544 0 68600 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 228716 0 228772 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 230188 0 230244 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 231660 0 231716 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 233132 0 233188 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 234604 0 234660 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 236076 0 236132 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 237548 0 237604 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 239020 0 239076 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 70016 0 70072 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 71488 0 71544 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 72960 0 73016 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 74432 0 74488 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 75904 0 75960 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 77376 0 77432 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 78848 0 78904 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 80320 0 80376 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 53824 0 53880 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 81792 0 81848 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 83264 0 83320 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 84736 0 84792 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 86208 0 86264 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 87680 0 87736 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 89152 0 89208 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 90624 0 90680 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 92096 0 92152 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 93476 0 93532 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 94948 0 95004 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 55296 0 55352 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 96420 0 96476 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 97892 0 97948 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 99364 0 99420 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 100836 0 100892 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 102308 0 102364 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 103780 0 103836 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 105252 0 105308 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 106724 0 106780 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 108196 0 108252 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 109668 0 109724 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 56768 0 56824 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 111140 0 111196 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 112612 0 112668 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 114084 0 114140 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 115556 0 115612 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 117028 0 117084 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 118500 0 118556 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 119972 0 120028 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 121444 0 121500 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 122916 0 122972 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 124388 0 124444 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 58240 0 58296 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 125860 0 125916 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 127332 0 127388 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 128804 0 128860 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 130276 0 130332 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 131748 0 131804 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 133220 0 133276 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 134692 0 134748 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 136164 0 136220 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 137636 0 137692 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 139108 0 139164 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 59712 0 59768 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 140580 0 140636 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 142052 0 142108 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 143524 0 143580 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 144996 0 145052 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 146468 0 146524 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 147848 0 147904 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 149320 0 149376 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 150792 0 150848 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 152264 0 152320 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 153736 0 153792 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 61184 0 61240 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 155208 0 155264 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 156680 0 156736 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 158152 0 158208 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 159624 0 159680 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 161096 0 161152 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 162568 0 162624 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 164040 0 164096 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 165512 0 165568 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 166984 0 167040 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 168456 0 168512 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 62656 0 62712 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 169928 0 169984 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 171400 0 171456 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 172872 0 172928 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 174344 0 174400 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 175816 0 175872 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 177288 0 177344 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 178760 0 178816 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 180232 0 180288 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 181704 0 181760 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 183176 0 183232 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 64128 0 64184 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 184648 0 184704 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 186120 0 186176 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 187592 0 187648 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 189064 0 189120 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 190536 0 190592 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 192008 0 192064 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 193480 0 193536 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 194952 0 195008 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 196424 0 196480 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 197896 0 197952 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 65600 0 65656 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 52904 0 52960 800 6 la_oen[0]
port 371 nsew signal input
rlabel metal2 s 199828 0 199884 800 6 la_oen[100]
port 372 nsew signal input
rlabel metal2 s 201300 0 201356 800 6 la_oen[101]
port 373 nsew signal input
rlabel metal2 s 202772 0 202828 800 6 la_oen[102]
port 374 nsew signal input
rlabel metal2 s 204244 0 204300 800 6 la_oen[103]
port 375 nsew signal input
rlabel metal2 s 205716 0 205772 800 6 la_oen[104]
port 376 nsew signal input
rlabel metal2 s 207188 0 207244 800 6 la_oen[105]
port 377 nsew signal input
rlabel metal2 s 208660 0 208716 800 6 la_oen[106]
port 378 nsew signal input
rlabel metal2 s 210132 0 210188 800 6 la_oen[107]
port 379 nsew signal input
rlabel metal2 s 211604 0 211660 800 6 la_oen[108]
port 380 nsew signal input
rlabel metal2 s 213076 0 213132 800 6 la_oen[109]
port 381 nsew signal input
rlabel metal2 s 67532 0 67588 800 6 la_oen[10]
port 382 nsew signal input
rlabel metal2 s 214548 0 214604 800 6 la_oen[110]
port 383 nsew signal input
rlabel metal2 s 216020 0 216076 800 6 la_oen[111]
port 384 nsew signal input
rlabel metal2 s 217492 0 217548 800 6 la_oen[112]
port 385 nsew signal input
rlabel metal2 s 218964 0 219020 800 6 la_oen[113]
port 386 nsew signal input
rlabel metal2 s 220436 0 220492 800 6 la_oen[114]
port 387 nsew signal input
rlabel metal2 s 221816 0 221872 800 6 la_oen[115]
port 388 nsew signal input
rlabel metal2 s 223288 0 223344 800 6 la_oen[116]
port 389 nsew signal input
rlabel metal2 s 224760 0 224816 800 6 la_oen[117]
port 390 nsew signal input
rlabel metal2 s 226232 0 226288 800 6 la_oen[118]
port 391 nsew signal input
rlabel metal2 s 227704 0 227760 800 6 la_oen[119]
port 392 nsew signal input
rlabel metal2 s 69004 0 69060 800 6 la_oen[11]
port 393 nsew signal input
rlabel metal2 s 229176 0 229232 800 6 la_oen[120]
port 394 nsew signal input
rlabel metal2 s 230648 0 230704 800 6 la_oen[121]
port 395 nsew signal input
rlabel metal2 s 232120 0 232176 800 6 la_oen[122]
port 396 nsew signal input
rlabel metal2 s 233592 0 233648 800 6 la_oen[123]
port 397 nsew signal input
rlabel metal2 s 235064 0 235120 800 6 la_oen[124]
port 398 nsew signal input
rlabel metal2 s 236536 0 236592 800 6 la_oen[125]
port 399 nsew signal input
rlabel metal2 s 238008 0 238064 800 6 la_oen[126]
port 400 nsew signal input
rlabel metal2 s 239480 0 239536 800 6 la_oen[127]
port 401 nsew signal input
rlabel metal2 s 70476 0 70532 800 6 la_oen[12]
port 402 nsew signal input
rlabel metal2 s 71948 0 72004 800 6 la_oen[13]
port 403 nsew signal input
rlabel metal2 s 73420 0 73476 800 6 la_oen[14]
port 404 nsew signal input
rlabel metal2 s 74892 0 74948 800 6 la_oen[15]
port 405 nsew signal input
rlabel metal2 s 76364 0 76420 800 6 la_oen[16]
port 406 nsew signal input
rlabel metal2 s 77836 0 77892 800 6 la_oen[17]
port 407 nsew signal input
rlabel metal2 s 79308 0 79364 800 6 la_oen[18]
port 408 nsew signal input
rlabel metal2 s 80780 0 80836 800 6 la_oen[19]
port 409 nsew signal input
rlabel metal2 s 54376 0 54432 800 6 la_oen[1]
port 410 nsew signal input
rlabel metal2 s 82252 0 82308 800 6 la_oen[20]
port 411 nsew signal input
rlabel metal2 s 83724 0 83780 800 6 la_oen[21]
port 412 nsew signal input
rlabel metal2 s 85196 0 85252 800 6 la_oen[22]
port 413 nsew signal input
rlabel metal2 s 86668 0 86724 800 6 la_oen[23]
port 414 nsew signal input
rlabel metal2 s 88140 0 88196 800 6 la_oen[24]
port 415 nsew signal input
rlabel metal2 s 89612 0 89668 800 6 la_oen[25]
port 416 nsew signal input
rlabel metal2 s 91084 0 91140 800 6 la_oen[26]
port 417 nsew signal input
rlabel metal2 s 92556 0 92612 800 6 la_oen[27]
port 418 nsew signal input
rlabel metal2 s 94028 0 94084 800 6 la_oen[28]
port 419 nsew signal input
rlabel metal2 s 95500 0 95556 800 6 la_oen[29]
port 420 nsew signal input
rlabel metal2 s 55756 0 55812 800 6 la_oen[2]
port 421 nsew signal input
rlabel metal2 s 96972 0 97028 800 6 la_oen[30]
port 422 nsew signal input
rlabel metal2 s 98444 0 98500 800 6 la_oen[31]
port 423 nsew signal input
rlabel metal2 s 99916 0 99972 800 6 la_oen[32]
port 424 nsew signal input
rlabel metal2 s 101388 0 101444 800 6 la_oen[33]
port 425 nsew signal input
rlabel metal2 s 102860 0 102916 800 6 la_oen[34]
port 426 nsew signal input
rlabel metal2 s 104332 0 104388 800 6 la_oen[35]
port 427 nsew signal input
rlabel metal2 s 105804 0 105860 800 6 la_oen[36]
port 428 nsew signal input
rlabel metal2 s 107276 0 107332 800 6 la_oen[37]
port 429 nsew signal input
rlabel metal2 s 108748 0 108804 800 6 la_oen[38]
port 430 nsew signal input
rlabel metal2 s 110220 0 110276 800 6 la_oen[39]
port 431 nsew signal input
rlabel metal2 s 57228 0 57284 800 6 la_oen[3]
port 432 nsew signal input
rlabel metal2 s 111600 0 111656 800 6 la_oen[40]
port 433 nsew signal input
rlabel metal2 s 113072 0 113128 800 6 la_oen[41]
port 434 nsew signal input
rlabel metal2 s 114544 0 114600 800 6 la_oen[42]
port 435 nsew signal input
rlabel metal2 s 116016 0 116072 800 6 la_oen[43]
port 436 nsew signal input
rlabel metal2 s 117488 0 117544 800 6 la_oen[44]
port 437 nsew signal input
rlabel metal2 s 118960 0 119016 800 6 la_oen[45]
port 438 nsew signal input
rlabel metal2 s 120432 0 120488 800 6 la_oen[46]
port 439 nsew signal input
rlabel metal2 s 121904 0 121960 800 6 la_oen[47]
port 440 nsew signal input
rlabel metal2 s 123376 0 123432 800 6 la_oen[48]
port 441 nsew signal input
rlabel metal2 s 124848 0 124904 800 6 la_oen[49]
port 442 nsew signal input
rlabel metal2 s 58700 0 58756 800 6 la_oen[4]
port 443 nsew signal input
rlabel metal2 s 126320 0 126376 800 6 la_oen[50]
port 444 nsew signal input
rlabel metal2 s 127792 0 127848 800 6 la_oen[51]
port 445 nsew signal input
rlabel metal2 s 129264 0 129320 800 6 la_oen[52]
port 446 nsew signal input
rlabel metal2 s 130736 0 130792 800 6 la_oen[53]
port 447 nsew signal input
rlabel metal2 s 132208 0 132264 800 6 la_oen[54]
port 448 nsew signal input
rlabel metal2 s 133680 0 133736 800 6 la_oen[55]
port 449 nsew signal input
rlabel metal2 s 135152 0 135208 800 6 la_oen[56]
port 450 nsew signal input
rlabel metal2 s 136624 0 136680 800 6 la_oen[57]
port 451 nsew signal input
rlabel metal2 s 138096 0 138152 800 6 la_oen[58]
port 452 nsew signal input
rlabel metal2 s 139568 0 139624 800 6 la_oen[59]
port 453 nsew signal input
rlabel metal2 s 60172 0 60228 800 6 la_oen[5]
port 454 nsew signal input
rlabel metal2 s 141040 0 141096 800 6 la_oen[60]
port 455 nsew signal input
rlabel metal2 s 142512 0 142568 800 6 la_oen[61]
port 456 nsew signal input
rlabel metal2 s 143984 0 144040 800 6 la_oen[62]
port 457 nsew signal input
rlabel metal2 s 145456 0 145512 800 6 la_oen[63]
port 458 nsew signal input
rlabel metal2 s 146928 0 146984 800 6 la_oen[64]
port 459 nsew signal input
rlabel metal2 s 148400 0 148456 800 6 la_oen[65]
port 460 nsew signal input
rlabel metal2 s 149872 0 149928 800 6 la_oen[66]
port 461 nsew signal input
rlabel metal2 s 151344 0 151400 800 6 la_oen[67]
port 462 nsew signal input
rlabel metal2 s 152816 0 152872 800 6 la_oen[68]
port 463 nsew signal input
rlabel metal2 s 154288 0 154344 800 6 la_oen[69]
port 464 nsew signal input
rlabel metal2 s 61644 0 61700 800 6 la_oen[6]
port 465 nsew signal input
rlabel metal2 s 155760 0 155816 800 6 la_oen[70]
port 466 nsew signal input
rlabel metal2 s 157232 0 157288 800 6 la_oen[71]
port 467 nsew signal input
rlabel metal2 s 158704 0 158760 800 6 la_oen[72]
port 468 nsew signal input
rlabel metal2 s 160176 0 160232 800 6 la_oen[73]
port 469 nsew signal input
rlabel metal2 s 161648 0 161704 800 6 la_oen[74]
port 470 nsew signal input
rlabel metal2 s 163120 0 163176 800 6 la_oen[75]
port 471 nsew signal input
rlabel metal2 s 164592 0 164648 800 6 la_oen[76]
port 472 nsew signal input
rlabel metal2 s 166064 0 166120 800 6 la_oen[77]
port 473 nsew signal input
rlabel metal2 s 167444 0 167500 800 6 la_oen[78]
port 474 nsew signal input
rlabel metal2 s 168916 0 168972 800 6 la_oen[79]
port 475 nsew signal input
rlabel metal2 s 63116 0 63172 800 6 la_oen[7]
port 476 nsew signal input
rlabel metal2 s 170388 0 170444 800 6 la_oen[80]
port 477 nsew signal input
rlabel metal2 s 171860 0 171916 800 6 la_oen[81]
port 478 nsew signal input
rlabel metal2 s 173332 0 173388 800 6 la_oen[82]
port 479 nsew signal input
rlabel metal2 s 174804 0 174860 800 6 la_oen[83]
port 480 nsew signal input
rlabel metal2 s 176276 0 176332 800 6 la_oen[84]
port 481 nsew signal input
rlabel metal2 s 177748 0 177804 800 6 la_oen[85]
port 482 nsew signal input
rlabel metal2 s 179220 0 179276 800 6 la_oen[86]
port 483 nsew signal input
rlabel metal2 s 180692 0 180748 800 6 la_oen[87]
port 484 nsew signal input
rlabel metal2 s 182164 0 182220 800 6 la_oen[88]
port 485 nsew signal input
rlabel metal2 s 183636 0 183692 800 6 la_oen[89]
port 486 nsew signal input
rlabel metal2 s 64588 0 64644 800 6 la_oen[8]
port 487 nsew signal input
rlabel metal2 s 185108 0 185164 800 6 la_oen[90]
port 488 nsew signal input
rlabel metal2 s 186580 0 186636 800 6 la_oen[91]
port 489 nsew signal input
rlabel metal2 s 188052 0 188108 800 6 la_oen[92]
port 490 nsew signal input
rlabel metal2 s 189524 0 189580 800 6 la_oen[93]
port 491 nsew signal input
rlabel metal2 s 190996 0 191052 800 6 la_oen[94]
port 492 nsew signal input
rlabel metal2 s 192468 0 192524 800 6 la_oen[95]
port 493 nsew signal input
rlabel metal2 s 193940 0 193996 800 6 la_oen[96]
port 494 nsew signal input
rlabel metal2 s 195412 0 195468 800 6 la_oen[97]
port 495 nsew signal input
rlabel metal2 s 196884 0 196940 800 6 la_oen[98]
port 496 nsew signal input
rlabel metal2 s 198356 0 198412 800 6 la_oen[99]
port 497 nsew signal input
rlabel metal2 s 66060 0 66116 800 6 la_oen[9]
port 498 nsew signal input
rlabel metal2 s 4 0 60 800 6 wb_clk_i
port 499 nsew signal input
rlabel metal2 s 464 0 520 800 6 wb_rst_i
port 500 nsew signal input
rlabel metal2 s 924 0 980 800 6 wbs_ack_o
port 501 nsew signal output
rlabel metal2 s 2856 0 2912 800 6 wbs_adr_i[0]
port 502 nsew signal input
rlabel metal2 s 19508 0 19564 800 6 wbs_adr_i[10]
port 503 nsew signal input
rlabel metal2 s 20980 0 21036 800 6 wbs_adr_i[11]
port 504 nsew signal input
rlabel metal2 s 22452 0 22508 800 6 wbs_adr_i[12]
port 505 nsew signal input
rlabel metal2 s 23924 0 23980 800 6 wbs_adr_i[13]
port 506 nsew signal input
rlabel metal2 s 25396 0 25452 800 6 wbs_adr_i[14]
port 507 nsew signal input
rlabel metal2 s 26868 0 26924 800 6 wbs_adr_i[15]
port 508 nsew signal input
rlabel metal2 s 28340 0 28396 800 6 wbs_adr_i[16]
port 509 nsew signal input
rlabel metal2 s 29812 0 29868 800 6 wbs_adr_i[17]
port 510 nsew signal input
rlabel metal2 s 31284 0 31340 800 6 wbs_adr_i[18]
port 511 nsew signal input
rlabel metal2 s 32756 0 32812 800 6 wbs_adr_i[19]
port 512 nsew signal input
rlabel metal2 s 4880 0 4936 800 6 wbs_adr_i[1]
port 513 nsew signal input
rlabel metal2 s 34228 0 34284 800 6 wbs_adr_i[20]
port 514 nsew signal input
rlabel metal2 s 35700 0 35756 800 6 wbs_adr_i[21]
port 515 nsew signal input
rlabel metal2 s 37172 0 37228 800 6 wbs_adr_i[22]
port 516 nsew signal input
rlabel metal2 s 38644 0 38700 800 6 wbs_adr_i[23]
port 517 nsew signal input
rlabel metal2 s 40116 0 40172 800 6 wbs_adr_i[24]
port 518 nsew signal input
rlabel metal2 s 41588 0 41644 800 6 wbs_adr_i[25]
port 519 nsew signal input
rlabel metal2 s 43060 0 43116 800 6 wbs_adr_i[26]
port 520 nsew signal input
rlabel metal2 s 44532 0 44588 800 6 wbs_adr_i[27]
port 521 nsew signal input
rlabel metal2 s 46004 0 46060 800 6 wbs_adr_i[28]
port 522 nsew signal input
rlabel metal2 s 47476 0 47532 800 6 wbs_adr_i[29]
port 523 nsew signal input
rlabel metal2 s 6812 0 6868 800 6 wbs_adr_i[2]
port 524 nsew signal input
rlabel metal2 s 48948 0 49004 800 6 wbs_adr_i[30]
port 525 nsew signal input
rlabel metal2 s 50420 0 50476 800 6 wbs_adr_i[31]
port 526 nsew signal input
rlabel metal2 s 8744 0 8800 800 6 wbs_adr_i[3]
port 527 nsew signal input
rlabel metal2 s 10768 0 10824 800 6 wbs_adr_i[4]
port 528 nsew signal input
rlabel metal2 s 12240 0 12296 800 6 wbs_adr_i[5]
port 529 nsew signal input
rlabel metal2 s 13712 0 13768 800 6 wbs_adr_i[6]
port 530 nsew signal input
rlabel metal2 s 15184 0 15240 800 6 wbs_adr_i[7]
port 531 nsew signal input
rlabel metal2 s 16656 0 16712 800 6 wbs_adr_i[8]
port 532 nsew signal input
rlabel metal2 s 18128 0 18184 800 6 wbs_adr_i[9]
port 533 nsew signal input
rlabel metal2 s 1384 0 1440 800 6 wbs_cyc_i
port 534 nsew signal input
rlabel metal2 s 3408 0 3464 800 6 wbs_dat_i[0]
port 535 nsew signal input
rlabel metal2 s 20060 0 20116 800 6 wbs_dat_i[10]
port 536 nsew signal input
rlabel metal2 s 21532 0 21588 800 6 wbs_dat_i[11]
port 537 nsew signal input
rlabel metal2 s 23004 0 23060 800 6 wbs_dat_i[12]
port 538 nsew signal input
rlabel metal2 s 24476 0 24532 800 6 wbs_dat_i[13]
port 539 nsew signal input
rlabel metal2 s 25948 0 26004 800 6 wbs_dat_i[14]
port 540 nsew signal input
rlabel metal2 s 27420 0 27476 800 6 wbs_dat_i[15]
port 541 nsew signal input
rlabel metal2 s 28892 0 28948 800 6 wbs_dat_i[16]
port 542 nsew signal input
rlabel metal2 s 30364 0 30420 800 6 wbs_dat_i[17]
port 543 nsew signal input
rlabel metal2 s 31836 0 31892 800 6 wbs_dat_i[18]
port 544 nsew signal input
rlabel metal2 s 33308 0 33364 800 6 wbs_dat_i[19]
port 545 nsew signal input
rlabel metal2 s 5340 0 5396 800 6 wbs_dat_i[1]
port 546 nsew signal input
rlabel metal2 s 34780 0 34836 800 6 wbs_dat_i[20]
port 547 nsew signal input
rlabel metal2 s 36252 0 36308 800 6 wbs_dat_i[21]
port 548 nsew signal input
rlabel metal2 s 37632 0 37688 800 6 wbs_dat_i[22]
port 549 nsew signal input
rlabel metal2 s 39104 0 39160 800 6 wbs_dat_i[23]
port 550 nsew signal input
rlabel metal2 s 40576 0 40632 800 6 wbs_dat_i[24]
port 551 nsew signal input
rlabel metal2 s 42048 0 42104 800 6 wbs_dat_i[25]
port 552 nsew signal input
rlabel metal2 s 43520 0 43576 800 6 wbs_dat_i[26]
port 553 nsew signal input
rlabel metal2 s 44992 0 45048 800 6 wbs_dat_i[27]
port 554 nsew signal input
rlabel metal2 s 46464 0 46520 800 6 wbs_dat_i[28]
port 555 nsew signal input
rlabel metal2 s 47936 0 47992 800 6 wbs_dat_i[29]
port 556 nsew signal input
rlabel metal2 s 7272 0 7328 800 6 wbs_dat_i[2]
port 557 nsew signal input
rlabel metal2 s 49408 0 49464 800 6 wbs_dat_i[30]
port 558 nsew signal input
rlabel metal2 s 50880 0 50936 800 6 wbs_dat_i[31]
port 559 nsew signal input
rlabel metal2 s 9296 0 9352 800 6 wbs_dat_i[3]
port 560 nsew signal input
rlabel metal2 s 11228 0 11284 800 6 wbs_dat_i[4]
port 561 nsew signal input
rlabel metal2 s 12700 0 12756 800 6 wbs_dat_i[5]
port 562 nsew signal input
rlabel metal2 s 14172 0 14228 800 6 wbs_dat_i[6]
port 563 nsew signal input
rlabel metal2 s 15644 0 15700 800 6 wbs_dat_i[7]
port 564 nsew signal input
rlabel metal2 s 17116 0 17172 800 6 wbs_dat_i[8]
port 565 nsew signal input
rlabel metal2 s 18588 0 18644 800 6 wbs_dat_i[9]
port 566 nsew signal input
rlabel metal2 s 3868 0 3924 800 6 wbs_dat_o[0]
port 567 nsew signal output
rlabel metal2 s 20520 0 20576 800 6 wbs_dat_o[10]
port 568 nsew signal output
rlabel metal2 s 21992 0 22048 800 6 wbs_dat_o[11]
port 569 nsew signal output
rlabel metal2 s 23464 0 23520 800 6 wbs_dat_o[12]
port 570 nsew signal output
rlabel metal2 s 24936 0 24992 800 6 wbs_dat_o[13]
port 571 nsew signal output
rlabel metal2 s 26408 0 26464 800 6 wbs_dat_o[14]
port 572 nsew signal output
rlabel metal2 s 27880 0 27936 800 6 wbs_dat_o[15]
port 573 nsew signal output
rlabel metal2 s 29352 0 29408 800 6 wbs_dat_o[16]
port 574 nsew signal output
rlabel metal2 s 30824 0 30880 800 6 wbs_dat_o[17]
port 575 nsew signal output
rlabel metal2 s 32296 0 32352 800 6 wbs_dat_o[18]
port 576 nsew signal output
rlabel metal2 s 33768 0 33824 800 6 wbs_dat_o[19]
port 577 nsew signal output
rlabel metal2 s 5800 0 5856 800 6 wbs_dat_o[1]
port 578 nsew signal output
rlabel metal2 s 35240 0 35296 800 6 wbs_dat_o[20]
port 579 nsew signal output
rlabel metal2 s 36712 0 36768 800 6 wbs_dat_o[21]
port 580 nsew signal output
rlabel metal2 s 38184 0 38240 800 6 wbs_dat_o[22]
port 581 nsew signal output
rlabel metal2 s 39656 0 39712 800 6 wbs_dat_o[23]
port 582 nsew signal output
rlabel metal2 s 41128 0 41184 800 6 wbs_dat_o[24]
port 583 nsew signal output
rlabel metal2 s 42600 0 42656 800 6 wbs_dat_o[25]
port 584 nsew signal output
rlabel metal2 s 44072 0 44128 800 6 wbs_dat_o[26]
port 585 nsew signal output
rlabel metal2 s 45544 0 45600 800 6 wbs_dat_o[27]
port 586 nsew signal output
rlabel metal2 s 47016 0 47072 800 6 wbs_dat_o[28]
port 587 nsew signal output
rlabel metal2 s 48488 0 48544 800 6 wbs_dat_o[29]
port 588 nsew signal output
rlabel metal2 s 7824 0 7880 800 6 wbs_dat_o[2]
port 589 nsew signal output
rlabel metal2 s 49960 0 50016 800 6 wbs_dat_o[30]
port 590 nsew signal output
rlabel metal2 s 51432 0 51488 800 6 wbs_dat_o[31]
port 591 nsew signal output
rlabel metal2 s 9756 0 9812 800 6 wbs_dat_o[3]
port 592 nsew signal output
rlabel metal2 s 11688 0 11744 800 6 wbs_dat_o[4]
port 593 nsew signal output
rlabel metal2 s 13160 0 13216 800 6 wbs_dat_o[5]
port 594 nsew signal output
rlabel metal2 s 14632 0 14688 800 6 wbs_dat_o[6]
port 595 nsew signal output
rlabel metal2 s 16104 0 16160 800 6 wbs_dat_o[7]
port 596 nsew signal output
rlabel metal2 s 17576 0 17632 800 6 wbs_dat_o[8]
port 597 nsew signal output
rlabel metal2 s 19048 0 19104 800 6 wbs_dat_o[9]
port 598 nsew signal output
rlabel metal2 s 4328 0 4384 800 6 wbs_sel_i[0]
port 599 nsew signal input
rlabel metal2 s 6352 0 6408 800 6 wbs_sel_i[1]
port 600 nsew signal input
rlabel metal2 s 8284 0 8340 800 6 wbs_sel_i[2]
port 601 nsew signal input
rlabel metal2 s 10216 0 10272 800 6 wbs_sel_i[3]
port 602 nsew signal input
rlabel metal2 s 1936 0 1992 800 6 wbs_stb_i
port 603 nsew signal input
rlabel metal2 s 2396 0 2452 800 6 wbs_we_i
port 604 nsew signal input
rlabel metal4 s 219050 2128 219370 237776 6 VPWR
port 605 nsew power bidirectional
rlabel metal4 s 188330 2128 188650 237776 6 VPWR
port 606 nsew power bidirectional
rlabel metal4 s 157610 2128 157930 237776 6 VPWR
port 607 nsew power bidirectional
rlabel metal4 s 126890 2128 127210 237776 6 VPWR
port 608 nsew power bidirectional
rlabel metal4 s 96170 2128 96490 237776 6 VPWR
port 609 nsew power bidirectional
rlabel metal4 s 65450 2128 65770 237776 6 VPWR
port 610 nsew power bidirectional
rlabel metal4 s 34730 2128 35050 237776 6 VPWR
port 611 nsew power bidirectional
rlabel metal4 s 4010 2128 4330 237776 6 VPWR
port 612 nsew power bidirectional
rlabel metal4 s 234410 2128 234730 237776 6 VGND
port 613 nsew ground bidirectional
rlabel metal4 s 203690 2128 204010 237776 6 VGND
port 614 nsew ground bidirectional
rlabel metal4 s 172970 2128 173290 237776 6 VGND
port 615 nsew ground bidirectional
rlabel metal4 s 142250 2128 142570 237776 6 VGND
port 616 nsew ground bidirectional
rlabel metal4 s 111530 2128 111850 237776 6 VGND
port 617 nsew ground bidirectional
rlabel metal4 s 80810 2128 81130 237776 6 VGND
port 618 nsew ground bidirectional
rlabel metal4 s 50090 2128 50410 237776 6 VGND
port 619 nsew ground bidirectional
rlabel metal4 s 19370 2128 19690 237776 6 VGND
port 620 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 239540 240000
string LEFview TRUE
<< end >>
