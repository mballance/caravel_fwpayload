magic
tech sky130A
magscale 1 2
timestamp 1607635834
<< locali >>
rect 429577 666587 429611 684437
rect 494069 666587 494103 676141
rect 559297 666587 559331 684437
rect 429485 647275 429519 656829
rect 559205 647275 559239 656829
rect 428105 639251 428139 639897
rect 436109 639183 436143 639897
rect 443837 639115 443871 639897
rect 451749 639047 451783 639897
rect 520289 638979 520323 639897
rect 234663 337705 235031 337739
rect 234997 337535 235031 337705
rect 236837 337603 236871 337705
rect 239413 337535 239447 337637
rect 228097 337399 228131 337501
rect 267473 337399 267507 337501
rect 228097 337365 228281 337399
rect 267565 328491 267599 337501
rect 326353 337195 326387 337909
rect 384313 337603 384347 337909
rect 389005 337535 389039 337841
rect 347789 336991 347823 337161
rect 357357 336991 357391 337297
rect 367109 336719 367143 337297
rect 377045 336787 377079 337501
rect 386429 337331 386463 337501
rect 379437 336787 379471 337297
rect 395353 336923 395387 337977
rect 398757 337331 398791 337909
rect 398849 337195 398883 337841
rect 404001 337331 404035 337841
rect 421021 336855 421055 337161
rect 422953 336923 422987 337909
rect 432521 337603 432555 337909
rect 432613 337807 432647 337909
rect 432705 337467 432739 337773
rect 499037 337603 499071 337977
rect 529063 337637 529431 337671
rect 423045 337263 423079 337433
rect 432521 337433 432739 337467
rect 432521 337399 432555 337433
rect 430497 337059 430531 337161
rect 431141 336991 431175 337365
rect 432613 337127 432647 337365
rect 433349 337195 433383 337297
rect 432521 336957 432797 336991
rect 432521 336787 432555 336957
rect 432613 336787 432647 336889
rect 433441 336855 433475 337297
rect 435833 337059 435867 337501
rect 441353 336991 441387 337569
rect 502349 337331 502383 337569
rect 526821 337535 526855 337637
rect 520197 336991 520231 337365
rect 524429 336787 524463 337365
rect 529305 337263 529339 337501
rect 529397 337263 529431 337637
rect 531421 337263 531455 337365
rect 531513 336787 531547 337229
rect 232329 314687 232363 324241
rect 249993 317475 250027 321657
rect 259653 318835 259687 321589
rect 232329 294899 232363 313225
rect 232421 282931 232455 292485
rect 236469 284359 236503 292485
rect 241805 289867 241839 299421
rect 243001 298231 243035 307717
rect 243001 280211 243035 298061
rect 249993 289867 250027 299421
rect 255513 298163 255547 315945
rect 267105 307819 267139 309145
rect 270693 299523 270727 309077
rect 277593 309043 277627 311933
rect 281641 307819 281675 317373
rect 283021 307819 283055 317373
rect 288633 309179 288667 318733
rect 292773 317475 292807 327029
rect 294061 325703 294095 335257
rect 356529 317475 356563 335257
rect 377045 327131 377079 335597
rect 381185 328491 381219 331109
rect 357541 317475 357575 327029
rect 382473 317543 382507 327029
rect 392317 318835 392351 328389
rect 393237 318835 393271 328389
rect 397837 318835 397871 328389
rect 400321 318835 400355 327029
rect 416881 318835 416915 328389
rect 422401 318835 422435 328389
rect 427921 318835 427955 328389
rect 433717 318835 433751 328389
rect 466561 318835 466595 321589
rect 472081 318835 472115 328389
rect 346593 309179 346627 311797
rect 371341 309111 371375 317373
rect 277593 298231 277627 307717
rect 252753 280211 252787 289765
rect 232145 262259 232179 271813
rect 236193 263687 236227 273105
rect 241805 270555 241839 280109
rect 254133 277423 254167 289765
rect 259653 277423 259687 289765
rect 265173 288439 265207 298061
rect 267013 280211 267047 298061
rect 277593 280211 277627 298061
rect 281641 289867 281675 299421
rect 283113 289867 283147 299421
rect 287253 298163 287287 307717
rect 288633 289867 288667 299421
rect 295533 298231 295567 307717
rect 309333 299523 309367 309077
rect 318993 299523 319027 309077
rect 342453 299591 342487 309009
rect 376953 307819 376987 317373
rect 382473 307819 382507 317373
rect 386705 309179 386739 318733
rect 292681 288439 292715 298061
rect 295625 293267 295659 298061
rect 298385 287079 298419 296633
rect 305193 289867 305227 299421
rect 310713 289867 310747 299421
rect 334265 296735 334299 298129
rect 346593 289867 346627 299421
rect 364533 298163 364567 307717
rect 400505 299455 400539 315945
rect 408785 302107 408819 315945
rect 416881 299523 416915 309077
rect 422493 299931 422527 309077
rect 428013 299523 428047 309077
rect 433441 299523 433475 309077
rect 451565 302107 451599 315945
rect 466561 299523 466595 309077
rect 472081 299523 472115 309077
rect 480361 307819 480395 317373
rect 309333 280211 309367 289697
rect 334265 282795 334299 289765
rect 347973 288439 348007 298061
rect 352113 287963 352147 298061
rect 364533 284971 364567 291329
rect 370053 288439 370087 298061
rect 375481 289799 375515 298061
rect 376953 289867 376987 299421
rect 397745 288439 397779 298061
rect 480361 288439 480395 298061
rect 342545 280279 342579 282897
rect 243093 260899 243127 270453
rect 252753 260899 252787 270453
rect 267105 260899 267139 270453
rect 270601 260899 270635 278681
rect 288633 270555 288667 280109
rect 236285 244375 236319 253861
rect 241805 251243 241839 260797
rect 254133 248523 254167 253997
rect 259653 248523 259687 253997
rect 265265 251243 265299 260797
rect 272073 251243 272107 260797
rect 281825 259471 281859 269025
rect 288633 251243 288667 260797
rect 292681 260763 292715 269025
rect 295441 263483 295475 273921
rect 305193 270555 305227 280109
rect 310713 270555 310747 280109
rect 321753 272187 321787 280109
rect 327273 272187 327307 280109
rect 334357 273207 334391 280109
rect 346593 270555 346627 280109
rect 356437 270487 356471 273309
rect 381093 270555 381127 280041
rect 382473 270555 382507 280109
rect 386613 278783 386647 287045
rect 408693 278783 408727 288337
rect 309333 260899 309367 270385
rect 324421 260899 324455 263585
rect 342545 260899 342579 263585
rect 381093 260899 381127 270385
rect 386613 269195 386647 273241
rect 397653 269127 397687 278545
rect 416881 270555 416915 280109
rect 433625 270555 433659 280109
rect 294153 251243 294187 260797
rect 295533 251243 295567 260797
rect 305193 251243 305227 260797
rect 309333 251243 309367 260729
rect 310713 251243 310747 260797
rect 321753 251243 321787 260797
rect 327273 251243 327307 260797
rect 334357 251311 334391 260797
rect 342453 251243 342487 260729
rect 346593 251243 346627 260797
rect 254133 244239 254167 248353
rect 236285 234651 236319 244205
rect 292773 240159 292807 251141
rect 324421 241587 324455 244273
rect 334357 244171 334391 251141
rect 348065 241519 348099 250053
rect 353585 241519 353619 251141
rect 370053 248523 370087 253997
rect 375573 248523 375607 253997
rect 382473 251243 382507 260797
rect 386521 259471 386555 264265
rect 392041 259471 392075 264265
rect 400505 260899 400539 270453
rect 451565 263483 451599 273717
rect 466561 270555 466595 280109
rect 472081 270555 472115 280109
rect 397561 249815 397595 253929
rect 416881 251243 416915 260797
rect 433625 251243 433659 260797
rect 375573 242811 375607 248353
rect 397561 240159 397595 244953
rect 400505 241519 400539 251141
rect 451565 244171 451599 259369
rect 466561 251243 466595 260797
rect 472081 251243 472115 260797
rect 236285 215339 236319 224825
rect 259653 222207 259687 231761
rect 292773 230503 292807 239989
rect 243093 212551 243127 222037
rect 270693 212483 270727 215373
rect 281733 212483 281767 229041
rect 309333 222207 309367 231761
rect 331321 227783 331355 231829
rect 451289 222207 451323 224961
rect 334357 212483 334391 219385
rect 243185 202895 243219 205649
rect 259653 202895 259687 212449
rect 265265 202895 265299 205649
rect 270693 205615 270727 211089
rect 295533 202827 295567 209729
rect 364165 208403 364199 212517
rect 364349 212415 364383 212789
rect 408785 212551 408819 215305
rect 336841 202895 336875 205649
rect 369961 202895 369995 212449
rect 243093 193239 243127 202725
rect 480269 201535 480303 202929
rect 255513 190519 255547 200073
rect 270601 193171 270635 196061
rect 281917 193171 281951 201433
rect 236285 178075 236319 187561
rect 270601 183515 270635 191777
rect 271981 183583 272015 186405
rect 295717 183515 295751 200073
rect 298293 183583 298327 186405
rect 309333 183583 309367 201433
rect 332793 189091 332827 198645
rect 352113 193171 352147 201433
rect 359197 187731 359231 197285
rect 369961 193171 369995 201433
rect 375573 193239 375607 196061
rect 321661 183583 321695 186405
rect 324421 183583 324455 186405
rect 252753 173927 252787 178789
rect 243001 162911 243035 167093
rect 254133 166991 254167 172465
rect 255513 166991 255547 180761
rect 267197 173315 267231 182121
rect 336841 176579 336875 182121
rect 259653 162911 259687 172465
rect 265173 154683 265207 164169
rect 271981 162911 272015 172465
rect 292773 164203 292807 172465
rect 342361 162911 342395 172465
rect 347973 162911 348007 180761
rect 352113 162911 352147 180761
rect 353493 162911 353527 180761
rect 357633 179435 357667 186405
rect 364533 186303 364567 190417
rect 386613 186303 386647 198645
rect 433717 193239 433751 196061
rect 397745 173927 397779 176613
rect 236377 143463 236411 151725
rect 243001 147611 243035 154513
rect 254409 143599 254443 153085
rect 271981 148631 272015 157981
rect 298293 157335 298327 162809
rect 292773 147611 292807 155873
rect 331413 147475 331447 154513
rect 334541 153187 334575 161381
rect 356437 151827 356471 161313
rect 370053 154615 370087 164169
rect 376953 154615 376987 164169
rect 382473 154615 382507 167637
rect 243277 124219 243311 133841
rect 254225 124219 254259 143497
rect 259653 133807 259687 143497
rect 283021 132515 283055 142069
rect 287253 133943 287287 143497
rect 292773 135303 292807 144857
rect 305101 133943 305135 143497
rect 321661 135235 321695 143497
rect 334449 142171 334483 151725
rect 375573 147611 375607 154513
rect 381093 147611 381127 154513
rect 392133 147611 392167 154513
rect 393237 145027 393271 162809
rect 397745 154615 397779 164169
rect 400505 157335 400539 164169
rect 422401 157335 422435 164169
rect 451565 147611 451599 162809
rect 466561 157335 466595 164169
rect 480269 153255 480303 164169
rect 381093 135303 381127 144789
rect 397745 143599 397779 144925
rect 393237 133943 393271 143497
rect 400505 137955 400539 144857
rect 422401 137955 422435 144857
rect 466561 137955 466595 144857
rect 240149 114563 240183 124117
rect 249993 114563 250027 124117
rect 267197 122859 267231 132413
rect 292773 125579 292807 133841
rect 304917 124219 304951 125681
rect 236285 103547 236319 113101
rect 240149 96679 240183 106233
rect 243093 106199 243127 109701
rect 252753 106335 252787 119357
rect 271981 115379 272015 124117
rect 287161 114563 287195 124117
rect 292865 113203 292899 124117
rect 236285 85595 236319 95149
rect 240149 85663 240183 95149
rect 254225 93891 254259 103445
rect 266461 92531 266495 102085
rect 281641 101371 281675 106233
rect 282929 95251 282963 104805
rect 295533 103547 295567 113101
rect 298201 111843 298235 118745
rect 310713 118643 310747 125545
rect 334449 124219 334483 133841
rect 353493 124219 353527 133841
rect 356437 124219 356471 133841
rect 298385 102187 298419 111673
rect 305101 106335 305135 115889
rect 321753 114563 321787 118813
rect 324513 114563 324547 118813
rect 327273 113203 327307 122757
rect 330033 106335 330067 120241
rect 342637 114563 342671 124117
rect 365913 118643 365947 124117
rect 381185 115991 381219 125545
rect 386613 122927 386647 133841
rect 348065 113203 348099 114529
rect 288633 96679 288667 99365
rect 236285 75939 236319 85425
rect 241805 77299 241839 86921
rect 287161 85663 287195 95149
rect 298385 93823 298419 99433
rect 308137 96679 308171 99365
rect 243185 67643 243219 80733
rect 249993 79339 250027 85493
rect 244473 67643 244507 70465
rect 254133 67643 254167 85493
rect 255513 74579 255547 79985
rect 259653 71111 259687 84133
rect 266461 64923 266495 77945
rect 270693 66283 270727 75837
rect 271981 73219 272015 82773
rect 281733 75939 281767 77265
rect 287253 75939 287287 85493
rect 288633 77299 288667 86921
rect 294153 84235 294187 93653
rect 309241 89675 309275 104805
rect 310713 96679 310747 99365
rect 319085 95251 319119 104805
rect 324513 96679 324547 106233
rect 353493 93891 353527 103445
rect 357633 96543 357667 106233
rect 386889 103547 386923 121397
rect 407773 114563 407807 124117
rect 433625 115991 433659 125545
rect 466653 114563 466687 124117
rect 397653 104975 397687 114461
rect 408693 104907 408727 114461
rect 393145 98719 393179 104805
rect 400505 95251 400539 104805
rect 298569 84235 298603 88961
rect 305193 77299 305227 86921
rect 308137 77299 308171 86921
rect 309333 77299 309367 80053
rect 310713 77299 310747 86921
rect 334265 79339 334299 85493
rect 342545 80019 342579 86921
rect 346593 80019 346627 86921
rect 364533 84235 364567 93789
rect 375573 85595 375607 93517
rect 381001 87023 381035 89777
rect 407773 87023 407807 104805
rect 408785 89675 408819 100045
rect 422401 99331 422435 106233
rect 427921 99331 427955 106233
rect 433625 99331 433659 106233
rect 480453 95251 480487 104805
rect 305193 67643 305227 70465
rect 249901 56559 249935 64821
rect 240241 46971 240275 56525
rect 255513 55267 255547 64821
rect 281733 61455 281767 67541
rect 283113 56627 283147 66181
rect 287253 56695 287287 66181
rect 249901 47039 249935 51153
rect 231961 37315 231995 46869
rect 236285 37315 236319 46869
rect 244473 37315 244507 46869
rect 249901 37315 249935 46869
rect 267013 45611 267047 55097
rect 271981 46971 272015 51765
rect 281641 46971 281675 56525
rect 287253 47039 287287 56525
rect 292773 47039 292807 66181
rect 310621 55267 310655 64821
rect 324513 56627 324547 66181
rect 334357 64991 334391 74477
rect 352021 66283 352055 77333
rect 356437 73219 356471 82773
rect 357725 74579 357759 84133
rect 359013 77979 359047 84133
rect 381001 75939 381035 85493
rect 382473 75939 382507 86921
rect 407773 75939 407807 85493
rect 408693 76007 408727 85493
rect 422401 77299 422435 86921
rect 433625 77299 433659 80189
rect 466469 77163 466503 85493
rect 364533 64923 364567 74477
rect 375573 66351 375607 75837
rect 321753 47039 321787 51153
rect 329941 46971 329975 55165
rect 331413 48331 331447 64821
rect 334357 48331 334391 64821
rect 231869 26299 231903 35853
rect 240241 26367 240275 31841
rect 252753 31671 252787 40137
rect 267105 29019 267139 42041
rect 272073 29019 272107 42925
rect 282929 35955 282963 45509
rect 292865 35955 292899 45509
rect 309333 37315 309367 46869
rect 342453 45611 342487 55165
rect 356529 45611 356563 63461
rect 359197 53839 359231 63461
rect 375481 56627 375515 66181
rect 381093 57987 381127 67541
rect 408693 66283 408727 75837
rect 427921 67643 427955 76313
rect 472081 67643 472115 85493
rect 480453 77163 480487 85493
rect 407773 56627 407807 66181
rect 375573 51731 375607 56457
rect 359105 45611 359139 48365
rect 382381 48331 382415 51085
rect 324513 29019 324547 40137
rect 236377 16643 236411 26197
rect 244289 16643 244323 19397
rect 252845 19363 252879 28917
rect 266645 19227 266679 27557
rect 270693 18003 270727 27557
rect 281733 19363 281767 28917
rect 252753 11747 252787 12529
rect 288541 10727 288575 19261
rect 305101 13447 305135 19261
rect 293969 11883 294003 12461
rect 308045 10115 308079 19261
rect 318993 18003 319027 27557
rect 324421 18003 324455 27557
rect 330033 26299 330067 44081
rect 353585 37247 353619 45509
rect 356621 35955 356655 40749
rect 357541 35955 357575 41429
rect 392133 35955 392167 48229
rect 397745 46971 397779 56525
rect 416881 48399 416915 57885
rect 433625 48331 433659 57885
rect 466561 48331 466595 57885
rect 472081 48331 472115 57885
rect 400597 45611 400631 47141
rect 400689 37179 400723 45441
rect 407773 37315 407807 46869
rect 342361 19363 342395 32385
rect 472173 31195 472207 38573
rect 346501 18003 346535 27557
rect 356529 26367 356563 31093
rect 347881 19431 347915 26197
rect 330125 9503 330159 17901
rect 334357 11339 334391 17901
rect 357541 9843 357575 26197
rect 364809 17459 364843 26197
rect 392225 16643 392259 26197
rect 393237 18003 393271 27557
rect 346501 8483 346535 9605
rect 369961 8279 369995 9605
rect 315221 5899 315255 6749
rect 371249 6103 371283 9605
rect 376861 6307 376895 9945
rect 322213 5831 322247 6001
rect 382381 5355 382415 13073
rect 397561 9707 397595 19261
rect 407773 9707 407807 27557
rect 427829 19431 427863 28917
rect 472173 19363 472207 22253
rect 427829 9707 427863 19261
rect 480361 18003 480395 27557
rect 282101 4029 282319 4063
rect 282101 3723 282135 4029
rect 282285 3995 282319 4029
rect 282193 3723 282227 3961
rect 238217 3519 238251 3621
rect 276765 3383 276799 3553
rect 292589 3315 292623 3553
rect 372813 3519 372847 3689
rect 302157 3315 302191 3485
rect 335185 3179 335219 3281
rect 82921 2975 82955 3145
rect 371525 2975 371559 3417
rect 372905 3179 372939 3485
rect 374653 3111 374687 3961
rect 392961 3927 392995 4029
rect 98653 2839 98687 2941
rect 121503 2873 121653 2907
rect 393053 595 393087 9605
rect 393881 3383 393915 4029
rect 393973 3859 394007 4097
rect 403541 3859 403575 4097
rect 403633 3723 403667 3961
rect 403725 3383 403759 3689
rect 403667 3349 403759 3383
rect 403817 3315 403851 3417
rect 406301 3383 406335 4233
rect 408359 4029 408451 4063
rect 408417 3655 408451 4029
rect 409245 3995 409279 4097
rect 408543 3621 408635 3655
rect 403541 3281 403851 3315
rect 403541 3111 403575 3281
rect 403909 3247 403943 3281
rect 408601 3247 408635 3621
rect 416237 3451 416271 4029
rect 423689 3655 423723 4097
rect 409613 3417 409889 3451
rect 409613 3383 409647 3417
rect 403759 3213 403943 3247
rect 403633 3111 403667 3213
rect 408509 3111 408543 3213
rect 408509 3077 408785 3111
rect 408877 3077 410717 3111
rect 408877 3043 408911 3077
rect 408509 3009 408911 3043
rect 408509 2907 408543 3009
rect 418169 2907 418203 3553
rect 423781 3519 423815 3621
rect 421113 2975 421147 3213
rect 421941 3179 421975 3349
rect 422953 3043 422987 3281
rect 426725 2907 426759 3621
rect 432705 3315 432739 3961
rect 447609 3247 447643 3349
rect 509801 3315 509835 3825
rect 516977 3247 517011 4029
rect 569141 3383 569175 3485
rect 540161 3043 540195 3281
<< viali >>
rect 429577 684437 429611 684471
rect 559297 684437 559331 684471
rect 429577 666553 429611 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 559297 666553 559331 666587
rect 429485 656829 429519 656863
rect 429485 647241 429519 647275
rect 559205 656829 559239 656863
rect 559205 647241 559239 647275
rect 428105 639897 428139 639931
rect 428105 639217 428139 639251
rect 436109 639897 436143 639931
rect 436109 639149 436143 639183
rect 443837 639897 443871 639931
rect 443837 639081 443871 639115
rect 451749 639897 451783 639931
rect 451749 639013 451783 639047
rect 520289 639897 520323 639931
rect 520289 638945 520323 638979
rect 395353 337977 395387 338011
rect 326353 337909 326387 337943
rect 234629 337705 234663 337739
rect 236837 337705 236871 337739
rect 236837 337569 236871 337603
rect 239413 337637 239447 337671
rect 228097 337501 228131 337535
rect 234997 337501 235031 337535
rect 239413 337501 239447 337535
rect 267473 337501 267507 337535
rect 228281 337365 228315 337399
rect 267473 337365 267507 337399
rect 267565 337501 267599 337535
rect 384313 337909 384347 337943
rect 384313 337569 384347 337603
rect 389005 337841 389039 337875
rect 377045 337501 377079 337535
rect 357357 337297 357391 337331
rect 326353 337161 326387 337195
rect 347789 337161 347823 337195
rect 347789 336957 347823 336991
rect 357357 336957 357391 336991
rect 367109 337297 367143 337331
rect 386429 337501 386463 337535
rect 389005 337501 389039 337535
rect 377045 336753 377079 336787
rect 379437 337297 379471 337331
rect 386429 337297 386463 337331
rect 499037 337977 499071 338011
rect 398757 337909 398791 337943
rect 422953 337909 422987 337943
rect 398757 337297 398791 337331
rect 398849 337841 398883 337875
rect 404001 337841 404035 337875
rect 404001 337297 404035 337331
rect 398849 337161 398883 337195
rect 421021 337161 421055 337195
rect 395353 336889 395387 336923
rect 432521 337909 432555 337943
rect 432613 337909 432647 337943
rect 432613 337773 432647 337807
rect 432705 337773 432739 337807
rect 432521 337569 432555 337603
rect 526821 337637 526855 337671
rect 529029 337637 529063 337671
rect 441353 337569 441387 337603
rect 499037 337569 499071 337603
rect 502349 337569 502383 337603
rect 423045 337433 423079 337467
rect 435833 337501 435867 337535
rect 423045 337229 423079 337263
rect 431141 337365 431175 337399
rect 432521 337365 432555 337399
rect 432613 337365 432647 337399
rect 430497 337161 430531 337195
rect 430497 337025 430531 337059
rect 433349 337297 433383 337331
rect 433349 337161 433383 337195
rect 433441 337297 433475 337331
rect 432613 337093 432647 337127
rect 431141 336957 431175 336991
rect 432797 336957 432831 336991
rect 422953 336889 422987 336923
rect 421021 336821 421055 336855
rect 379437 336753 379471 336787
rect 432521 336753 432555 336787
rect 432613 336889 432647 336923
rect 435833 337025 435867 337059
rect 526821 337501 526855 337535
rect 529305 337501 529339 337535
rect 502349 337297 502383 337331
rect 520197 337365 520231 337399
rect 441353 336957 441387 336991
rect 520197 336957 520231 336991
rect 524429 337365 524463 337399
rect 433441 336821 433475 336855
rect 432613 336753 432647 336787
rect 529305 337229 529339 337263
rect 529397 337229 529431 337263
rect 531421 337365 531455 337399
rect 531421 337229 531455 337263
rect 531513 337229 531547 337263
rect 524429 336753 524463 336787
rect 531513 336753 531547 336787
rect 367109 336685 367143 336719
rect 377045 335597 377079 335631
rect 267565 328457 267599 328491
rect 294061 335257 294095 335291
rect 292773 327029 292807 327063
rect 232329 324241 232363 324275
rect 249993 321657 250027 321691
rect 259653 321589 259687 321623
rect 259653 318801 259687 318835
rect 249993 317441 250027 317475
rect 288633 318733 288667 318767
rect 281641 317373 281675 317407
rect 232329 314653 232363 314687
rect 255513 315945 255547 315979
rect 232329 313225 232363 313259
rect 243001 307717 243035 307751
rect 232329 294865 232363 294899
rect 241805 299421 241839 299455
rect 232421 292485 232455 292519
rect 236469 292485 236503 292519
rect 243001 298197 243035 298231
rect 249993 299421 250027 299455
rect 241805 289833 241839 289867
rect 243001 298061 243035 298095
rect 236469 284325 236503 284359
rect 232421 282897 232455 282931
rect 277593 311933 277627 311967
rect 267105 309145 267139 309179
rect 267105 307785 267139 307819
rect 270693 309077 270727 309111
rect 277593 309009 277627 309043
rect 281641 307785 281675 307819
rect 283021 317373 283055 317407
rect 294061 325669 294095 325703
rect 356529 335257 356563 335291
rect 292773 317441 292807 317475
rect 381185 331109 381219 331143
rect 381185 328457 381219 328491
rect 377045 327097 377079 327131
rect 392317 328389 392351 328423
rect 356529 317441 356563 317475
rect 357541 327029 357575 327063
rect 382473 327029 382507 327063
rect 392317 318801 392351 318835
rect 393237 328389 393271 328423
rect 393237 318801 393271 318835
rect 397837 328389 397871 328423
rect 416881 328389 416915 328423
rect 397837 318801 397871 318835
rect 400321 327029 400355 327063
rect 400321 318801 400355 318835
rect 416881 318801 416915 318835
rect 422401 328389 422435 328423
rect 422401 318801 422435 318835
rect 427921 328389 427955 328423
rect 427921 318801 427955 318835
rect 433717 328389 433751 328423
rect 472081 328389 472115 328423
rect 433717 318801 433751 318835
rect 466561 321589 466595 321623
rect 466561 318801 466595 318835
rect 472081 318801 472115 318835
rect 382473 317509 382507 317543
rect 386705 318733 386739 318767
rect 357541 317441 357575 317475
rect 371341 317373 371375 317407
rect 288633 309145 288667 309179
rect 346593 311797 346627 311831
rect 346593 309145 346627 309179
rect 283021 307785 283055 307819
rect 309333 309077 309367 309111
rect 270693 299489 270727 299523
rect 277593 307717 277627 307751
rect 287253 307717 287287 307751
rect 277593 298197 277627 298231
rect 281641 299421 281675 299455
rect 255513 298129 255547 298163
rect 249993 289833 250027 289867
rect 265173 298061 265207 298095
rect 243001 280177 243035 280211
rect 252753 289765 252787 289799
rect 252753 280177 252787 280211
rect 254133 289765 254167 289799
rect 241805 280109 241839 280143
rect 236193 273105 236227 273139
rect 232145 271813 232179 271847
rect 254133 277389 254167 277423
rect 259653 289765 259687 289799
rect 265173 288405 265207 288439
rect 267013 298061 267047 298095
rect 267013 280177 267047 280211
rect 277593 298061 277627 298095
rect 281641 289833 281675 289867
rect 283113 299421 283147 299455
rect 295533 307717 295567 307751
rect 287253 298129 287287 298163
rect 288633 299421 288667 299455
rect 283113 289833 283147 289867
rect 309333 299489 309367 299523
rect 318993 309077 319027 309111
rect 371341 309077 371375 309111
rect 376953 317373 376987 317407
rect 342453 309009 342487 309043
rect 376953 307785 376987 307819
rect 382473 317373 382507 317407
rect 480361 317373 480395 317407
rect 386705 309145 386739 309179
rect 400505 315945 400539 315979
rect 382473 307785 382507 307819
rect 342453 299557 342487 299591
rect 364533 307717 364567 307751
rect 318993 299489 319027 299523
rect 295533 298197 295567 298231
rect 305193 299421 305227 299455
rect 288633 289833 288667 289867
rect 292681 298061 292715 298095
rect 295625 298061 295659 298095
rect 295625 293233 295659 293267
rect 298385 296633 298419 296667
rect 292681 288405 292715 288439
rect 305193 289833 305227 289867
rect 310713 299421 310747 299455
rect 346593 299421 346627 299455
rect 334265 298129 334299 298163
rect 334265 296701 334299 296735
rect 310713 289833 310747 289867
rect 408785 315945 408819 315979
rect 451565 315945 451599 315979
rect 408785 302073 408819 302107
rect 416881 309077 416915 309111
rect 422493 309077 422527 309111
rect 422493 299897 422527 299931
rect 428013 309077 428047 309111
rect 416881 299489 416915 299523
rect 428013 299489 428047 299523
rect 433441 309077 433475 309111
rect 451565 302073 451599 302107
rect 466561 309077 466595 309111
rect 433441 299489 433475 299523
rect 466561 299489 466595 299523
rect 472081 309077 472115 309111
rect 480361 307785 480395 307819
rect 472081 299489 472115 299523
rect 364533 298129 364567 298163
rect 376953 299421 376987 299455
rect 400505 299421 400539 299455
rect 346593 289833 346627 289867
rect 347973 298061 348007 298095
rect 334265 289765 334299 289799
rect 298385 287045 298419 287079
rect 309333 289697 309367 289731
rect 277593 280177 277627 280211
rect 347973 288405 348007 288439
rect 352113 298061 352147 298095
rect 370053 298061 370087 298095
rect 352113 287929 352147 287963
rect 364533 291329 364567 291363
rect 375481 298061 375515 298095
rect 376953 289833 376987 289867
rect 397745 298061 397779 298095
rect 375481 289765 375515 289799
rect 370053 288405 370087 288439
rect 397745 288405 397779 288439
rect 480361 298061 480395 298095
rect 480361 288405 480395 288439
rect 408693 288337 408727 288371
rect 364533 284937 364567 284971
rect 386613 287045 386647 287079
rect 334265 282761 334299 282795
rect 342545 282897 342579 282931
rect 342545 280245 342579 280279
rect 309333 280177 309367 280211
rect 288633 280109 288667 280143
rect 259653 277389 259687 277423
rect 270601 278681 270635 278715
rect 241805 270521 241839 270555
rect 236193 263653 236227 263687
rect 243093 270453 243127 270487
rect 232145 262225 232179 262259
rect 243093 260865 243127 260899
rect 252753 270453 252787 270487
rect 252753 260865 252787 260899
rect 267105 270453 267139 270487
rect 267105 260865 267139 260899
rect 305193 280109 305227 280143
rect 288633 270521 288667 270555
rect 295441 273921 295475 273955
rect 270601 260865 270635 260899
rect 281825 269025 281859 269059
rect 241805 260797 241839 260831
rect 236285 253861 236319 253895
rect 265265 260797 265299 260831
rect 241805 251209 241839 251243
rect 254133 253997 254167 254031
rect 254133 248489 254167 248523
rect 259653 253997 259687 254031
rect 265265 251209 265299 251243
rect 272073 260797 272107 260831
rect 292681 269025 292715 269059
rect 281825 259437 281859 259471
rect 288633 260797 288667 260831
rect 272073 251209 272107 251243
rect 305193 270521 305227 270555
rect 310713 280109 310747 280143
rect 321753 280109 321787 280143
rect 321753 272153 321787 272187
rect 327273 280109 327307 280143
rect 334357 280109 334391 280143
rect 334357 273173 334391 273207
rect 346593 280109 346627 280143
rect 327273 272153 327307 272187
rect 310713 270521 310747 270555
rect 382473 280109 382507 280143
rect 381093 280041 381127 280075
rect 346593 270521 346627 270555
rect 356437 273309 356471 273343
rect 381093 270521 381127 270555
rect 386613 278749 386647 278783
rect 408693 278749 408727 278783
rect 416881 280109 416915 280143
rect 397653 278545 397687 278579
rect 382473 270521 382507 270555
rect 386613 273241 386647 273275
rect 356437 270453 356471 270487
rect 295441 263449 295475 263483
rect 309333 270385 309367 270419
rect 381093 270385 381127 270419
rect 309333 260865 309367 260899
rect 324421 263585 324455 263619
rect 324421 260865 324455 260899
rect 342545 263585 342579 263619
rect 342545 260865 342579 260899
rect 386613 269161 386647 269195
rect 416881 270521 416915 270555
rect 433625 280109 433659 280143
rect 466561 280109 466595 280143
rect 433625 270521 433659 270555
rect 451565 273717 451599 273751
rect 397653 269093 397687 269127
rect 400505 270453 400539 270487
rect 381093 260865 381127 260899
rect 386521 264265 386555 264299
rect 292681 260729 292715 260763
rect 294153 260797 294187 260831
rect 288633 251209 288667 251243
rect 294153 251209 294187 251243
rect 295533 260797 295567 260831
rect 295533 251209 295567 251243
rect 305193 260797 305227 260831
rect 310713 260797 310747 260831
rect 305193 251209 305227 251243
rect 309333 260729 309367 260763
rect 309333 251209 309367 251243
rect 310713 251209 310747 251243
rect 321753 260797 321787 260831
rect 321753 251209 321787 251243
rect 327273 260797 327307 260831
rect 334357 260797 334391 260831
rect 346593 260797 346627 260831
rect 334357 251277 334391 251311
rect 342453 260729 342487 260763
rect 327273 251209 327307 251243
rect 342453 251209 342487 251243
rect 382473 260797 382507 260831
rect 346593 251209 346627 251243
rect 370053 253997 370087 254031
rect 259653 248489 259687 248523
rect 292773 251141 292807 251175
rect 236285 244341 236319 244375
rect 254133 248353 254167 248387
rect 236285 244205 236319 244239
rect 254133 244205 254167 244239
rect 334357 251141 334391 251175
rect 324421 244273 324455 244307
rect 353585 251141 353619 251175
rect 334357 244137 334391 244171
rect 348065 250053 348099 250087
rect 324421 241553 324455 241587
rect 348065 241485 348099 241519
rect 370053 248489 370087 248523
rect 375573 253997 375607 254031
rect 386521 259437 386555 259471
rect 392041 264265 392075 264299
rect 466561 270521 466595 270555
rect 472081 280109 472115 280143
rect 472081 270521 472115 270555
rect 451565 263449 451599 263483
rect 400505 260865 400539 260899
rect 392041 259437 392075 259471
rect 416881 260797 416915 260831
rect 382473 251209 382507 251243
rect 397561 253929 397595 253963
rect 416881 251209 416915 251243
rect 433625 260797 433659 260831
rect 466561 260797 466595 260831
rect 433625 251209 433659 251243
rect 451565 259369 451599 259403
rect 397561 249781 397595 249815
rect 400505 251141 400539 251175
rect 375573 248489 375607 248523
rect 375573 248353 375607 248387
rect 375573 242777 375607 242811
rect 397561 244953 397595 244987
rect 353585 241485 353619 241519
rect 292773 240125 292807 240159
rect 466561 251209 466595 251243
rect 472081 260797 472115 260831
rect 472081 251209 472115 251243
rect 451565 244137 451599 244171
rect 400505 241485 400539 241519
rect 397561 240125 397595 240159
rect 236285 234617 236319 234651
rect 292773 239989 292807 240023
rect 259653 231761 259687 231795
rect 236285 224825 236319 224859
rect 331321 231829 331355 231863
rect 292773 230469 292807 230503
rect 309333 231761 309367 231795
rect 259653 222173 259687 222207
rect 281733 229041 281767 229075
rect 236285 215305 236319 215339
rect 243093 222037 243127 222071
rect 243093 212517 243127 212551
rect 270693 215373 270727 215407
rect 259653 212449 259687 212483
rect 270693 212449 270727 212483
rect 331321 227749 331355 227783
rect 309333 222173 309367 222207
rect 451289 224961 451323 224995
rect 451289 222173 451323 222207
rect 281733 212449 281767 212483
rect 334357 219385 334391 219419
rect 408785 215305 408819 215339
rect 364349 212789 364383 212823
rect 334357 212449 334391 212483
rect 364165 212517 364199 212551
rect 243185 205649 243219 205683
rect 243185 202861 243219 202895
rect 270693 211089 270727 211123
rect 259653 202861 259687 202895
rect 265265 205649 265299 205683
rect 270693 205581 270727 205615
rect 295533 209729 295567 209763
rect 265265 202861 265299 202895
rect 408785 212517 408819 212551
rect 364349 212381 364383 212415
rect 369961 212449 369995 212483
rect 364165 208369 364199 208403
rect 336841 205649 336875 205683
rect 336841 202861 336875 202895
rect 369961 202861 369995 202895
rect 480269 202929 480303 202963
rect 295533 202793 295567 202827
rect 243093 202725 243127 202759
rect 480269 201501 480303 201535
rect 281917 201433 281951 201467
rect 243093 193205 243127 193239
rect 255513 200073 255547 200107
rect 270601 196061 270635 196095
rect 270601 193137 270635 193171
rect 309333 201433 309367 201467
rect 281917 193137 281951 193171
rect 295717 200073 295751 200107
rect 255513 190485 255547 190519
rect 270601 191777 270635 191811
rect 236285 187561 236319 187595
rect 271981 186405 272015 186439
rect 271981 183549 272015 183583
rect 270601 183481 270635 183515
rect 298293 186405 298327 186439
rect 298293 183549 298327 183583
rect 352113 201433 352147 201467
rect 332793 198645 332827 198679
rect 369961 201433 369995 201467
rect 352113 193137 352147 193171
rect 359197 197285 359231 197319
rect 332793 189057 332827 189091
rect 386613 198645 386647 198679
rect 375573 196061 375607 196095
rect 375573 193205 375607 193239
rect 369961 193137 369995 193171
rect 359197 187697 359231 187731
rect 364533 190417 364567 190451
rect 309333 183549 309367 183583
rect 321661 186405 321695 186439
rect 321661 183549 321695 183583
rect 324421 186405 324455 186439
rect 324421 183549 324455 183583
rect 357633 186405 357667 186439
rect 295717 183481 295751 183515
rect 267197 182121 267231 182155
rect 255513 180761 255547 180795
rect 236285 178041 236319 178075
rect 252753 178789 252787 178823
rect 252753 173893 252787 173927
rect 254133 172465 254167 172499
rect 243001 167093 243035 167127
rect 254133 166957 254167 166991
rect 336841 182121 336875 182155
rect 336841 176545 336875 176579
rect 347973 180761 348007 180795
rect 267197 173281 267231 173315
rect 255513 166957 255547 166991
rect 259653 172465 259687 172499
rect 243001 162877 243035 162911
rect 271981 172465 272015 172499
rect 259653 162877 259687 162911
rect 265173 164169 265207 164203
rect 292773 172465 292807 172499
rect 292773 164169 292807 164203
rect 342361 172465 342395 172499
rect 271981 162877 272015 162911
rect 342361 162877 342395 162911
rect 347973 162877 348007 162911
rect 352113 180761 352147 180795
rect 352113 162877 352147 162911
rect 353493 180761 353527 180795
rect 364533 186269 364567 186303
rect 433717 196061 433751 196095
rect 433717 193205 433751 193239
rect 386613 186269 386647 186303
rect 357633 179401 357667 179435
rect 397745 176613 397779 176647
rect 397745 173893 397779 173927
rect 382473 167637 382507 167671
rect 353493 162877 353527 162911
rect 370053 164169 370087 164203
rect 298293 162809 298327 162843
rect 265173 154649 265207 154683
rect 271981 157981 272015 158015
rect 243001 154513 243035 154547
rect 236377 151725 236411 151759
rect 243001 147577 243035 147611
rect 254409 153085 254443 153119
rect 298293 157301 298327 157335
rect 334541 161381 334575 161415
rect 271981 148597 272015 148631
rect 292773 155873 292807 155907
rect 292773 147577 292807 147611
rect 331413 154513 331447 154547
rect 334541 153153 334575 153187
rect 356437 161313 356471 161347
rect 370053 154581 370087 154615
rect 376953 164169 376987 164203
rect 376953 154581 376987 154615
rect 397745 164169 397779 164203
rect 382473 154581 382507 154615
rect 393237 162809 393271 162843
rect 356437 151793 356471 151827
rect 375573 154513 375607 154547
rect 331413 147441 331447 147475
rect 334449 151725 334483 151759
rect 254409 143565 254443 143599
rect 292773 144857 292807 144891
rect 236377 143429 236411 143463
rect 254225 143497 254259 143531
rect 243277 133841 243311 133875
rect 243277 124185 243311 124219
rect 259653 143497 259687 143531
rect 287253 143497 287287 143531
rect 259653 133773 259687 133807
rect 283021 142069 283055 142103
rect 292773 135269 292807 135303
rect 305101 143497 305135 143531
rect 287253 133909 287287 133943
rect 321661 143497 321695 143531
rect 375573 147577 375607 147611
rect 381093 154513 381127 154547
rect 381093 147577 381127 147611
rect 392133 154513 392167 154547
rect 392133 147577 392167 147611
rect 400505 164169 400539 164203
rect 400505 157301 400539 157335
rect 422401 164169 422435 164203
rect 466561 164169 466595 164203
rect 422401 157301 422435 157335
rect 451565 162809 451599 162843
rect 397745 154581 397779 154615
rect 466561 157301 466595 157335
rect 480269 164169 480303 164203
rect 480269 153221 480303 153255
rect 451565 147577 451599 147611
rect 393237 144993 393271 145027
rect 397745 144925 397779 144959
rect 334449 142137 334483 142171
rect 381093 144789 381127 144823
rect 397745 143565 397779 143599
rect 400505 144857 400539 144891
rect 381093 135269 381127 135303
rect 393237 143497 393271 143531
rect 321661 135201 321695 135235
rect 305101 133909 305135 133943
rect 400505 137921 400539 137955
rect 422401 144857 422435 144891
rect 422401 137921 422435 137955
rect 466561 144857 466595 144891
rect 466561 137921 466595 137955
rect 393237 133909 393271 133943
rect 283021 132481 283055 132515
rect 292773 133841 292807 133875
rect 254225 124185 254259 124219
rect 267197 132413 267231 132447
rect 240149 124117 240183 124151
rect 240149 114529 240183 114563
rect 249993 124117 250027 124151
rect 334449 133841 334483 133875
rect 292773 125545 292807 125579
rect 304917 125681 304951 125715
rect 304917 124185 304951 124219
rect 310713 125545 310747 125579
rect 267197 122825 267231 122859
rect 271981 124117 272015 124151
rect 249993 114529 250027 114563
rect 252753 119357 252787 119391
rect 236285 113101 236319 113135
rect 243093 109701 243127 109735
rect 236285 103513 236319 103547
rect 240149 106233 240183 106267
rect 271981 115345 272015 115379
rect 287161 124117 287195 124151
rect 287161 114529 287195 114563
rect 292865 124117 292899 124151
rect 292865 113169 292899 113203
rect 298201 118745 298235 118779
rect 252753 106301 252787 106335
rect 295533 113101 295567 113135
rect 243093 106165 243127 106199
rect 281641 106233 281675 106267
rect 240149 96645 240183 96679
rect 254225 103445 254259 103479
rect 236285 95149 236319 95183
rect 240149 95149 240183 95183
rect 254225 93857 254259 93891
rect 266461 102085 266495 102119
rect 281641 101337 281675 101371
rect 282929 104805 282963 104839
rect 334449 124185 334483 124219
rect 353493 133841 353527 133875
rect 353493 124185 353527 124219
rect 356437 133841 356471 133875
rect 386613 133841 386647 133875
rect 356437 124185 356471 124219
rect 381185 125545 381219 125579
rect 342637 124117 342671 124151
rect 327273 122757 327307 122791
rect 310713 118609 310747 118643
rect 321753 118813 321787 118847
rect 298201 111809 298235 111843
rect 305101 115889 305135 115923
rect 295533 103513 295567 103547
rect 298385 111673 298419 111707
rect 321753 114529 321787 114563
rect 324513 118813 324547 118847
rect 324513 114529 324547 114563
rect 327273 113169 327307 113203
rect 330033 120241 330067 120275
rect 305101 106301 305135 106335
rect 365913 124117 365947 124151
rect 365913 118609 365947 118643
rect 433625 125545 433659 125579
rect 386613 122893 386647 122927
rect 407773 124117 407807 124151
rect 381185 115957 381219 115991
rect 386889 121397 386923 121431
rect 342637 114529 342671 114563
rect 348065 114529 348099 114563
rect 348065 113169 348099 113203
rect 330033 106301 330067 106335
rect 324513 106233 324547 106267
rect 298385 102153 298419 102187
rect 309241 104805 309275 104839
rect 298385 99433 298419 99467
rect 288633 99365 288667 99399
rect 288633 96645 288667 96679
rect 282929 95217 282963 95251
rect 266461 92497 266495 92531
rect 287161 95149 287195 95183
rect 240149 85629 240183 85663
rect 241805 86921 241839 86955
rect 236285 85561 236319 85595
rect 236285 85425 236319 85459
rect 308137 99365 308171 99399
rect 308137 96645 308171 96679
rect 298385 93789 298419 93823
rect 294153 93653 294187 93687
rect 287161 85629 287195 85663
rect 288633 86921 288667 86955
rect 249993 85493 250027 85527
rect 241805 77265 241839 77299
rect 243185 80733 243219 80767
rect 236285 75905 236319 75939
rect 249993 79305 250027 79339
rect 254133 85493 254167 85527
rect 243185 67609 243219 67643
rect 244473 70465 244507 70499
rect 244473 67609 244507 67643
rect 287253 85493 287287 85527
rect 259653 84133 259687 84167
rect 255513 79985 255547 80019
rect 255513 74545 255547 74579
rect 271981 82773 272015 82807
rect 259653 71077 259687 71111
rect 266461 77945 266495 77979
rect 254133 67609 254167 67643
rect 270693 75837 270727 75871
rect 281733 77265 281767 77299
rect 281733 75905 281767 75939
rect 319085 104805 319119 104839
rect 310713 99365 310747 99399
rect 310713 96645 310747 96679
rect 357633 106233 357667 106267
rect 324513 96645 324547 96679
rect 353493 103445 353527 103479
rect 319085 95217 319119 95251
rect 433625 115957 433659 115991
rect 466653 124117 466687 124151
rect 407773 114529 407807 114563
rect 466653 114529 466687 114563
rect 397653 114461 397687 114495
rect 397653 104941 397687 104975
rect 408693 114461 408727 114495
rect 408693 104873 408727 104907
rect 422401 106233 422435 106267
rect 386889 103513 386923 103547
rect 393145 104805 393179 104839
rect 393145 98685 393179 98719
rect 400505 104805 400539 104839
rect 357633 96509 357667 96543
rect 400505 95217 400539 95251
rect 407773 104805 407807 104839
rect 353493 93857 353527 93891
rect 309241 89641 309275 89675
rect 364533 93789 364567 93823
rect 294153 84201 294187 84235
rect 298569 88961 298603 88995
rect 298569 84201 298603 84235
rect 305193 86921 305227 86955
rect 288633 77265 288667 77299
rect 305193 77265 305227 77299
rect 308137 86921 308171 86955
rect 310713 86921 310747 86955
rect 308137 77265 308171 77299
rect 309333 80053 309367 80087
rect 309333 77265 309367 77299
rect 342545 86921 342579 86955
rect 334265 85493 334299 85527
rect 342545 79985 342579 80019
rect 346593 86921 346627 86955
rect 375573 93517 375607 93551
rect 381001 89777 381035 89811
rect 381001 86989 381035 87023
rect 408785 100045 408819 100079
rect 422401 99297 422435 99331
rect 427921 106233 427955 106267
rect 427921 99297 427955 99331
rect 433625 106233 433659 106267
rect 433625 99297 433659 99331
rect 480453 104805 480487 104839
rect 480453 95217 480487 95251
rect 408785 89641 408819 89675
rect 407773 86989 407807 87023
rect 375573 85561 375607 85595
rect 382473 86921 382507 86955
rect 364533 84201 364567 84235
rect 381001 85493 381035 85527
rect 357725 84133 357759 84167
rect 346593 79985 346627 80019
rect 356437 82773 356471 82807
rect 334265 79305 334299 79339
rect 310713 77265 310747 77299
rect 352021 77333 352055 77367
rect 287253 75905 287287 75939
rect 271981 73185 272015 73219
rect 334357 74477 334391 74511
rect 305193 70465 305227 70499
rect 305193 67609 305227 67643
rect 270693 66249 270727 66283
rect 281733 67541 281767 67575
rect 266461 64889 266495 64923
rect 249901 64821 249935 64855
rect 240241 56525 240275 56559
rect 249901 56525 249935 56559
rect 255513 64821 255547 64855
rect 281733 61421 281767 61455
rect 283113 66181 283147 66215
rect 287253 66181 287287 66215
rect 287253 56661 287287 56695
rect 292773 66181 292807 66215
rect 283113 56593 283147 56627
rect 255513 55233 255547 55267
rect 281641 56525 281675 56559
rect 267013 55097 267047 55131
rect 249901 51153 249935 51187
rect 249901 47005 249935 47039
rect 240241 46937 240275 46971
rect 231961 46869 231995 46903
rect 231961 37281 231995 37315
rect 236285 46869 236319 46903
rect 236285 37281 236319 37315
rect 244473 46869 244507 46903
rect 244473 37281 244507 37315
rect 249901 46869 249935 46903
rect 271981 51765 272015 51799
rect 271981 46937 272015 46971
rect 287253 56525 287287 56559
rect 287253 47005 287287 47039
rect 324513 66181 324547 66215
rect 310621 64821 310655 64855
rect 359013 84133 359047 84167
rect 359013 77945 359047 77979
rect 381001 75905 381035 75939
rect 422401 86921 422435 86955
rect 382473 75905 382507 75939
rect 407773 85493 407807 85527
rect 408693 85493 408727 85527
rect 466469 85493 466503 85527
rect 422401 77265 422435 77299
rect 433625 80189 433659 80223
rect 433625 77265 433659 77299
rect 466469 77129 466503 77163
rect 472081 85493 472115 85527
rect 408693 75973 408727 76007
rect 427921 76313 427955 76347
rect 407773 75905 407807 75939
rect 357725 74545 357759 74579
rect 375573 75837 375607 75871
rect 356437 73185 356471 73219
rect 364533 74477 364567 74511
rect 352021 66249 352055 66283
rect 334357 64957 334391 64991
rect 408693 75837 408727 75871
rect 375573 66317 375607 66351
rect 381093 67541 381127 67575
rect 364533 64889 364567 64923
rect 375481 66181 375515 66215
rect 324513 56593 324547 56627
rect 331413 64821 331447 64855
rect 310621 55233 310655 55267
rect 329941 55165 329975 55199
rect 292773 47005 292807 47039
rect 321753 51153 321787 51187
rect 321753 47005 321787 47039
rect 281641 46937 281675 46971
rect 331413 48297 331447 48331
rect 334357 64821 334391 64855
rect 356529 63461 356563 63495
rect 334357 48297 334391 48331
rect 342453 55165 342487 55199
rect 329941 46937 329975 46971
rect 267013 45577 267047 45611
rect 309333 46869 309367 46903
rect 282929 45509 282963 45543
rect 272073 42925 272107 42959
rect 267105 42041 267139 42075
rect 249901 37281 249935 37315
rect 252753 40137 252787 40171
rect 231869 35853 231903 35887
rect 240241 31841 240275 31875
rect 252753 31637 252787 31671
rect 267105 28985 267139 29019
rect 282929 35921 282963 35955
rect 292865 45509 292899 45543
rect 342453 45577 342487 45611
rect 359197 63461 359231 63495
rect 427921 67609 427955 67643
rect 480453 85493 480487 85527
rect 480453 77129 480487 77163
rect 472081 67609 472115 67643
rect 408693 66249 408727 66283
rect 381093 57953 381127 57987
rect 407773 66181 407807 66215
rect 375481 56593 375515 56627
rect 407773 56593 407807 56627
rect 416881 57885 416915 57919
rect 397745 56525 397779 56559
rect 359197 53805 359231 53839
rect 375573 56457 375607 56491
rect 375573 51697 375607 51731
rect 382381 51085 382415 51119
rect 356529 45577 356563 45611
rect 359105 48365 359139 48399
rect 382381 48297 382415 48331
rect 359105 45577 359139 45611
rect 392133 48229 392167 48263
rect 353585 45509 353619 45543
rect 330033 44081 330067 44115
rect 309333 37281 309367 37315
rect 324513 40137 324547 40171
rect 292865 35921 292899 35955
rect 272073 28985 272107 29019
rect 324513 28985 324547 29019
rect 240241 26333 240275 26367
rect 252845 28917 252879 28951
rect 231869 26265 231903 26299
rect 236377 26197 236411 26231
rect 236377 16609 236411 16643
rect 244289 19397 244323 19431
rect 281733 28917 281767 28951
rect 252845 19329 252879 19363
rect 266645 27557 266679 27591
rect 266645 19193 266679 19227
rect 270693 27557 270727 27591
rect 281733 19329 281767 19363
rect 318993 27557 319027 27591
rect 270693 17969 270727 18003
rect 288541 19261 288575 19295
rect 244289 16609 244323 16643
rect 252753 12529 252787 12563
rect 252753 11713 252787 11747
rect 305101 19261 305135 19295
rect 305101 13413 305135 13447
rect 308045 19261 308079 19295
rect 293969 12461 294003 12495
rect 293969 11849 294003 11883
rect 288541 10693 288575 10727
rect 318993 17969 319027 18003
rect 324421 27557 324455 27591
rect 357541 41429 357575 41463
rect 353585 37213 353619 37247
rect 356621 40749 356655 40783
rect 356621 35921 356655 35955
rect 357541 35921 357575 35955
rect 416881 48365 416915 48399
rect 433625 57885 433659 57919
rect 433625 48297 433659 48331
rect 466561 57885 466595 57919
rect 466561 48297 466595 48331
rect 472081 57885 472115 57919
rect 472081 48297 472115 48331
rect 397745 46937 397779 46971
rect 400597 47141 400631 47175
rect 400597 45577 400631 45611
rect 407773 46869 407807 46903
rect 400689 45441 400723 45475
rect 407773 37281 407807 37315
rect 472173 38573 472207 38607
rect 400689 37145 400723 37179
rect 392133 35921 392167 35955
rect 330033 26265 330067 26299
rect 342361 32385 342395 32419
rect 472173 31161 472207 31195
rect 356529 31093 356563 31127
rect 342361 19329 342395 19363
rect 346501 27557 346535 27591
rect 324421 17969 324455 18003
rect 427829 28917 427863 28951
rect 356529 26333 356563 26367
rect 393237 27557 393271 27591
rect 347881 26197 347915 26231
rect 347881 19397 347915 19431
rect 357541 26197 357575 26231
rect 346501 17969 346535 18003
rect 308045 10081 308079 10115
rect 330125 17901 330159 17935
rect 334357 17901 334391 17935
rect 334357 11305 334391 11339
rect 364809 26197 364843 26231
rect 364809 17425 364843 17459
rect 392225 26197 392259 26231
rect 407773 27557 407807 27591
rect 393237 17969 393271 18003
rect 397561 19261 397595 19295
rect 392225 16609 392259 16643
rect 382381 13073 382415 13107
rect 357541 9809 357575 9843
rect 376861 9945 376895 9979
rect 330125 9469 330159 9503
rect 346501 9605 346535 9639
rect 346501 8449 346535 8483
rect 369961 9605 369995 9639
rect 369961 8245 369995 8279
rect 371249 9605 371283 9639
rect 315221 6749 315255 6783
rect 376861 6273 376895 6307
rect 371249 6069 371283 6103
rect 315221 5865 315255 5899
rect 322213 6001 322247 6035
rect 322213 5797 322247 5831
rect 397561 9673 397595 9707
rect 480361 27557 480395 27591
rect 427829 19397 427863 19431
rect 472173 22253 472207 22287
rect 472173 19329 472207 19363
rect 407773 9673 407807 9707
rect 427829 19261 427863 19295
rect 480361 17969 480395 18003
rect 427829 9673 427863 9707
rect 382381 5321 382415 5355
rect 393053 9605 393087 9639
rect 392961 4029 392995 4063
rect 282101 3689 282135 3723
rect 282193 3961 282227 3995
rect 282285 3961 282319 3995
rect 374653 3961 374687 3995
rect 282193 3689 282227 3723
rect 372813 3689 372847 3723
rect 238217 3621 238251 3655
rect 238217 3485 238251 3519
rect 276765 3553 276799 3587
rect 276765 3349 276799 3383
rect 292589 3553 292623 3587
rect 292589 3281 292623 3315
rect 302157 3485 302191 3519
rect 372813 3485 372847 3519
rect 372905 3485 372939 3519
rect 371525 3417 371559 3451
rect 302157 3281 302191 3315
rect 335185 3281 335219 3315
rect 82921 3145 82955 3179
rect 335185 3145 335219 3179
rect 372905 3145 372939 3179
rect 392961 3893 392995 3927
rect 374653 3077 374687 3111
rect 82921 2941 82955 2975
rect 98653 2941 98687 2975
rect 371525 2941 371559 2975
rect 121469 2873 121503 2907
rect 121653 2873 121687 2907
rect 98653 2805 98687 2839
rect 406301 4233 406335 4267
rect 393973 4097 394007 4131
rect 393881 4029 393915 4063
rect 393973 3825 394007 3859
rect 403541 4097 403575 4131
rect 403541 3825 403575 3859
rect 403633 3961 403667 3995
rect 403633 3689 403667 3723
rect 403725 3689 403759 3723
rect 393881 3349 393915 3383
rect 403633 3349 403667 3383
rect 403817 3417 403851 3451
rect 409245 4097 409279 4131
rect 408325 4029 408359 4063
rect 423689 4097 423723 4131
rect 409245 3961 409279 3995
rect 416237 4029 416271 4063
rect 408417 3621 408451 3655
rect 408509 3621 408543 3655
rect 406301 3349 406335 3383
rect 403909 3281 403943 3315
rect 516977 4029 517011 4063
rect 432705 3961 432739 3995
rect 423689 3621 423723 3655
rect 423781 3621 423815 3655
rect 409889 3417 409923 3451
rect 416237 3417 416271 3451
rect 418169 3553 418203 3587
rect 409613 3349 409647 3383
rect 403541 3077 403575 3111
rect 403633 3213 403667 3247
rect 403725 3213 403759 3247
rect 408509 3213 408543 3247
rect 408601 3213 408635 3247
rect 403633 3077 403667 3111
rect 408785 3077 408819 3111
rect 410717 3077 410751 3111
rect 408509 2873 408543 2907
rect 423781 3485 423815 3519
rect 426725 3621 426759 3655
rect 421941 3349 421975 3383
rect 421113 3213 421147 3247
rect 421941 3145 421975 3179
rect 422953 3281 422987 3315
rect 422953 3009 422987 3043
rect 421113 2941 421147 2975
rect 418169 2873 418203 2907
rect 509801 3825 509835 3859
rect 432705 3281 432739 3315
rect 447609 3349 447643 3383
rect 509801 3281 509835 3315
rect 447609 3213 447643 3247
rect 569141 3485 569175 3519
rect 569141 3349 569175 3383
rect 516977 3213 517011 3247
rect 540161 3281 540195 3315
rect 540161 3009 540195 3043
rect 426725 2873 426759 2907
rect 393053 561 393087 595
<< metal1 >>
rect 218974 700952 218980 701004
rect 219032 700992 219038 701004
rect 393314 700992 393320 701004
rect 219032 700964 393320 700992
rect 219032 700952 219038 700964
rect 393314 700952 393320 700964
rect 393372 700952 393378 701004
rect 355962 700884 355968 700936
rect 356020 700924 356026 700936
rect 543458 700924 543464 700936
rect 356020 700896 543464 700924
rect 356020 700884 356026 700896
rect 543458 700884 543464 700896
rect 543516 700884 543522 700936
rect 202782 700816 202788 700868
rect 202840 700856 202846 700868
rect 390554 700856 390560 700868
rect 202840 700828 390560 700856
rect 202840 700816 202846 700828
rect 390554 700816 390560 700828
rect 390612 700816 390618 700868
rect 170306 700748 170312 700800
rect 170364 700788 170370 700800
rect 396074 700788 396080 700800
rect 170364 700760 396080 700788
rect 170364 700748 170370 700760
rect 396074 700748 396080 700760
rect 396132 700748 396138 700800
rect 154114 700680 154120 700732
rect 154172 700720 154178 700732
rect 401594 700720 401600 700732
rect 154172 700692 401600 700720
rect 154172 700680 154178 700692
rect 401594 700680 401600 700692
rect 401652 700680 401658 700732
rect 137830 700612 137836 700664
rect 137888 700652 137894 700664
rect 398834 700652 398840 700664
rect 137888 700624 398840 700652
rect 137888 700612 137894 700624
rect 398834 700612 398840 700624
rect 398892 700612 398898 700664
rect 105446 700544 105452 700596
rect 105504 700584 105510 700596
rect 404354 700584 404360 700596
rect 105504 700556 404360 700584
rect 105504 700544 105510 700556
rect 404354 700544 404360 700556
rect 404412 700544 404418 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 409874 700516 409880 700528
rect 89220 700488 409880 700516
rect 89220 700476 89226 700488
rect 409874 700476 409880 700488
rect 409932 700476 409938 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 407114 700448 407120 700460
rect 73028 700420 407120 700448
rect 73028 700408 73034 700420
rect 407114 700408 407120 700420
rect 407172 700408 407178 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 411254 700380 411260 700392
rect 40552 700352 411260 700380
rect 40552 700340 40558 700352
rect 411254 700340 411260 700352
rect 411312 700340 411318 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 416774 700312 416780 700324
rect 24360 700284 416780 700312
rect 24360 700272 24366 700284
rect 416774 700272 416780 700284
rect 416832 700272 416838 700324
rect 353202 700204 353208 700256
rect 353260 700244 353266 700256
rect 527174 700244 527180 700256
rect 353260 700216 527180 700244
rect 353260 700204 353266 700216
rect 527174 700204 527180 700216
rect 527232 700204 527238 700256
rect 267642 700136 267648 700188
rect 267700 700176 267706 700188
rect 383654 700176 383660 700188
rect 267700 700148 383660 700176
rect 267700 700136 267706 700148
rect 383654 700136 383660 700148
rect 383712 700136 383718 700188
rect 362862 700068 362868 700120
rect 362920 700108 362926 700120
rect 478506 700108 478512 700120
rect 362920 700080 478512 700108
rect 362920 700068 362926 700080
rect 478506 700068 478512 700080
rect 478564 700068 478570 700120
rect 360102 700000 360108 700052
rect 360160 700040 360166 700052
rect 462314 700040 462320 700052
rect 360160 700012 462320 700040
rect 360160 700000 360166 700012
rect 462314 700000 462320 700012
rect 462372 700000 462378 700052
rect 283834 699932 283840 699984
rect 283892 699972 283898 699984
rect 385034 699972 385040 699984
rect 283892 699944 385040 699972
rect 283892 699932 283898 699944
rect 385034 699932 385040 699944
rect 385092 699932 385098 699984
rect 332502 699864 332508 699916
rect 332560 699904 332566 699916
rect 375374 699904 375380 699916
rect 332560 699876 375380 699904
rect 332560 699864 332566 699876
rect 375374 699864 375380 699876
rect 375432 699864 375438 699916
rect 371142 699796 371148 699848
rect 371200 699836 371206 699848
rect 413646 699836 413652 699848
rect 371200 699808 413652 699836
rect 371200 699796 371206 699808
rect 413646 699796 413652 699808
rect 413704 699796 413710 699848
rect 348786 699728 348792 699780
rect 348844 699768 348850 699780
rect 378134 699768 378140 699780
rect 348844 699740 378140 699768
rect 348844 699728 348850 699740
rect 378134 699728 378140 699740
rect 378192 699728 378198 699780
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 364978 699660 364984 699712
rect 365036 699700 365042 699712
rect 365622 699700 365628 699712
rect 365036 699672 365628 699700
rect 365036 699660 365042 699672
rect 365622 699660 365628 699672
rect 365680 699660 365686 699712
rect 368382 699660 368388 699712
rect 368440 699700 368446 699712
rect 397454 699700 397460 699712
rect 368440 699672 397460 699700
rect 368440 699660 368446 699672
rect 397454 699660 397460 699672
rect 397512 699660 397518 699712
rect 344922 696940 344928 696992
rect 344980 696980 344986 696992
rect 580166 696980 580172 696992
rect 344980 696952 580172 696980
rect 344980 696940 344986 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 429378 688576 429384 688628
rect 429436 688616 429442 688628
rect 429838 688616 429844 688628
rect 429436 688588 429844 688616
rect 429436 688576 429442 688588
rect 429838 688576 429844 688588
rect 429896 688576 429902 688628
rect 559098 688576 559104 688628
rect 559156 688616 559162 688628
rect 559650 688616 559656 688628
rect 559156 688588 559656 688616
rect 559156 688576 559162 688588
rect 559650 688576 559656 688588
rect 559708 688576 559714 688628
rect 429212 685936 429976 685964
rect 347682 685856 347688 685908
rect 347740 685896 347746 685908
rect 429212 685896 429240 685936
rect 347740 685868 429240 685896
rect 429948 685896 429976 685936
rect 552584 685936 559788 685964
rect 552584 685896 552612 685936
rect 429948 685868 552612 685896
rect 559760 685896 559788 685936
rect 580166 685896 580172 685908
rect 559760 685868 580172 685896
rect 347740 685856 347746 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 429286 684428 429292 684480
rect 429344 684468 429350 684480
rect 429565 684471 429623 684477
rect 429565 684468 429577 684471
rect 429344 684440 429577 684468
rect 429344 684428 429350 684440
rect 429565 684437 429577 684440
rect 429611 684437 429623 684471
rect 429565 684431 429623 684437
rect 559006 684428 559012 684480
rect 559064 684468 559070 684480
rect 559285 684471 559343 684477
rect 559285 684468 559297 684471
rect 559064 684440 559297 684468
rect 559064 684428 559070 684440
rect 559285 684437 559297 684440
rect 559331 684437 559343 684471
rect 559285 684431 559343 684437
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 419534 681748 419540 681760
rect 3568 681720 419540 681748
rect 3568 681708 3574 681720
rect 419534 681708 419540 681720
rect 419592 681708 419598 681760
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 342162 673480 342168 673532
rect 342220 673520 342226 673532
rect 580166 673520 580172 673532
rect 342220 673492 580172 673520
rect 342220 673480 342226 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 425054 667944 425060 667956
rect 3476 667916 425060 667944
rect 3476 667904 3482 667916
rect 425054 667904 425060 667916
rect 425112 667904 425118 667956
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 429470 656860 429476 656872
rect 429431 656832 429476 656860
rect 429470 656820 429476 656832
rect 429528 656820 429534 656872
rect 559190 656860 559196 656872
rect 559151 656832 559196 656860
rect 559190 656820 559196 656832
rect 559248 656820 559254 656872
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 422294 652780 422300 652792
rect 3108 652752 422300 652780
rect 3108 652740 3114 652752
rect 422294 652740 422300 652752
rect 422352 652740 422358 652792
rect 336642 650020 336648 650072
rect 336700 650060 336706 650072
rect 580166 650060 580172 650072
rect 336700 650032 580172 650060
rect 336700 650020 336706 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 429473 647275 429531 647281
rect 429473 647241 429485 647275
rect 429519 647272 429531 647275
rect 429562 647272 429568 647284
rect 429519 647244 429568 647272
rect 429519 647241 429531 647244
rect 429473 647235 429531 647241
rect 429562 647232 429568 647244
rect 429620 647232 429626 647284
rect 559193 647275 559251 647281
rect 559193 647241 559205 647275
rect 559239 647272 559251 647275
rect 559282 647272 559288 647284
rect 559239 647244 559288 647272
rect 559239 647241 559251 647244
rect 559193 647235 559251 647241
rect 559282 647232 559288 647244
rect 559340 647232 559346 647284
rect 365162 643968 365168 644020
rect 365220 644008 365226 644020
rect 429562 644008 429568 644020
rect 365220 643980 429568 644008
rect 365220 643968 365226 643980
rect 429562 643968 429568 643980
rect 429620 643968 429626 644020
rect 300762 643900 300768 643952
rect 300820 643940 300826 643952
rect 380986 643940 380992 643952
rect 300820 643912 380992 643940
rect 300820 643900 300826 643912
rect 380986 643900 380992 643912
rect 381044 643900 381050 643952
rect 357342 643832 357348 643884
rect 357400 643872 357406 643884
rect 494238 643872 494244 643884
rect 357400 643844 494244 643872
rect 357400 643832 357406 643844
rect 494238 643832 494244 643844
rect 494296 643832 494302 643884
rect 235902 643764 235908 643816
rect 235960 643804 235966 643816
rect 388898 643804 388904 643816
rect 235960 643776 388904 643804
rect 235960 643764 235966 643776
rect 388898 643764 388904 643776
rect 388956 643764 388962 643816
rect 349430 643696 349436 643748
rect 349488 643736 349494 643748
rect 559282 643736 559288 643748
rect 349488 643708 559288 643736
rect 349488 643696 349494 643708
rect 559282 643696 559288 643708
rect 559340 643696 559346 643748
rect 365622 643084 365628 643136
rect 365680 643124 365686 643136
rect 373074 643124 373080 643136
rect 365680 643096 373080 643124
rect 365680 643084 365686 643096
rect 373074 643084 373080 643096
rect 373132 643084 373138 643136
rect 331030 643016 331036 643068
rect 331088 643056 331094 643068
rect 530394 643056 530400 643068
rect 331088 643028 530400 643056
rect 331088 643016 331094 643028
rect 530394 643016 530400 643028
rect 530452 643016 530458 643068
rect 323118 642948 323124 643000
rect 323176 642988 323182 643000
rect 531222 642988 531228 643000
rect 323176 642960 531228 642988
rect 323176 642948 323182 642960
rect 531222 642948 531228 642960
rect 531280 642948 531286 643000
rect 315206 642880 315212 642932
rect 315264 642920 315270 642932
rect 531038 642920 531044 642932
rect 315264 642892 531044 642920
rect 315264 642880 315270 642892
rect 531038 642880 531044 642892
rect 531096 642880 531102 642932
rect 296806 642812 296812 642864
rect 296864 642852 296870 642864
rect 530762 642852 530768 642864
rect 296864 642824 530768 642852
rect 296864 642812 296870 642824
rect 530762 642812 530768 642824
rect 530820 642812 530826 642864
rect 309962 642744 309968 642796
rect 310020 642784 310026 642796
rect 580166 642784 580172 642796
rect 310020 642756 580172 642784
rect 310020 642744 310026 642756
rect 580166 642744 580172 642756
rect 580224 642744 580230 642796
rect 270494 642676 270500 642728
rect 270552 642716 270558 642728
rect 580442 642716 580448 642728
rect 270552 642688 580448 642716
rect 270552 642676 270558 642688
rect 580442 642676 580448 642688
rect 580500 642676 580506 642728
rect 5442 642608 5448 642660
rect 5500 642648 5506 642660
rect 433610 642648 433616 642660
rect 5500 642620 433616 642648
rect 5500 642608 5506 642620
rect 433610 642608 433616 642620
rect 433668 642608 433674 642660
rect 5350 642540 5356 642592
rect 5408 642580 5414 642592
rect 441522 642580 441528 642592
rect 5408 642552 441528 642580
rect 5408 642540 5414 642552
rect 441522 642540 441528 642552
rect 441580 642540 441586 642592
rect 3234 642472 3240 642524
rect 3292 642512 3298 642524
rect 438854 642512 438860 642524
rect 3292 642484 438860 642512
rect 3292 642472 3298 642484
rect 438854 642472 438860 642484
rect 438912 642472 438918 642524
rect 8018 642404 8024 642456
rect 8076 642444 8082 642456
rect 446766 642444 446772 642456
rect 8076 642416 446772 642444
rect 8076 642404 8082 642416
rect 446766 642404 446772 642416
rect 446824 642404 446830 642456
rect 5166 642336 5172 642388
rect 5224 642376 5230 642388
rect 449434 642376 449440 642388
rect 5224 642348 449440 642376
rect 5224 642336 5230 642348
rect 449434 642336 449440 642348
rect 449492 642336 449498 642388
rect 7926 642268 7932 642320
rect 7984 642308 7990 642320
rect 454678 642308 454684 642320
rect 7984 642280 454684 642308
rect 7984 642268 7990 642280
rect 454678 642268 454684 642280
rect 454736 642268 454742 642320
rect 3326 642200 3332 642252
rect 3384 642240 3390 642252
rect 459922 642240 459928 642252
rect 3384 642212 459928 642240
rect 3384 642200 3390 642212
rect 459922 642200 459928 642212
rect 459980 642200 459986 642252
rect 6362 642132 6368 642184
rect 6420 642172 6426 642184
rect 465166 642172 465172 642184
rect 6420 642144 465172 642172
rect 6420 642132 6426 642144
rect 465166 642132 465172 642144
rect 465224 642132 465230 642184
rect 4982 642064 4988 642116
rect 5040 642104 5046 642116
rect 470502 642104 470508 642116
rect 5040 642076 470508 642104
rect 5040 642064 5046 642076
rect 470502 642064 470508 642076
rect 470560 642064 470566 642116
rect 6270 641996 6276 642048
rect 6328 642036 6334 642048
rect 480990 642036 480996 642048
rect 6328 642008 480996 642036
rect 6328 641996 6334 642008
rect 480990 641996 480996 642008
rect 481048 641996 481054 642048
rect 4062 641928 4068 641980
rect 4120 641968 4126 641980
rect 486234 641968 486240 641980
rect 4120 641940 486240 641968
rect 4120 641928 4126 641940
rect 486234 641928 486240 641940
rect 486292 641928 486298 641980
rect 3970 641860 3976 641912
rect 4028 641900 4034 641912
rect 496814 641900 496820 641912
rect 4028 641872 496820 641900
rect 4028 641860 4034 641872
rect 496814 641860 496820 641872
rect 496872 641860 496878 641912
rect 3878 641792 3884 641844
rect 3936 641832 3942 641844
rect 502058 641832 502064 641844
rect 3936 641804 502064 641832
rect 3936 641792 3942 641804
rect 502058 641792 502064 641804
rect 502116 641792 502122 641844
rect 3786 641724 3792 641776
rect 3844 641764 3850 641776
rect 512546 641764 512552 641776
rect 3844 641736 512552 641764
rect 3844 641724 3850 641736
rect 512546 641724 512552 641736
rect 512604 641724 512610 641776
rect 320450 641112 320456 641164
rect 320508 641152 320514 641164
rect 530486 641152 530492 641164
rect 320508 641124 530492 641152
rect 320508 641112 320514 641124
rect 530486 641112 530492 641124
rect 530544 641112 530550 641164
rect 312538 641044 312544 641096
rect 312596 641084 312602 641096
rect 531130 641084 531136 641096
rect 312596 641056 531136 641084
rect 312596 641044 312602 641056
rect 531130 641044 531136 641056
rect 531188 641044 531194 641096
rect 302050 640976 302056 641028
rect 302108 641016 302114 641028
rect 530854 641016 530860 641028
rect 302108 640988 530860 641016
rect 302108 640976 302114 640988
rect 530854 640976 530860 640988
rect 530912 640976 530918 641028
rect 294138 640908 294144 640960
rect 294196 640948 294202 640960
rect 529566 640948 529572 640960
rect 294196 640920 529572 640948
rect 294196 640908 294202 640920
rect 529566 640908 529572 640920
rect 529624 640908 529630 640960
rect 286226 640840 286232 640892
rect 286284 640880 286290 640892
rect 529474 640880 529480 640892
rect 286284 640852 529480 640880
rect 286284 640840 286290 640852
rect 529474 640840 529480 640852
rect 529532 640840 529538 640892
rect 278314 640772 278320 640824
rect 278372 640812 278378 640824
rect 530578 640812 530584 640824
rect 278372 640784 530584 640812
rect 278372 640772 278378 640784
rect 530578 640772 530584 640784
rect 530636 640772 530642 640824
rect 265158 640704 265164 640756
rect 265216 640744 265222 640756
rect 580350 640744 580356 640756
rect 265216 640716 580356 640744
rect 265216 640704 265222 640716
rect 580350 640704 580356 640716
rect 580408 640704 580414 640756
rect 7834 640636 7840 640688
rect 7892 640676 7898 640688
rect 467834 640676 467840 640688
rect 7892 640648 467840 640676
rect 7892 640636 7898 640648
rect 467834 640636 467840 640648
rect 467892 640636 467898 640688
rect 7742 640568 7748 640620
rect 7800 640608 7806 640620
rect 475746 640608 475752 640620
rect 7800 640580 475752 640608
rect 7800 640568 7806 640580
rect 475746 640568 475752 640580
rect 475804 640568 475810 640620
rect 4798 640500 4804 640552
rect 4856 640540 4862 640552
rect 499390 640540 499396 640552
rect 4856 640512 499396 640540
rect 4856 640500 4862 640512
rect 499390 640500 499396 640512
rect 499448 640500 499454 640552
rect 6178 640432 6184 640484
rect 6236 640472 6242 640484
rect 507302 640472 507308 640484
rect 6236 640444 507308 640472
rect 6236 640432 6242 640444
rect 507302 640432 507308 640444
rect 507360 640432 507366 640484
rect 7650 640364 7656 640416
rect 7708 640404 7714 640416
rect 515214 640404 515220 640416
rect 7708 640376 515220 640404
rect 7708 640364 7714 640376
rect 515214 640364 515220 640376
rect 515272 640364 515278 640416
rect 7558 640296 7564 640348
rect 7616 640336 7622 640348
rect 523126 640336 523132 640348
rect 7616 640308 523132 640336
rect 7616 640296 7622 640308
rect 523126 640296 523132 640308
rect 523184 640296 523190 640348
rect 428090 639928 428096 639940
rect 428051 639900 428096 639928
rect 428090 639888 428096 639900
rect 428148 639888 428154 639940
rect 436094 639928 436100 639940
rect 436055 639900 436100 639928
rect 436094 639888 436100 639900
rect 436152 639888 436158 639940
rect 443822 639928 443828 639940
rect 443783 639900 443828 639928
rect 443822 639888 443828 639900
rect 443880 639888 443886 639940
rect 451734 639928 451740 639940
rect 451695 639900 451740 639928
rect 451734 639888 451740 639900
rect 451792 639888 451798 639940
rect 520274 639928 520280 639940
rect 520235 639900 520280 639928
rect 520274 639888 520280 639900
rect 520332 639888 520338 639940
rect 333882 639820 333888 639872
rect 333940 639860 333946 639872
rect 529750 639860 529756 639872
rect 333940 639832 529756 639860
rect 333940 639820 333946 639832
rect 529750 639820 529756 639832
rect 529808 639820 529814 639872
rect 325970 639752 325976 639804
rect 326028 639792 326034 639804
rect 529658 639792 529664 639804
rect 326028 639764 529664 639792
rect 326028 639752 326034 639764
rect 529658 639752 529664 639764
rect 529716 639752 529722 639804
rect 328454 639684 328460 639736
rect 328512 639724 328518 639736
rect 338022 639724 338028 639736
rect 328512 639696 338028 639724
rect 328512 639684 328518 639696
rect 338022 639684 338028 639696
rect 338080 639684 338086 639736
rect 339218 639684 339224 639736
rect 339276 639724 339282 639736
rect 579798 639724 579804 639736
rect 339276 639696 579804 639724
rect 339276 639684 339282 639696
rect 579798 639684 579804 639696
rect 579856 639684 579862 639736
rect 307570 639616 307576 639668
rect 307628 639656 307634 639668
rect 580902 639656 580908 639668
rect 307628 639628 580908 639656
rect 307628 639616 307634 639628
rect 580902 639616 580908 639628
rect 580960 639616 580966 639668
rect 299474 639548 299480 639600
rect 299532 639588 299538 639600
rect 580810 639588 580816 639600
rect 299532 639560 580816 639588
rect 299532 639548 299538 639560
rect 580810 639548 580816 639560
rect 580868 639548 580874 639600
rect 291746 639480 291752 639532
rect 291804 639520 291810 639532
rect 580718 639520 580724 639532
rect 291804 639492 580724 639520
rect 291804 639480 291810 639492
rect 580718 639480 580724 639492
rect 580776 639480 580782 639532
rect 284018 639412 284024 639464
rect 284076 639452 284082 639464
rect 580626 639452 580632 639464
rect 284076 639424 580632 639452
rect 284076 639412 284082 639424
rect 580626 639412 580632 639424
rect 580684 639412 580690 639464
rect 275922 639344 275928 639396
rect 275980 639384 275986 639396
rect 580534 639384 580540 639396
rect 275980 639356 580540 639384
rect 275980 639344 275986 639356
rect 580534 639344 580540 639356
rect 580592 639344 580598 639396
rect 268194 639276 268200 639328
rect 268252 639316 268258 639328
rect 580258 639316 580264 639328
rect 268252 639288 580264 639316
rect 268252 639276 268258 639288
rect 580258 639276 580264 639288
rect 580316 639276 580322 639328
rect 6730 639208 6736 639260
rect 6788 639248 6794 639260
rect 428093 639251 428151 639257
rect 428093 639248 428105 639251
rect 6788 639220 428105 639248
rect 6788 639208 6794 639220
rect 428093 639217 428105 639220
rect 428139 639217 428151 639251
rect 428093 639211 428151 639217
rect 6638 639140 6644 639192
rect 6696 639180 6702 639192
rect 436097 639183 436155 639189
rect 436097 639180 436109 639183
rect 6696 639152 436109 639180
rect 6696 639140 6702 639152
rect 436097 639149 436109 639152
rect 436143 639149 436155 639183
rect 436097 639143 436155 639149
rect 6546 639072 6552 639124
rect 6604 639112 6610 639124
rect 443825 639115 443883 639121
rect 443825 639112 443837 639115
rect 6604 639084 443837 639112
rect 6604 639072 6610 639084
rect 443825 639081 443837 639084
rect 443871 639081 443883 639115
rect 443825 639075 443883 639081
rect 6454 639004 6460 639056
rect 6512 639044 6518 639056
rect 451737 639047 451795 639053
rect 451737 639044 451749 639047
rect 6512 639016 451749 639044
rect 6512 639004 6518 639016
rect 451737 639013 451749 639016
rect 451783 639013 451795 639047
rect 451737 639007 451795 639013
rect 3602 638936 3608 638988
rect 3660 638976 3666 638988
rect 520277 638979 520335 638985
rect 520277 638976 520289 638979
rect 3660 638948 520289 638976
rect 3660 638936 3666 638948
rect 520277 638945 520289 638948
rect 520323 638945 520335 638979
rect 520277 638939 520335 638945
rect 529750 627852 529756 627904
rect 529808 627892 529814 627904
rect 580074 627892 580080 627904
rect 529808 627864 580080 627892
rect 529808 627852 529814 627864
rect 580074 627852 580080 627864
rect 580132 627852 580138 627904
rect 3142 624928 3148 624980
rect 3200 624968 3206 624980
rect 6730 624968 6736 624980
rect 3200 624940 6736 624968
rect 3200 624928 3206 624940
rect 6730 624928 6736 624940
rect 6788 624928 6794 624980
rect 2774 610512 2780 610564
rect 2832 610552 2838 610564
rect 5442 610552 5448 610564
rect 2832 610524 5448 610552
rect 2832 610512 2838 610524
rect 5442 610512 5448 610524
rect 5500 610512 5506 610564
rect 530302 604392 530308 604444
rect 530360 604432 530366 604444
rect 580074 604432 580080 604444
rect 530360 604404 580080 604432
rect 530360 604392 530366 604404
rect 580074 604392 580080 604404
rect 580132 604392 580138 604444
rect 3142 596028 3148 596080
rect 3200 596068 3206 596080
rect 8110 596068 8116 596080
rect 3200 596040 8116 596068
rect 3200 596028 3206 596040
rect 8110 596028 8116 596040
rect 8168 596028 8174 596080
rect 530394 593308 530400 593360
rect 530452 593348 530458 593360
rect 580074 593348 580080 593360
rect 530452 593320 580080 593348
rect 530452 593308 530458 593320
rect 580074 593308 580080 593320
rect 580132 593308 580138 593360
rect 529658 580932 529664 580984
rect 529716 580972 529722 580984
rect 580074 580972 580080 580984
rect 529716 580944 580080 580972
rect 529716 580932 529722 580944
rect 580074 580932 580080 580944
rect 580132 580932 580138 580984
rect 3142 567536 3148 567588
rect 3200 567576 3206 567588
rect 6638 567576 6644 567588
rect 3200 567548 6644 567576
rect 3200 567536 3206 567548
rect 6638 567536 6644 567548
rect 6696 567536 6702 567588
rect 530486 557472 530492 557524
rect 530544 557512 530550 557524
rect 580074 557512 580080 557524
rect 530544 557484 580080 557512
rect 530544 557472 530550 557484
rect 580074 557472 580080 557484
rect 580132 557472 580138 557524
rect 2774 553052 2780 553104
rect 2832 553092 2838 553104
rect 5350 553092 5356 553104
rect 2832 553064 5356 553092
rect 2832 553052 2838 553064
rect 5350 553052 5356 553064
rect 5408 553052 5414 553104
rect 531222 546388 531228 546440
rect 531280 546428 531286 546440
rect 580074 546428 580080 546440
rect 531280 546400 580080 546428
rect 531280 546388 531286 546400
rect 580074 546388 580080 546400
rect 580132 546388 580138 546440
rect 531130 510552 531136 510604
rect 531188 510592 531194 510604
rect 580074 510592 580080 510604
rect 531188 510564 580080 510592
rect 531188 510552 531194 510564
rect 580074 510552 580080 510564
rect 580132 510552 580138 510604
rect 3234 510348 3240 510400
rect 3292 510388 3298 510400
rect 6546 510388 6552 510400
rect 3292 510360 6552 510388
rect 3292 510348 3298 510360
rect 6546 510348 6552 510360
rect 6604 510348 6610 510400
rect 531038 499468 531044 499520
rect 531096 499508 531102 499520
rect 580074 499508 580080 499520
rect 531096 499480 580080 499508
rect 531096 499468 531102 499480
rect 580074 499468 580080 499480
rect 580132 499468 580138 499520
rect 2774 496408 2780 496460
rect 2832 496448 2838 496460
rect 5166 496448 5172 496460
rect 2832 496420 5172 496448
rect 2832 496408 2838 496420
rect 5166 496408 5172 496420
rect 5224 496408 5230 496460
rect 3234 481244 3240 481296
rect 3292 481284 3298 481296
rect 8018 481284 8024 481296
rect 3292 481256 8024 481284
rect 3292 481244 3298 481256
rect 8018 481244 8024 481256
rect 8076 481244 8082 481296
rect 530946 463632 530952 463684
rect 531004 463672 531010 463684
rect 579798 463672 579804 463684
rect 531004 463644 579804 463672
rect 531004 463632 531010 463644
rect 579798 463632 579804 463644
rect 579856 463632 579862 463684
rect 3142 452412 3148 452464
rect 3200 452452 3206 452464
rect 6454 452452 6460 452464
rect 3200 452424 6460 452452
rect 3200 452412 3206 452424
rect 6454 452412 6460 452424
rect 6512 452412 6518 452464
rect 530854 440172 530860 440224
rect 530912 440212 530918 440224
rect 580166 440212 580172 440224
rect 530912 440184 580172 440212
rect 530912 440172 530918 440184
rect 580166 440172 580172 440184
rect 580224 440172 580230 440224
rect 2774 437996 2780 438048
rect 2832 438036 2838 438048
rect 5258 438036 5264 438048
rect 2832 438008 5264 438036
rect 2832 437996 2838 438008
rect 5258 437996 5264 438008
rect 5316 437996 5322 438048
rect 3234 424260 3240 424312
rect 3292 424300 3298 424312
rect 7926 424300 7932 424312
rect 3292 424272 7932 424300
rect 3292 424260 3298 424272
rect 7926 424260 7932 424272
rect 7984 424260 7990 424312
rect 530762 416712 530768 416764
rect 530820 416752 530826 416764
rect 580166 416752 580172 416764
rect 530820 416724 580172 416752
rect 530820 416712 530826 416724
rect 580166 416712 580172 416724
rect 580224 416712 580230 416764
rect 529566 393252 529572 393304
rect 529624 393292 529630 393304
rect 579614 393292 579620 393304
rect 529624 393264 579620 393292
rect 529624 393252 529630 393264
rect 579614 393252 579620 393264
rect 579672 393252 579678 393304
rect 3234 380604 3240 380656
rect 3292 380644 3298 380656
rect 6362 380644 6368 380656
rect 3292 380616 6368 380644
rect 3292 380604 3298 380616
rect 6362 380604 6368 380616
rect 6420 380604 6426 380656
rect 2774 366732 2780 366784
rect 2832 366772 2838 366784
rect 5074 366772 5080 366784
rect 2832 366744 5080 366772
rect 2832 366732 2838 366744
rect 5074 366732 5080 366744
rect 5132 366732 5138 366784
rect 529658 346332 529664 346384
rect 529716 346372 529722 346384
rect 580166 346372 580172 346384
rect 529716 346344 580172 346372
rect 529716 346332 529722 346344
rect 580166 346332 580172 346344
rect 580224 346332 580230 346384
rect 356698 338376 356704 338428
rect 356756 338416 356762 338428
rect 357342 338416 357348 338428
rect 356756 338388 357348 338416
rect 356756 338376 356762 338388
rect 357342 338376 357348 338388
rect 357400 338376 357406 338428
rect 71038 338036 71044 338088
rect 71096 338076 71102 338088
rect 264882 338076 264888 338088
rect 71096 338048 264888 338076
rect 71096 338036 71102 338048
rect 264882 338036 264888 338048
rect 264940 338036 264946 338088
rect 332502 338036 332508 338088
rect 332560 338076 332566 338088
rect 400214 338076 400220 338088
rect 332560 338048 400220 338076
rect 332560 338036 332566 338048
rect 400214 338036 400220 338048
rect 400272 338036 400278 338088
rect 412082 338036 412088 338088
rect 412140 338076 412146 338088
rect 419166 338076 419172 338088
rect 412140 338048 419172 338076
rect 412140 338036 412146 338048
rect 419166 338036 419172 338048
rect 419224 338036 419230 338088
rect 420270 338036 420276 338088
rect 420328 338076 420334 338088
rect 445478 338076 445484 338088
rect 420328 338048 445484 338076
rect 420328 338036 420334 338048
rect 445478 338036 445484 338048
rect 445536 338036 445542 338088
rect 512270 338036 512276 338088
rect 512328 338076 512334 338088
rect 547138 338076 547144 338088
rect 512328 338048 547144 338076
rect 512328 338036 512334 338048
rect 547138 338036 547144 338048
rect 547196 338036 547202 338088
rect 66898 337968 66904 338020
rect 66956 338008 66962 338020
rect 261202 338008 261208 338020
rect 66956 337980 261208 338008
rect 66956 337968 66962 337980
rect 261202 337968 261208 337980
rect 261260 337968 261266 338020
rect 322750 337968 322756 338020
rect 322808 338008 322814 338020
rect 395246 338008 395252 338020
rect 322808 337980 395252 338008
rect 322808 337968 322814 337980
rect 395246 337968 395252 337980
rect 395304 337968 395310 338020
rect 395341 338011 395399 338017
rect 395341 337977 395353 338011
rect 395387 338008 395399 338011
rect 402606 338008 402612 338020
rect 395387 337980 402612 338008
rect 395387 337977 395399 337980
rect 395341 337971 395399 337977
rect 402606 337968 402612 337980
rect 402664 337968 402670 338020
rect 416682 337968 416688 338020
rect 416740 338008 416746 338020
rect 443638 338008 443644 338020
rect 416740 337980 443644 338008
rect 416740 337968 416746 337980
rect 443638 337968 443644 337980
rect 443696 337968 443702 338020
rect 451918 337968 451924 338020
rect 451976 338008 451982 338020
rect 459002 338008 459008 338020
rect 451976 337980 459008 338008
rect 451976 337968 451982 337980
rect 459002 337968 459008 337980
rect 459060 337968 459066 338020
rect 490834 337968 490840 338020
rect 490892 338008 490898 338020
rect 499025 338011 499083 338017
rect 499025 338008 499037 338011
rect 490892 337980 499037 338008
rect 490892 337968 490898 337980
rect 499025 337977 499037 337980
rect 499071 337977 499083 338011
rect 499025 337971 499083 337977
rect 512822 337968 512828 338020
rect 512880 338008 512886 338020
rect 547230 338008 547236 338020
rect 512880 337980 547236 338008
rect 512880 337968 512886 337980
rect 547230 337968 547236 337980
rect 547288 337968 547294 338020
rect 57238 337900 57244 337952
rect 57296 337940 57302 337952
rect 257522 337940 257528 337952
rect 57296 337912 257528 337940
rect 57296 337900 57302 337912
rect 257522 337900 257528 337912
rect 257580 337900 257586 337952
rect 309778 337900 309784 337952
rect 309836 337940 309842 337952
rect 309836 337912 315528 337940
rect 309836 337900 309842 337912
rect 50338 337832 50344 337884
rect 50396 337872 50402 337884
rect 251358 337872 251364 337884
rect 50396 337844 251364 337872
rect 50396 337832 50402 337844
rect 251358 337832 251364 337844
rect 251416 337832 251422 337884
rect 268378 337832 268384 337884
rect 268436 337872 268442 337884
rect 288710 337872 288716 337884
rect 268436 337844 288716 337872
rect 268436 337832 268442 337844
rect 288710 337832 288716 337844
rect 288768 337832 288774 337884
rect 311894 337832 311900 337884
rect 311952 337872 311958 337884
rect 312262 337872 312268 337884
rect 311952 337844 312268 337872
rect 311952 337832 311958 337844
rect 312262 337832 312268 337844
rect 312320 337832 312326 337884
rect 313458 337832 313464 337884
rect 313516 337872 313522 337884
rect 314102 337872 314108 337884
rect 313516 337844 314108 337872
rect 313516 337832 313522 337844
rect 314102 337832 314108 337844
rect 314160 337832 314166 337884
rect 314654 337832 314660 337884
rect 314712 337872 314718 337884
rect 315390 337872 315396 337884
rect 314712 337844 315396 337872
rect 314712 337832 314718 337844
rect 315390 337832 315396 337844
rect 315448 337832 315454 337884
rect 315500 337872 315528 337912
rect 316034 337900 316040 337952
rect 316092 337940 316098 337952
rect 316678 337940 316684 337952
rect 316092 337912 316684 337940
rect 316092 337900 316098 337912
rect 316678 337900 316684 337912
rect 316736 337900 316742 337952
rect 317598 337900 317604 337952
rect 317656 337940 317662 337952
rect 318334 337940 318340 337952
rect 317656 337912 318340 337940
rect 317656 337900 317662 337912
rect 318334 337900 318340 337912
rect 318392 337900 318398 337952
rect 320174 337900 320180 337952
rect 320232 337940 320238 337952
rect 320910 337940 320916 337952
rect 320232 337912 320916 337940
rect 320232 337900 320238 337912
rect 320910 337900 320916 337912
rect 320968 337900 320974 337952
rect 326341 337943 326399 337949
rect 326341 337909 326353 337943
rect 326387 337940 326399 337943
rect 384301 337943 384359 337949
rect 384301 337940 384313 337943
rect 326387 337912 384313 337940
rect 326387 337909 326399 337912
rect 326341 337903 326399 337909
rect 384301 337909 384313 337912
rect 384347 337909 384359 337943
rect 384301 337903 384359 337909
rect 385678 337900 385684 337952
rect 385736 337940 385742 337952
rect 389726 337940 389732 337952
rect 385736 337912 389732 337940
rect 385736 337900 385742 337912
rect 389726 337900 389732 337912
rect 389784 337900 389790 337952
rect 398745 337943 398803 337949
rect 398745 337940 398757 337943
rect 389836 337912 398757 337940
rect 387978 337872 387984 337884
rect 315500 337844 387984 337872
rect 387978 337832 387984 337844
rect 388036 337832 388042 337884
rect 388993 337875 389051 337881
rect 388993 337841 389005 337875
rect 389039 337872 389051 337875
rect 389836 337872 389864 337912
rect 398745 337909 398757 337912
rect 398791 337909 398803 337943
rect 398745 337903 398803 337909
rect 407758 337900 407764 337952
rect 407816 337940 407822 337952
rect 415486 337940 415492 337952
rect 407816 337912 415492 337940
rect 407816 337900 407822 337912
rect 415486 337900 415492 337912
rect 415544 337900 415550 337952
rect 420362 337940 420368 337952
rect 415596 337912 420368 337940
rect 389039 337844 389864 337872
rect 389039 337841 389051 337844
rect 388993 337835 389051 337841
rect 391198 337832 391204 337884
rect 391256 337872 391262 337884
rect 397086 337872 397092 337884
rect 391256 337844 397092 337872
rect 391256 337832 391262 337844
rect 397086 337832 397092 337844
rect 397144 337832 397150 337884
rect 398837 337875 398895 337881
rect 398837 337841 398849 337875
rect 398883 337872 398895 337875
rect 403989 337875 404047 337881
rect 403989 337872 404001 337875
rect 398883 337844 404001 337872
rect 398883 337841 398895 337844
rect 398837 337835 398895 337841
rect 403989 337841 404001 337844
rect 404035 337841 404047 337875
rect 403989 337835 404047 337841
rect 404998 337832 405004 337884
rect 405056 337872 405062 337884
rect 411806 337872 411812 337884
rect 405056 337844 411812 337872
rect 405056 337832 405062 337844
rect 411806 337832 411812 337844
rect 411864 337832 411870 337884
rect 413278 337832 413284 337884
rect 413336 337872 413342 337884
rect 415596 337872 415624 337912
rect 420362 337900 420368 337912
rect 420420 337900 420426 337952
rect 422941 337943 422999 337949
rect 422941 337909 422953 337943
rect 422987 337940 422999 337943
rect 432509 337943 432567 337949
rect 432509 337940 432521 337943
rect 422987 337912 432521 337940
rect 422987 337909 422999 337912
rect 422941 337903 422999 337909
rect 432509 337909 432521 337912
rect 432555 337909 432567 337943
rect 432509 337903 432567 337909
rect 432601 337943 432659 337949
rect 432601 337909 432613 337943
rect 432647 337940 432659 337943
rect 439958 337940 439964 337952
rect 432647 337912 439964 337940
rect 432647 337909 432659 337912
rect 432601 337903 432659 337909
rect 439958 337900 439964 337912
rect 440016 337900 440022 337952
rect 442258 337900 442264 337952
rect 442316 337940 442322 337952
rect 449802 337940 449808 337952
rect 442316 337912 449808 337940
rect 442316 337900 442322 337912
rect 449802 337900 449808 337912
rect 449860 337900 449866 337952
rect 453390 337900 453396 337952
rect 453448 337940 453454 337952
rect 462038 337940 462044 337952
rect 453448 337912 462044 337940
rect 453448 337900 453454 337912
rect 462038 337900 462044 337912
rect 462096 337900 462102 337952
rect 490190 337900 490196 337952
rect 490248 337940 490254 337952
rect 501598 337940 501604 337952
rect 490248 337912 501604 337940
rect 490248 337900 490254 337912
rect 501598 337900 501604 337912
rect 501656 337900 501662 337952
rect 503438 337900 503444 337952
rect 503496 337940 503502 337952
rect 503622 337940 503628 337952
rect 503496 337912 503628 337940
rect 503496 337900 503502 337912
rect 503622 337900 503628 337912
rect 503680 337900 503686 337952
rect 520826 337900 520832 337952
rect 520884 337940 520890 337952
rect 556798 337940 556804 337952
rect 520884 337912 556804 337940
rect 520884 337900 520890 337912
rect 556798 337900 556804 337912
rect 556856 337900 556862 337952
rect 413336 337844 415624 337872
rect 413336 337832 413342 337844
rect 416130 337832 416136 337884
rect 416188 337872 416194 337884
rect 442994 337872 443000 337884
rect 416188 337844 443000 337872
rect 416188 337832 416194 337844
rect 442994 337832 443000 337844
rect 443052 337832 443058 337884
rect 449250 337832 449256 337884
rect 449308 337872 449314 337884
rect 457162 337872 457168 337884
rect 449308 337844 457168 337872
rect 449308 337832 449314 337844
rect 457162 337832 457168 337844
rect 457220 337832 457226 337884
rect 497550 337832 497556 337884
rect 497608 337872 497614 337884
rect 509878 337872 509884 337884
rect 497608 337844 509884 337872
rect 497608 337832 497614 337844
rect 509878 337832 509884 337844
rect 509936 337832 509942 337884
rect 514662 337832 514668 337884
rect 514720 337872 514726 337884
rect 553394 337872 553400 337884
rect 514720 337844 553400 337872
rect 514720 337832 514726 337844
rect 553394 337832 553400 337844
rect 553452 337832 553458 337884
rect 46198 337764 46204 337816
rect 46256 337804 46262 337816
rect 247678 337804 247684 337816
rect 46256 337776 247684 337804
rect 46256 337764 46262 337776
rect 247678 337764 247684 337776
rect 247736 337764 247742 337816
rect 269758 337764 269764 337816
rect 269816 337804 269822 337816
rect 292390 337804 292396 337816
rect 269816 337776 292396 337804
rect 269816 337764 269822 337776
rect 292390 337764 292396 337776
rect 292448 337764 292454 337816
rect 294598 337764 294604 337816
rect 294656 337804 294662 337816
rect 375098 337804 375104 337816
rect 294656 337776 375104 337804
rect 294656 337764 294662 337776
rect 375098 337764 375104 337776
rect 375156 337764 375162 337816
rect 376018 337764 376024 337816
rect 376076 337804 376082 337816
rect 406286 337804 406292 337816
rect 376076 337776 406292 337804
rect 376076 337764 376082 337776
rect 406286 337764 406292 337776
rect 406344 337764 406350 337816
rect 409782 337764 409788 337816
rect 409840 337804 409846 337816
rect 432601 337807 432659 337813
rect 432601 337804 432613 337807
rect 409840 337776 432613 337804
rect 409840 337764 409846 337776
rect 432601 337773 432613 337776
rect 432647 337773 432659 337807
rect 432601 337767 432659 337773
rect 432693 337807 432751 337813
rect 432693 337773 432705 337807
rect 432739 337804 432751 337807
rect 436922 337804 436928 337816
rect 432739 337776 436928 337804
rect 432739 337773 432751 337776
rect 432693 337767 432751 337773
rect 436922 337764 436928 337776
rect 436980 337764 436986 337816
rect 437474 337764 437480 337816
rect 437532 337804 437538 337816
rect 438762 337804 438768 337816
rect 437532 337776 438768 337804
rect 437532 337764 437538 337776
rect 438762 337764 438768 337776
rect 438820 337764 438826 337816
rect 445018 337764 445024 337816
rect 445076 337804 445082 337816
rect 456518 337804 456524 337816
rect 445076 337776 456524 337804
rect 445076 337764 445082 337776
rect 456518 337764 456524 337776
rect 456576 337764 456582 337816
rect 463602 337764 463608 337816
rect 463660 337804 463666 337816
rect 468110 337804 468116 337816
rect 463660 337776 468116 337804
rect 463660 337764 463666 337776
rect 468110 337764 468116 337776
rect 468168 337764 468174 337816
rect 488994 337764 489000 337816
rect 489052 337804 489058 337816
rect 502610 337804 502616 337816
rect 489052 337776 502616 337804
rect 489052 337764 489058 337776
rect 502610 337764 502616 337776
rect 502668 337764 502674 337816
rect 504266 337764 504272 337816
rect 504324 337804 504330 337816
rect 505002 337804 505008 337816
rect 504324 337776 505008 337804
rect 504324 337764 504330 337776
rect 505002 337764 505008 337776
rect 505060 337764 505066 337816
rect 505388 337776 506520 337804
rect 39298 337696 39304 337748
rect 39356 337736 39362 337748
rect 234617 337739 234675 337745
rect 234617 337736 234629 337739
rect 39356 337708 234629 337736
rect 39356 337696 39362 337708
rect 234617 337705 234629 337708
rect 234663 337705 234675 337739
rect 234617 337699 234675 337705
rect 236825 337739 236883 337745
rect 236825 337705 236837 337739
rect 236871 337736 236883 337739
rect 240410 337736 240416 337748
rect 236871 337708 240416 337736
rect 236871 337705 236883 337708
rect 236825 337699 236883 337705
rect 240410 337696 240416 337708
rect 240468 337696 240474 337748
rect 258718 337696 258724 337748
rect 258776 337736 258782 337748
rect 266722 337736 266728 337748
rect 258776 337708 266728 337736
rect 258776 337696 258782 337708
rect 266722 337696 266728 337708
rect 266780 337696 266786 337748
rect 287698 337696 287704 337748
rect 287756 337736 287762 337748
rect 369578 337736 369584 337748
rect 287756 337708 369584 337736
rect 287756 337696 287762 337708
rect 369578 337696 369584 337708
rect 369636 337696 369642 337748
rect 374638 337696 374644 337748
rect 374696 337736 374702 337748
rect 409966 337736 409972 337748
rect 374696 337708 409972 337736
rect 374696 337696 374702 337708
rect 409966 337696 409972 337708
rect 410024 337696 410030 337748
rect 412542 337696 412548 337748
rect 412600 337736 412606 337748
rect 441798 337736 441804 337748
rect 412600 337708 441804 337736
rect 412600 337696 412606 337708
rect 441798 337696 441804 337708
rect 441856 337696 441862 337748
rect 442350 337696 442356 337748
rect 442408 337736 442414 337748
rect 454678 337736 454684 337748
rect 442408 337708 454684 337736
rect 442408 337696 442414 337708
rect 454678 337696 454684 337708
rect 454736 337696 454742 337748
rect 487154 337696 487160 337748
rect 487212 337736 487218 337748
rect 499758 337736 499764 337748
rect 487212 337708 499764 337736
rect 487212 337696 487218 337708
rect 499758 337696 499764 337708
rect 499816 337696 499822 337748
rect 499942 337696 499948 337748
rect 500000 337736 500006 337748
rect 500862 337736 500868 337748
rect 500000 337708 500868 337736
rect 500000 337696 500006 337708
rect 500862 337696 500868 337708
rect 500920 337696 500926 337748
rect 501230 337696 501236 337748
rect 501288 337736 501294 337748
rect 505388 337736 505416 337776
rect 501288 337708 505416 337736
rect 501288 337696 501294 337708
rect 505462 337696 505468 337748
rect 505520 337736 505526 337748
rect 506382 337736 506388 337748
rect 505520 337708 506388 337736
rect 505520 337696 505526 337708
rect 506382 337696 506388 337708
rect 506440 337696 506446 337748
rect 506492 337736 506520 337776
rect 507946 337764 507952 337816
rect 508004 337804 508010 337816
rect 509142 337804 509148 337816
rect 508004 337776 509148 337804
rect 508004 337764 508010 337776
rect 509142 337764 509148 337776
rect 509200 337764 509206 337816
rect 515858 337764 515864 337816
rect 515916 337804 515922 337816
rect 554866 337804 554872 337816
rect 515916 337776 554872 337804
rect 515916 337764 515922 337776
rect 554866 337764 554872 337776
rect 554924 337764 554930 337816
rect 506492 337708 513052 337736
rect 32398 337628 32404 337680
rect 32456 337668 32462 337680
rect 239401 337671 239459 337677
rect 239401 337668 239413 337671
rect 32456 337640 239413 337668
rect 32456 337628 32462 337640
rect 239401 337637 239413 337640
rect 239447 337637 239459 337671
rect 239401 337631 239459 337637
rect 253382 337628 253388 337680
rect 253440 337668 253446 337680
rect 255682 337668 255688 337680
rect 253440 337640 255688 337668
rect 253440 337628 253446 337640
rect 255682 337628 255688 337640
rect 255740 337628 255746 337680
rect 264330 337628 264336 337680
rect 264388 337668 264394 337680
rect 281442 337668 281448 337680
rect 264388 337640 281448 337668
rect 264388 337628 264394 337640
rect 281442 337628 281448 337640
rect 281500 337628 281506 337680
rect 283558 337628 283564 337680
rect 283616 337668 283622 337680
rect 365898 337668 365904 337680
rect 283616 337640 365904 337668
rect 283616 337628 283622 337640
rect 365898 337628 365904 337640
rect 365956 337628 365962 337680
rect 366910 337628 366916 337680
rect 366968 337668 366974 337680
rect 418522 337668 418528 337680
rect 366968 337640 418528 337668
rect 366968 337628 366974 337640
rect 418522 337628 418528 337640
rect 418580 337628 418586 337680
rect 420822 337628 420828 337680
rect 420880 337668 420886 337680
rect 446122 337668 446128 337680
rect 420880 337640 446128 337668
rect 420880 337628 420886 337640
rect 446122 337628 446128 337640
rect 446180 337628 446186 337680
rect 456058 337628 456064 337680
rect 456116 337668 456122 337680
rect 463878 337668 463884 337680
rect 456116 337640 463884 337668
rect 456116 337628 456122 337640
rect 463878 337628 463884 337640
rect 463936 337628 463942 337680
rect 466362 337628 466368 337680
rect 466420 337668 466426 337680
rect 469398 337668 469404 337680
rect 466420 337640 469404 337668
rect 466420 337628 466426 337640
rect 469398 337628 469404 337640
rect 469456 337628 469462 337680
rect 475470 337628 475476 337680
rect 475528 337668 475534 337680
rect 477678 337668 477684 337680
rect 475528 337640 477684 337668
rect 475528 337628 475534 337640
rect 477678 337628 477684 337640
rect 477736 337628 477742 337680
rect 485866 337628 485872 337680
rect 485924 337668 485930 337680
rect 489178 337668 489184 337680
rect 485924 337640 489184 337668
rect 485924 337628 485930 337640
rect 489178 337628 489184 337640
rect 489236 337628 489242 337680
rect 491386 337628 491392 337680
rect 491444 337668 491450 337680
rect 492490 337668 492496 337680
rect 491444 337640 492496 337668
rect 491444 337628 491450 337640
rect 492490 337628 492496 337640
rect 492548 337628 492554 337680
rect 495066 337628 495072 337680
rect 495124 337668 495130 337680
rect 496078 337668 496084 337680
rect 495124 337640 496084 337668
rect 495124 337628 495130 337640
rect 496078 337628 496084 337640
rect 496136 337628 496142 337680
rect 496906 337628 496912 337680
rect 496964 337668 496970 337680
rect 498838 337668 498844 337680
rect 496964 337640 498844 337668
rect 496964 337628 496970 337640
rect 498838 337628 498844 337640
rect 498896 337628 498902 337680
rect 510798 337668 510804 337680
rect 498948 337640 510804 337668
rect 28258 337560 28264 337612
rect 28316 337600 28322 337612
rect 236825 337603 236883 337609
rect 236825 337600 236837 337603
rect 28316 337572 236837 337600
rect 28316 337560 28322 337572
rect 236825 337569 236837 337572
rect 236871 337569 236883 337603
rect 248322 337600 248328 337612
rect 236825 337563 236883 337569
rect 237576 337572 248328 337600
rect 3326 337492 3332 337544
rect 3384 337532 3390 337544
rect 7834 337532 7840 337544
rect 3384 337504 7840 337532
rect 3384 337492 3390 337504
rect 7834 337492 7840 337504
rect 7892 337492 7898 337544
rect 17218 337492 17224 337544
rect 17276 337532 17282 337544
rect 228085 337535 228143 337541
rect 228085 337532 228097 337535
rect 17276 337504 228097 337532
rect 17276 337492 17282 337504
rect 228085 337501 228097 337504
rect 228131 337501 228143 337535
rect 228085 337495 228143 337501
rect 228174 337492 228180 337544
rect 228232 337532 228238 337544
rect 234890 337532 234896 337544
rect 228232 337504 234896 337532
rect 228232 337492 228238 337504
rect 234890 337492 234896 337504
rect 234948 337492 234954 337544
rect 234985 337535 235043 337541
rect 234985 337501 234997 337535
rect 235031 337532 235043 337535
rect 237576 337532 237604 337572
rect 248322 337560 248328 337572
rect 248380 337560 248386 337612
rect 289998 337600 290004 337612
rect 248432 337572 290004 337600
rect 235031 337504 237604 337532
rect 239401 337535 239459 337541
rect 235031 337501 235043 337504
rect 234985 337495 235043 337501
rect 239401 337501 239413 337535
rect 239447 337532 239459 337535
rect 244642 337532 244648 337544
rect 239447 337504 244648 337532
rect 239447 337501 239459 337504
rect 239401 337495 239459 337501
rect 244642 337492 244648 337504
rect 244700 337492 244706 337544
rect 246298 337492 246304 337544
rect 246356 337532 246362 337544
rect 248432 337532 248460 337572
rect 289998 337560 290004 337572
rect 290056 337560 290062 337612
rect 293862 337560 293868 337612
rect 293920 337600 293926 337612
rect 380618 337600 380624 337612
rect 293920 337572 380624 337600
rect 293920 337560 293926 337572
rect 380618 337560 380624 337572
rect 380676 337560 380682 337612
rect 384301 337603 384359 337609
rect 384301 337569 384313 337603
rect 384347 337600 384359 337603
rect 391566 337600 391572 337612
rect 384347 337572 391572 337600
rect 384347 337569 384359 337572
rect 384301 337563 384359 337569
rect 391566 337560 391572 337572
rect 391624 337560 391630 337612
rect 393222 337560 393228 337612
rect 393280 337600 393286 337612
rect 432046 337600 432052 337612
rect 393280 337572 432052 337600
rect 393280 337560 393286 337572
rect 432046 337560 432052 337572
rect 432104 337560 432110 337612
rect 432509 337603 432567 337609
rect 432509 337569 432521 337603
rect 432555 337600 432567 337603
rect 441246 337600 441252 337612
rect 432555 337572 441252 337600
rect 432555 337569 432567 337572
rect 432509 337563 432567 337569
rect 441246 337560 441252 337572
rect 441304 337560 441310 337612
rect 441341 337603 441399 337609
rect 441341 337569 441353 337603
rect 441387 337600 441399 337603
rect 452838 337600 452844 337612
rect 441387 337572 452844 337600
rect 441387 337569 441399 337572
rect 441341 337563 441399 337569
rect 452838 337560 452844 337572
rect 452896 337560 452902 337612
rect 453942 337560 453948 337612
rect 454000 337600 454006 337612
rect 463234 337600 463240 337612
rect 454000 337572 463240 337600
rect 454000 337560 454006 337572
rect 463234 337560 463240 337572
rect 463292 337560 463298 337612
rect 492674 337560 492680 337612
rect 492732 337600 492738 337612
rect 498948 337600 498976 337640
rect 510798 337628 510804 337640
rect 510856 337628 510862 337680
rect 513024 337668 513052 337708
rect 518342 337696 518348 337748
rect 518400 337736 518406 337748
rect 560294 337736 560300 337748
rect 518400 337708 560300 337736
rect 518400 337696 518406 337708
rect 560294 337696 560300 337708
rect 560352 337696 560358 337748
rect 516778 337668 516784 337680
rect 513024 337640 516784 337668
rect 516778 337628 516784 337640
rect 516836 337628 516842 337680
rect 526809 337671 526867 337677
rect 526809 337668 526821 337671
rect 519556 337640 526821 337668
rect 492732 337572 498976 337600
rect 499025 337603 499083 337609
rect 492732 337560 492738 337572
rect 499025 337569 499037 337603
rect 499071 337600 499083 337603
rect 502337 337603 502395 337609
rect 502337 337600 502349 337603
rect 499071 337572 502349 337600
rect 499071 337569 499083 337572
rect 499025 337563 499083 337569
rect 502337 337569 502349 337572
rect 502383 337569 502395 337603
rect 502337 337563 502395 337569
rect 502426 337560 502432 337612
rect 502484 337600 502490 337612
rect 503530 337600 503536 337612
rect 502484 337572 503536 337600
rect 502484 337560 502490 337572
rect 503530 337560 503536 337572
rect 503588 337560 503594 337612
rect 508590 337560 508596 337612
rect 508648 337600 508654 337612
rect 519556 337600 519584 337640
rect 526809 337637 526821 337640
rect 526855 337637 526867 337671
rect 526809 337631 526867 337637
rect 526898 337628 526904 337680
rect 526956 337668 526962 337680
rect 529017 337671 529075 337677
rect 529017 337668 529029 337671
rect 526956 337640 529029 337668
rect 526956 337628 526962 337640
rect 529017 337637 529029 337640
rect 529063 337637 529075 337671
rect 563146 337668 563152 337680
rect 529017 337631 529075 337637
rect 529216 337640 563152 337668
rect 508648 337572 519584 337600
rect 508648 337560 508654 337572
rect 246356 337504 248460 337532
rect 246356 337492 246362 337504
rect 262858 337492 262864 337544
rect 262916 337532 262922 337544
rect 267461 337535 267519 337541
rect 267461 337532 267473 337535
rect 262916 337504 267473 337532
rect 262916 337492 262922 337504
rect 267461 337501 267473 337504
rect 267507 337501 267519 337535
rect 267461 337495 267519 337501
rect 267553 337535 267611 337541
rect 267553 337501 267565 337535
rect 267599 337532 267611 337535
rect 285030 337532 285036 337544
rect 267599 337504 285036 337532
rect 267599 337501 267611 337504
rect 267553 337495 267611 337501
rect 285030 337492 285036 337504
rect 285088 337492 285094 337544
rect 286962 337492 286968 337544
rect 287020 337532 287026 337544
rect 376938 337532 376944 337544
rect 287020 337504 376944 337532
rect 287020 337492 287026 337504
rect 376938 337492 376944 337504
rect 376996 337492 377002 337544
rect 377033 337535 377091 337541
rect 377033 337501 377045 337535
rect 377079 337532 377091 337535
rect 384022 337532 384028 337544
rect 377079 337504 384028 337532
rect 377079 337501 377091 337504
rect 377033 337495 377091 337501
rect 384022 337492 384028 337504
rect 384080 337492 384086 337544
rect 386417 337535 386475 337541
rect 386417 337501 386429 337535
rect 386463 337532 386475 337535
rect 388993 337535 389051 337541
rect 388993 337532 389005 337535
rect 386463 337504 389005 337532
rect 386463 337501 386475 337504
rect 386417 337495 386475 337501
rect 388993 337501 389005 337504
rect 389039 337501 389051 337535
rect 388993 337495 389051 337501
rect 389082 337492 389088 337544
rect 389140 337532 389146 337544
rect 389140 337504 422984 337532
rect 389140 337492 389146 337504
rect 24118 337424 24124 337476
rect 24176 337464 24182 337476
rect 24176 337436 237236 337464
rect 24176 337424 24182 337436
rect 15838 337356 15844 337408
rect 15896 337396 15902 337408
rect 228174 337396 228180 337408
rect 15896 337368 228180 337396
rect 15896 337356 15902 337368
rect 228174 337356 228180 337368
rect 228232 337356 228238 337408
rect 228269 337399 228327 337405
rect 228269 337365 228281 337399
rect 228315 337396 228327 337399
rect 235442 337396 235448 337408
rect 228315 337368 235448 337396
rect 228315 337365 228327 337368
rect 228269 337359 228327 337365
rect 235442 337356 235448 337368
rect 235500 337356 235506 337408
rect 237208 337396 237236 337436
rect 261478 337424 261484 337476
rect 261536 337464 261542 337476
rect 261536 337436 264192 337464
rect 261536 337424 261542 337436
rect 239766 337396 239772 337408
rect 237208 337368 239772 337396
rect 239766 337356 239772 337368
rect 239824 337356 239830 337408
rect 257338 337356 257344 337408
rect 257396 337396 257402 337408
rect 263042 337396 263048 337408
rect 257396 337368 263048 337396
rect 257396 337356 257402 337368
rect 263042 337356 263048 337368
rect 263100 337356 263106 337408
rect 61378 337288 61384 337340
rect 61436 337328 61442 337340
rect 251726 337328 251732 337340
rect 61436 337300 251732 337328
rect 61436 337288 61442 337300
rect 251726 337288 251732 337300
rect 251784 337288 251790 337340
rect 251818 337288 251824 337340
rect 251876 337328 251882 337340
rect 253198 337328 253204 337340
rect 251876 337300 253204 337328
rect 251876 337288 251882 337300
rect 253198 337288 253204 337300
rect 253256 337288 253262 337340
rect 255958 337288 255964 337340
rect 256016 337328 256022 337340
rect 259362 337328 259368 337340
rect 256016 337300 259368 337328
rect 256016 337288 256022 337300
rect 259362 337288 259368 337300
rect 259420 337288 259426 337340
rect 264164 337328 264192 337436
rect 264238 337424 264244 337476
rect 264296 337464 264302 337476
rect 279602 337464 279608 337476
rect 264296 337436 279608 337464
rect 264296 337424 264302 337436
rect 279602 337424 279608 337436
rect 279660 337424 279666 337476
rect 280062 337424 280068 337476
rect 280120 337464 280126 337476
rect 373258 337464 373264 337476
rect 280120 337436 373264 337464
rect 280120 337424 280126 337436
rect 373258 337424 373264 337436
rect 373316 337424 373322 337476
rect 375282 337424 375288 337476
rect 375340 337464 375346 337476
rect 422202 337464 422208 337476
rect 375340 337436 422208 337464
rect 375340 337424 375346 337436
rect 422202 337424 422208 337436
rect 422260 337424 422266 337476
rect 267461 337399 267519 337405
rect 267461 337365 267473 337399
rect 267507 337396 267519 337399
rect 275922 337396 275928 337408
rect 267507 337368 275928 337396
rect 267507 337365 267519 337368
rect 267461 337359 267519 337365
rect 275922 337356 275928 337368
rect 275980 337356 275986 337408
rect 276658 337356 276664 337408
rect 276716 337396 276722 337408
rect 371418 337396 371424 337408
rect 276716 337368 371424 337396
rect 276716 337356 276722 337368
rect 371418 337356 371424 337368
rect 371476 337356 371482 337408
rect 372522 337356 372528 337408
rect 372580 337396 372586 337408
rect 421006 337396 421012 337408
rect 372580 337368 421012 337396
rect 372580 337356 372586 337368
rect 421006 337356 421012 337368
rect 421064 337356 421070 337408
rect 422956 337396 422984 337504
rect 432598 337492 432604 337544
rect 432656 337532 432662 337544
rect 435726 337532 435732 337544
rect 432656 337504 435732 337532
rect 432656 337492 432662 337504
rect 435726 337492 435732 337504
rect 435784 337492 435790 337544
rect 435821 337535 435879 337541
rect 435821 337501 435833 337535
rect 435867 337532 435879 337535
rect 450998 337532 451004 337544
rect 435867 337504 451004 337532
rect 435867 337501 435879 337504
rect 435821 337495 435879 337501
rect 450998 337492 451004 337504
rect 451056 337492 451062 337544
rect 451182 337492 451188 337544
rect 451240 337532 451246 337544
rect 461394 337532 461400 337544
rect 451240 337504 461400 337532
rect 451240 337492 451246 337504
rect 461394 337492 461400 337504
rect 461452 337492 461458 337544
rect 479794 337492 479800 337544
rect 479852 337532 479858 337544
rect 485958 337532 485964 337544
rect 479852 337504 485964 337532
rect 479852 337492 479858 337504
rect 485958 337492 485964 337504
rect 486016 337492 486022 337544
rect 494514 337492 494520 337544
rect 494572 337532 494578 337544
rect 513558 337532 513564 337544
rect 494572 337504 513564 337532
rect 494572 337492 494578 337504
rect 513558 337492 513564 337504
rect 513616 337492 513622 337544
rect 526809 337535 526867 337541
rect 526809 337501 526821 337535
rect 526855 337532 526867 337535
rect 528922 337532 528928 337544
rect 526855 337504 528928 337532
rect 526855 337501 526867 337504
rect 526809 337495 526867 337501
rect 528922 337492 528928 337504
rect 528980 337492 528986 337544
rect 529216 337532 529244 337640
rect 563146 337628 563152 337640
rect 563204 337628 563210 337680
rect 529382 337560 529388 337612
rect 529440 337600 529446 337612
rect 573358 337600 573364 337612
rect 529440 337572 573364 337600
rect 529440 337560 529446 337572
rect 573358 337560 573364 337572
rect 573416 337560 573422 337612
rect 529032 337504 529244 337532
rect 529293 337535 529351 337541
rect 423033 337467 423091 337473
rect 423033 337433 423045 337467
rect 423079 337464 423091 337467
rect 446398 337464 446404 337476
rect 423079 337436 446404 337464
rect 423079 337433 423091 337436
rect 423033 337427 423091 337433
rect 446398 337424 446404 337436
rect 446456 337424 446462 337476
rect 446490 337424 446496 337476
rect 446548 337464 446554 337476
rect 458358 337464 458364 337476
rect 446548 337436 458364 337464
rect 446548 337424 446554 337436
rect 458358 337424 458364 337436
rect 458416 337424 458422 337476
rect 485314 337424 485320 337476
rect 485372 337464 485378 337476
rect 493318 337464 493324 337476
rect 485372 337436 493324 337464
rect 485372 337424 485378 337436
rect 493318 337424 493324 337436
rect 493376 337424 493382 337476
rect 496262 337424 496268 337476
rect 496320 337464 496326 337476
rect 496320 337436 510936 337464
rect 496320 337424 496326 337436
rect 429562 337396 429568 337408
rect 422956 337368 429568 337396
rect 429562 337356 429568 337368
rect 429620 337356 429626 337408
rect 431129 337399 431187 337405
rect 431129 337365 431141 337399
rect 431175 337396 431187 337399
rect 432509 337399 432567 337405
rect 432509 337396 432521 337399
rect 431175 337368 432521 337396
rect 431175 337365 431187 337368
rect 431129 337359 431187 337365
rect 432509 337365 432521 337368
rect 432555 337365 432567 337399
rect 432509 337359 432567 337365
rect 432601 337399 432659 337405
rect 432601 337365 432613 337399
rect 432647 337396 432659 337399
rect 447318 337396 447324 337408
rect 432647 337368 447324 337396
rect 432647 337365 432659 337368
rect 432601 337359 432659 337365
rect 447318 337356 447324 337368
rect 447376 337356 447382 337408
rect 453298 337356 453304 337408
rect 453356 337396 453362 337408
rect 460750 337396 460756 337408
rect 453356 337368 460756 337396
rect 453356 337356 453362 337368
rect 460750 337356 460756 337368
rect 460808 337356 460814 337408
rect 460842 337356 460848 337408
rect 460900 337396 460906 337408
rect 466914 337396 466920 337408
rect 460900 337368 466920 337396
rect 460900 337356 460906 337368
rect 466914 337356 466920 337368
rect 466972 337356 466978 337408
rect 482830 337356 482836 337408
rect 482888 337396 482894 337408
rect 491478 337396 491484 337408
rect 482888 337368 491484 337396
rect 482888 337356 482894 337368
rect 491478 337356 491484 337368
rect 491536 337356 491542 337408
rect 510908 337396 510936 337436
rect 510982 337424 510988 337476
rect 511040 337464 511046 337476
rect 511810 337464 511816 337476
rect 511040 337436 511816 337464
rect 511040 337424 511046 337436
rect 511810 337424 511816 337436
rect 511868 337424 511874 337476
rect 515306 337424 515312 337476
rect 515364 337464 515370 337476
rect 515364 337436 519492 337464
rect 515364 337424 515370 337436
rect 517606 337396 517612 337408
rect 510908 337368 517612 337396
rect 517606 337356 517612 337368
rect 517664 337356 517670 337408
rect 519464 337396 519492 337436
rect 519538 337424 519544 337476
rect 519596 337464 519602 337476
rect 529032 337464 529060 337504
rect 529293 337501 529305 337535
rect 529339 337532 529351 337535
rect 567194 337532 567200 337544
rect 529339 337504 567200 337532
rect 529339 337501 529351 337504
rect 529293 337495 529351 337501
rect 567194 337492 567200 337504
rect 567252 337492 567258 337544
rect 519596 337436 529060 337464
rect 519596 337424 519602 337436
rect 529474 337424 529480 337476
rect 529532 337464 529538 337476
rect 569218 337464 569224 337476
rect 529532 337436 569224 337464
rect 529532 337424 529538 337436
rect 569218 337424 569224 337436
rect 569276 337424 569282 337476
rect 520185 337399 520243 337405
rect 520185 337396 520197 337399
rect 519464 337368 520197 337396
rect 520185 337365 520197 337368
rect 520231 337365 520243 337399
rect 520185 337359 520243 337365
rect 524417 337399 524475 337405
rect 524417 337365 524429 337399
rect 524463 337396 524475 337399
rect 531314 337396 531320 337408
rect 524463 337368 531320 337396
rect 524463 337365 524475 337368
rect 524417 337359 524475 337365
rect 531314 337356 531320 337368
rect 531372 337356 531378 337408
rect 531409 337399 531467 337405
rect 531409 337365 531421 337399
rect 531455 337396 531467 337399
rect 571978 337396 571984 337408
rect 531455 337368 571984 337396
rect 531455 337365 531467 337368
rect 531409 337359 531467 337365
rect 571978 337356 571984 337368
rect 572036 337356 572042 337408
rect 270402 337328 270408 337340
rect 264164 337300 270408 337328
rect 270402 337288 270408 337300
rect 270460 337288 270466 337340
rect 284938 337288 284944 337340
rect 284996 337328 285002 337340
rect 338942 337328 338948 337340
rect 284996 337300 338948 337328
rect 284996 337288 285002 337300
rect 338942 337288 338948 337300
rect 339000 337288 339006 337340
rect 357345 337331 357403 337337
rect 357345 337297 357357 337331
rect 357391 337328 357403 337331
rect 367097 337331 367155 337337
rect 367097 337328 367109 337331
rect 357391 337300 367109 337328
rect 357391 337297 357403 337300
rect 357345 337291 357403 337297
rect 367097 337297 367109 337300
rect 367143 337297 367155 337331
rect 367097 337291 367155 337297
rect 379425 337331 379483 337337
rect 379425 337297 379437 337331
rect 379471 337328 379483 337331
rect 386417 337331 386475 337337
rect 386417 337328 386429 337331
rect 379471 337300 386429 337328
rect 379471 337297 379483 337300
rect 379425 337291 379483 337297
rect 386417 337297 386429 337300
rect 386463 337297 386475 337331
rect 386417 337291 386475 337297
rect 398745 337331 398803 337337
rect 398745 337297 398757 337331
rect 398791 337328 398803 337331
rect 403894 337328 403900 337340
rect 398791 337300 403900 337328
rect 398791 337297 398803 337300
rect 398745 337291 398803 337297
rect 403894 337288 403900 337300
rect 403952 337288 403958 337340
rect 403989 337331 404047 337337
rect 403989 337297 404001 337331
rect 404035 337328 404047 337331
rect 411162 337328 411168 337340
rect 404035 337300 411168 337328
rect 404035 337297 404047 337300
rect 403989 337291 404047 337297
rect 411162 337288 411168 337300
rect 411220 337288 411226 337340
rect 428366 337328 428372 337340
rect 411272 337300 428372 337328
rect 84838 337220 84844 337272
rect 84896 337260 84902 337272
rect 272242 337260 272248 337272
rect 84896 337232 272248 337260
rect 84896 337220 84902 337232
rect 272242 337220 272248 337232
rect 272300 337220 272306 337272
rect 283650 337220 283656 337272
rect 283708 337260 283714 337272
rect 337102 337260 337108 337272
rect 283708 337232 337108 337260
rect 283708 337220 283714 337232
rect 337102 337220 337108 337232
rect 337160 337220 337166 337272
rect 339402 337220 339408 337272
rect 339460 337260 339466 337272
rect 339460 337232 345704 337260
rect 339460 337220 339466 337232
rect 97258 337152 97264 337204
rect 97316 337192 97322 337204
rect 277762 337192 277768 337204
rect 97316 337164 277768 337192
rect 97316 337152 97322 337164
rect 277762 337152 277768 337164
rect 277820 337152 277826 337204
rect 316678 337152 316684 337204
rect 316736 337192 316742 337204
rect 326341 337195 326399 337201
rect 326341 337192 326353 337195
rect 316736 337164 326353 337192
rect 316736 337152 316742 337164
rect 326341 337161 326353 337164
rect 326387 337161 326399 337195
rect 345676 337192 345704 337232
rect 346302 337220 346308 337272
rect 346360 337260 346366 337272
rect 407482 337260 407488 337272
rect 346360 337232 407488 337260
rect 346360 337220 346366 337232
rect 407482 337220 407488 337232
rect 407540 337220 407546 337272
rect 409138 337220 409144 337272
rect 409196 337260 409202 337272
rect 411272 337260 411300 337300
rect 428366 337288 428372 337300
rect 428424 337288 428430 337340
rect 428550 337288 428556 337340
rect 428608 337328 428614 337340
rect 433337 337331 433395 337337
rect 433337 337328 433349 337331
rect 428608 337300 433349 337328
rect 428608 337288 428614 337300
rect 433337 337297 433349 337300
rect 433383 337297 433395 337331
rect 433337 337291 433395 337297
rect 433429 337331 433487 337337
rect 433429 337297 433441 337331
rect 433475 337328 433487 337331
rect 450354 337328 450360 337340
rect 433475 337300 450360 337328
rect 433475 337297 433487 337300
rect 433429 337291 433487 337297
rect 450354 337288 450360 337300
rect 450412 337288 450418 337340
rect 502337 337331 502395 337337
rect 502337 337297 502349 337331
rect 502383 337328 502395 337331
rect 506658 337328 506664 337340
rect 502383 337300 506664 337328
rect 502383 337297 502395 337300
rect 502337 337291 502395 337297
rect 506658 337288 506664 337300
rect 506716 337288 506722 337340
rect 520366 337328 520372 337340
rect 507872 337300 520372 337328
rect 409196 337232 411300 337260
rect 409196 337220 409202 337232
rect 413462 337220 413468 337272
rect 413520 337260 413526 337272
rect 413520 337232 421144 337260
rect 413520 337220 413526 337232
rect 347777 337195 347835 337201
rect 347777 337192 347789 337195
rect 345676 337164 347789 337192
rect 326341 337155 326399 337161
rect 347777 337161 347789 337164
rect 347823 337161 347835 337195
rect 398837 337195 398895 337201
rect 398837 337192 398849 337195
rect 347777 337155 347835 337161
rect 354600 337164 398849 337192
rect 104802 337084 104808 337136
rect 104860 337124 104866 337136
rect 283190 337124 283196 337136
rect 104860 337096 283196 337124
rect 104860 337084 104866 337096
rect 283190 337084 283196 337096
rect 283248 337084 283254 337136
rect 353202 337084 353208 337136
rect 353260 337124 353266 337136
rect 354600 337124 354628 337164
rect 398837 337161 398849 337164
rect 398883 337161 398895 337195
rect 398837 337155 398895 337161
rect 417602 337152 417608 337204
rect 417660 337192 417666 337204
rect 421009 337195 421067 337201
rect 421009 337192 421021 337195
rect 417660 337164 421021 337192
rect 417660 337152 417666 337164
rect 421009 337161 421021 337164
rect 421055 337161 421067 337195
rect 421116 337192 421144 337232
rect 422202 337220 422208 337272
rect 422260 337260 422266 337272
rect 423033 337263 423091 337269
rect 423033 337260 423045 337263
rect 422260 337232 423045 337260
rect 422260 337220 422266 337232
rect 423033 337229 423045 337232
rect 423079 337229 423091 337263
rect 423033 337223 423091 337229
rect 424962 337220 424968 337272
rect 425020 337260 425026 337272
rect 447962 337260 447968 337272
rect 425020 337232 447968 337260
rect 425020 337220 425026 337232
rect 447962 337220 447968 337232
rect 448020 337220 448026 337272
rect 448422 337220 448428 337272
rect 448480 337260 448486 337272
rect 460198 337260 460204 337272
rect 448480 337232 460204 337260
rect 448480 337220 448486 337232
rect 460198 337220 460204 337232
rect 460256 337220 460262 337272
rect 495710 337220 495716 337272
rect 495768 337260 495774 337272
rect 496722 337260 496728 337272
rect 495768 337232 496728 337260
rect 495768 337220 495774 337232
rect 496722 337220 496728 337232
rect 496780 337220 496786 337272
rect 506750 337220 506756 337272
rect 506808 337260 506814 337272
rect 507762 337260 507768 337272
rect 506808 337232 507768 337260
rect 506808 337220 506814 337232
rect 507762 337220 507768 337232
rect 507820 337220 507826 337272
rect 424042 337192 424048 337204
rect 421116 337164 424048 337192
rect 421009 337155 421067 337161
rect 424042 337152 424048 337164
rect 424100 337152 424106 337204
rect 430485 337195 430543 337201
rect 430485 337161 430497 337195
rect 430531 337192 430543 337195
rect 433242 337192 433248 337204
rect 430531 337164 433248 337192
rect 430531 337161 430543 337164
rect 430485 337155 430543 337161
rect 433242 337152 433248 337164
rect 433300 337152 433306 337204
rect 433337 337195 433395 337201
rect 433337 337161 433349 337195
rect 433383 337192 433395 337195
rect 449158 337192 449164 337204
rect 433383 337164 449164 337192
rect 433383 337161 433395 337164
rect 433337 337155 433395 337161
rect 449158 337152 449164 337164
rect 449216 337152 449222 337204
rect 498102 337152 498108 337204
rect 498160 337192 498166 337204
rect 507872 337192 507900 337300
rect 520366 337288 520372 337300
rect 520424 337288 520430 337340
rect 549898 337328 549904 337340
rect 520752 337300 549904 337328
rect 517146 337220 517152 337272
rect 517204 337260 517210 337272
rect 520752 337260 520780 337300
rect 549898 337288 549904 337300
rect 549956 337288 549962 337340
rect 517204 337232 520780 337260
rect 517204 337220 517210 337232
rect 522022 337220 522028 337272
rect 522080 337260 522086 337272
rect 529293 337263 529351 337269
rect 529293 337260 529305 337263
rect 522080 337232 529305 337260
rect 522080 337220 522086 337232
rect 529293 337229 529305 337232
rect 529339 337229 529351 337263
rect 529293 337223 529351 337229
rect 529385 337263 529443 337269
rect 529385 337229 529397 337263
rect 529431 337260 529443 337263
rect 531409 337263 531467 337269
rect 531409 337260 531421 337263
rect 529431 337232 531421 337260
rect 529431 337229 529443 337232
rect 529385 337223 529443 337229
rect 531409 337229 531421 337232
rect 531455 337229 531467 337263
rect 531409 337223 531467 337229
rect 531501 337263 531559 337269
rect 531501 337229 531513 337263
rect 531547 337260 531559 337263
rect 558178 337260 558184 337272
rect 531547 337232 558184 337260
rect 531547 337229 531559 337232
rect 531501 337223 531559 337229
rect 558178 337220 558184 337232
rect 558236 337220 558242 337272
rect 498160 337164 507900 337192
rect 498160 337152 498166 337164
rect 509050 337152 509056 337204
rect 509108 337192 509114 337204
rect 540238 337192 540244 337204
rect 509108 337164 540244 337192
rect 509108 337152 509114 337164
rect 540238 337152 540244 337164
rect 540296 337152 540302 337204
rect 353260 337096 354628 337124
rect 353260 337084 353266 337096
rect 357342 337084 357348 337136
rect 357400 337124 357406 337136
rect 413646 337124 413652 337136
rect 357400 337096 413652 337124
rect 357400 337084 357406 337096
rect 413646 337084 413652 337096
rect 413704 337084 413710 337136
rect 414658 337084 414664 337136
rect 414716 337124 414722 337136
rect 422846 337124 422852 337136
rect 414716 337096 422852 337124
rect 414716 337084 414722 337096
rect 422846 337084 422852 337096
rect 422904 337084 422910 337136
rect 423582 337084 423588 337136
rect 423640 337124 423646 337136
rect 432601 337127 432659 337133
rect 432601 337124 432613 337127
rect 423640 337096 432613 337124
rect 423640 337084 423646 337096
rect 432601 337093 432613 337096
rect 432647 337093 432659 337127
rect 451642 337124 451648 337136
rect 432601 337087 432659 337093
rect 432800 337096 451648 337124
rect 111702 337016 111708 337068
rect 111760 337056 111766 337068
rect 286870 337056 286876 337068
rect 111760 337028 286876 337056
rect 111760 337016 111766 337028
rect 286870 337016 286876 337028
rect 286928 337016 286934 337068
rect 360102 337016 360108 337068
rect 360160 337056 360166 337068
rect 414842 337056 414848 337068
rect 360160 337028 414848 337056
rect 360160 337016 360166 337028
rect 414842 337016 414848 337028
rect 414900 337016 414906 337068
rect 420178 337016 420184 337068
rect 420236 337056 420242 337068
rect 430485 337059 430543 337065
rect 430485 337056 430497 337059
rect 420236 337028 430497 337056
rect 420236 337016 420242 337028
rect 430485 337025 430497 337028
rect 430531 337025 430543 337059
rect 430485 337019 430543 337025
rect 431862 337016 431868 337068
rect 431920 337056 431926 337068
rect 432800 337056 432828 337096
rect 451642 337084 451648 337096
rect 451700 337084 451706 337136
rect 507302 337084 507308 337136
rect 507360 337124 507366 337136
rect 538214 337124 538220 337136
rect 507360 337096 538220 337124
rect 507360 337084 507366 337096
rect 538214 337084 538220 337096
rect 538272 337084 538278 337136
rect 435821 337059 435879 337065
rect 435821 337056 435833 337059
rect 431920 337028 432828 337056
rect 432892 337028 435833 337056
rect 431920 337016 431926 337028
rect 118602 336948 118608 337000
rect 118660 336988 118666 337000
rect 290550 336988 290556 337000
rect 118660 336960 290556 336988
rect 118660 336948 118666 336960
rect 290550 336948 290556 336960
rect 290608 336948 290614 337000
rect 347777 336991 347835 336997
rect 347777 336957 347789 336991
rect 347823 336988 347835 336991
rect 357345 336991 357403 336997
rect 357345 336988 357357 336991
rect 347823 336960 357357 336988
rect 347823 336957 347835 336960
rect 347777 336951 347835 336957
rect 357345 336957 357357 336960
rect 357391 336957 357403 336991
rect 357345 336951 357403 336957
rect 366450 336948 366456 337000
rect 366508 336988 366514 337000
rect 417326 336988 417332 337000
rect 366508 336960 417332 336988
rect 366508 336948 366514 336960
rect 417326 336948 417332 336960
rect 417384 336948 417390 337000
rect 424410 336948 424416 337000
rect 424468 336988 424474 337000
rect 431129 336991 431187 336997
rect 431129 336988 431141 336991
rect 424468 336960 431141 336988
rect 424468 336948 424474 336960
rect 431129 336957 431141 336960
rect 431175 336957 431187 336991
rect 431129 336951 431187 336957
rect 431218 336948 431224 337000
rect 431276 336988 431282 337000
rect 432785 336991 432843 336997
rect 431276 336960 432736 336988
rect 431276 336948 431282 336960
rect 125502 336880 125508 336932
rect 125560 336920 125566 336932
rect 294230 336920 294236 336932
rect 125560 336892 294236 336920
rect 125560 336880 125566 336892
rect 294230 336880 294236 336892
rect 294288 336880 294294 336932
rect 366358 336880 366364 336932
rect 366416 336920 366422 336932
rect 395341 336923 395399 336929
rect 395341 336920 395353 336923
rect 366416 336892 395353 336920
rect 366416 336880 366422 336892
rect 395341 336889 395353 336892
rect 395387 336889 395399 336923
rect 395341 336883 395399 336889
rect 395430 336880 395436 336932
rect 395488 336920 395494 336932
rect 400766 336920 400772 336932
rect 395488 336892 400772 336920
rect 395488 336880 395494 336892
rect 400766 336880 400772 336892
rect 400824 336880 400830 336932
rect 413370 336880 413376 336932
rect 413428 336920 413434 336932
rect 422941 336923 422999 336929
rect 422941 336920 422953 336923
rect 413428 336892 422953 336920
rect 413428 336880 413434 336892
rect 422941 336889 422953 336892
rect 422987 336889 422999 336923
rect 422941 336883 422999 336889
rect 427078 336880 427084 336932
rect 427136 336920 427142 336932
rect 432601 336923 432659 336929
rect 432601 336920 432613 336923
rect 427136 336892 432613 336920
rect 427136 336880 427142 336892
rect 432601 336889 432613 336892
rect 432647 336889 432659 336923
rect 432708 336920 432736 336960
rect 432785 336957 432797 336991
rect 432831 336988 432843 336991
rect 432892 336988 432920 337028
rect 435821 337025 435833 337028
rect 435867 337025 435879 337059
rect 435821 337019 435879 337025
rect 436002 337016 436008 337068
rect 436060 337056 436066 337068
rect 454034 337056 454040 337068
rect 436060 337028 454040 337056
rect 436060 337016 436066 337028
rect 454034 337016 454040 337028
rect 454092 337016 454098 337068
rect 482186 337016 482192 337068
rect 482244 337056 482250 337068
rect 482830 337056 482836 337068
rect 482244 337028 482836 337056
rect 482244 337016 482250 337028
rect 482830 337016 482836 337028
rect 482888 337016 482894 337068
rect 509786 337016 509792 337068
rect 509844 337056 509850 337068
rect 540330 337056 540336 337068
rect 509844 337028 540336 337056
rect 509844 337016 509850 337028
rect 540330 337016 540336 337028
rect 540388 337016 540394 337068
rect 432831 336960 432920 336988
rect 432831 336957 432843 336960
rect 432785 336951 432843 336957
rect 434622 336948 434628 337000
rect 434680 336988 434686 337000
rect 441341 336991 441399 336997
rect 441341 336988 441353 336991
rect 434680 336960 441353 336988
rect 434680 336948 434686 336960
rect 441341 336957 441353 336960
rect 441387 336957 441399 336991
rect 441341 336951 441399 336957
rect 464338 336948 464344 337000
rect 464396 336988 464402 337000
rect 466270 336988 466276 337000
rect 464396 336960 466276 336988
rect 464396 336948 464402 336960
rect 466270 336948 466276 336960
rect 466328 336948 466334 337000
rect 479150 336948 479156 337000
rect 479208 336988 479214 337000
rect 484578 336988 484584 337000
rect 479208 336960 484584 336988
rect 479208 336948 479214 336960
rect 484578 336948 484584 336960
rect 484636 336948 484642 337000
rect 516502 336948 516508 337000
rect 516560 336988 516566 337000
rect 517422 336988 517428 337000
rect 516560 336960 517428 336988
rect 516560 336948 516566 336960
rect 517422 336948 517428 336960
rect 517480 336948 517486 337000
rect 517698 336948 517704 337000
rect 517756 336988 517762 337000
rect 518802 336988 518808 337000
rect 517756 336960 518808 336988
rect 517756 336948 517762 336960
rect 518802 336948 518808 336960
rect 518860 336948 518866 337000
rect 518986 336948 518992 337000
rect 519044 336988 519050 337000
rect 520090 336988 520096 337000
rect 519044 336960 520096 336988
rect 519044 336948 519050 336960
rect 520090 336948 520096 336960
rect 520148 336948 520154 337000
rect 520185 336991 520243 336997
rect 520185 336957 520197 336991
rect 520231 336988 520243 336991
rect 545758 336988 545764 337000
rect 520231 336960 545764 336988
rect 520231 336957 520243 336960
rect 520185 336951 520243 336957
rect 545758 336948 545764 336960
rect 545816 336948 545822 337000
rect 440602 336920 440608 336932
rect 432708 336892 440608 336920
rect 432601 336883 432659 336889
rect 440602 336880 440608 336892
rect 440660 336880 440666 336932
rect 453482 336920 453488 336932
rect 447152 336892 453488 336920
rect 105538 336812 105544 336864
rect 105596 336852 105602 336864
rect 274082 336852 274088 336864
rect 105596 336824 274088 336852
rect 105596 336812 105602 336824
rect 274082 336812 274088 336824
rect 274140 336812 274146 336864
rect 363598 336812 363604 336864
rect 363656 336852 363662 336864
rect 398926 336852 398932 336864
rect 363656 336824 398932 336852
rect 363656 336812 363662 336824
rect 398926 336812 398932 336824
rect 398984 336812 398990 336864
rect 404446 336852 404452 336864
rect 400876 336824 404452 336852
rect 106918 336744 106924 336796
rect 106976 336784 106982 336796
rect 268562 336784 268568 336796
rect 106976 336756 267044 336784
rect 106976 336744 106982 336756
rect 267016 336716 267044 336756
rect 267660 336756 268568 336784
rect 267660 336716 267688 336756
rect 268562 336744 268568 336756
rect 268620 336744 268626 336796
rect 347958 336744 347964 336796
rect 348016 336784 348022 336796
rect 348786 336784 348792 336796
rect 348016 336756 348792 336784
rect 348016 336744 348022 336756
rect 348786 336744 348792 336756
rect 348844 336744 348850 336796
rect 363690 336744 363696 336796
rect 363748 336784 363754 336796
rect 377033 336787 377091 336793
rect 377033 336784 377045 336787
rect 363748 336756 377045 336784
rect 363748 336744 363754 336756
rect 377033 336753 377045 336756
rect 377079 336753 377091 336787
rect 379425 336787 379483 336793
rect 379425 336784 379437 336787
rect 377033 336747 377091 336753
rect 377140 336756 379437 336784
rect 267016 336688 267688 336716
rect 356514 336676 356520 336728
rect 356572 336716 356578 336728
rect 356698 336716 356704 336728
rect 356572 336688 356704 336716
rect 356572 336676 356578 336688
rect 356698 336676 356704 336688
rect 356756 336676 356762 336728
rect 367097 336719 367155 336725
rect 367097 336685 367109 336719
rect 367143 336716 367155 336719
rect 377140 336716 377168 336756
rect 379425 336753 379437 336756
rect 379471 336753 379483 336787
rect 379425 336747 379483 336753
rect 381538 336744 381544 336796
rect 381596 336784 381602 336796
rect 382458 336784 382464 336796
rect 381596 336756 382464 336784
rect 381596 336744 381602 336756
rect 382458 336744 382464 336756
rect 382516 336744 382522 336796
rect 382918 336744 382924 336796
rect 382976 336784 382982 336796
rect 386138 336784 386144 336796
rect 382976 336756 386144 336784
rect 382976 336744 382982 336756
rect 386138 336744 386144 336756
rect 386196 336744 386202 336796
rect 389910 336744 389916 336796
rect 389968 336784 389974 336796
rect 393406 336784 393412 336796
rect 389968 336756 393412 336784
rect 389968 336744 389974 336756
rect 393406 336744 393412 336756
rect 393464 336744 393470 336796
rect 396718 336744 396724 336796
rect 396776 336784 396782 336796
rect 400876 336784 400904 336824
rect 404446 336812 404452 336824
rect 404504 336812 404510 336864
rect 410610 336812 410616 336864
rect 410668 336852 410674 336864
rect 416406 336852 416412 336864
rect 410668 336824 416412 336852
rect 410668 336812 410674 336824
rect 416406 336812 416412 336824
rect 416464 336812 416470 336864
rect 421009 336855 421067 336861
rect 421009 336821 421021 336855
rect 421055 336852 421067 336855
rect 427722 336852 427728 336864
rect 421055 336824 427728 336852
rect 421055 336821 421067 336824
rect 421009 336815 421067 336821
rect 427722 336812 427728 336824
rect 427780 336812 427786 336864
rect 429102 336812 429108 336864
rect 429160 336852 429166 336864
rect 433429 336855 433487 336861
rect 433429 336852 433441 336855
rect 429160 336824 433441 336852
rect 429160 336812 429166 336824
rect 433429 336821 433441 336824
rect 433475 336821 433487 336855
rect 433429 336815 433487 336821
rect 435358 336812 435364 336864
rect 435416 336852 435422 336864
rect 442442 336852 442448 336864
rect 435416 336824 442448 336852
rect 435416 336812 435422 336824
rect 442442 336812 442448 336824
rect 442500 336812 442506 336864
rect 396776 336756 400904 336784
rect 396776 336744 396782 336756
rect 401042 336744 401048 336796
rect 401100 336784 401106 336796
rect 408126 336784 408132 336796
rect 401100 336756 408132 336784
rect 401100 336744 401106 336756
rect 408126 336744 408132 336756
rect 408184 336744 408190 336796
rect 410518 336744 410524 336796
rect 410576 336784 410582 336796
rect 413002 336784 413008 336796
rect 410576 336756 413008 336784
rect 410576 336744 410582 336756
rect 413002 336744 413008 336756
rect 413060 336744 413066 336796
rect 416038 336744 416044 336796
rect 416096 336784 416102 336796
rect 424226 336784 424232 336796
rect 416096 336756 424232 336784
rect 416096 336744 416102 336756
rect 424226 336744 424232 336756
rect 424284 336744 424290 336796
rect 424318 336744 424324 336796
rect 424376 336784 424382 336796
rect 425882 336784 425888 336796
rect 424376 336756 425888 336784
rect 424376 336744 424382 336756
rect 425882 336744 425888 336756
rect 425940 336744 425946 336796
rect 430482 336744 430488 336796
rect 430540 336784 430546 336796
rect 432509 336787 432567 336793
rect 432509 336784 432521 336787
rect 430540 336756 432521 336784
rect 430540 336744 430546 336756
rect 432509 336753 432521 336756
rect 432555 336753 432567 336787
rect 432509 336747 432567 336753
rect 432601 336787 432659 336793
rect 432601 336753 432613 336787
rect 432647 336784 432659 336787
rect 437474 336784 437480 336796
rect 432647 336756 437480 336784
rect 432647 336753 432659 336756
rect 432601 336747 432659 336753
rect 437474 336744 437480 336756
rect 437532 336744 437538 336796
rect 438118 336744 438124 336796
rect 438176 336784 438182 336796
rect 444282 336784 444288 336796
rect 438176 336756 444288 336784
rect 438176 336744 438182 336756
rect 444282 336744 444288 336756
rect 444340 336744 444346 336796
rect 446398 336744 446404 336796
rect 446456 336784 446462 336796
rect 447152 336784 447180 336892
rect 453482 336880 453488 336892
rect 453540 336880 453546 336932
rect 462958 336880 462964 336932
rect 463016 336920 463022 336932
rect 464430 336920 464436 336932
rect 463016 336892 464436 336920
rect 463016 336880 463022 336892
rect 464430 336880 464436 336892
rect 464488 336880 464494 336932
rect 468754 336920 468760 336932
rect 467576 336892 468760 336920
rect 464982 336812 464988 336864
rect 465040 336852 465046 336864
rect 467576 336852 467604 336892
rect 468754 336880 468760 336892
rect 468812 336880 468818 336932
rect 476758 336880 476764 336932
rect 476816 336920 476822 336932
rect 477402 336920 477408 336932
rect 476816 336892 477408 336920
rect 476816 336880 476822 336892
rect 477402 336880 477408 336892
rect 477460 336880 477466 336932
rect 478506 336880 478512 336932
rect 478564 336920 478570 336932
rect 483198 336920 483204 336932
rect 478564 336892 483204 336920
rect 478564 336880 478570 336892
rect 483198 336880 483204 336892
rect 483256 336880 483262 336932
rect 498746 336880 498752 336932
rect 498804 336920 498810 336932
rect 499482 336920 499488 336932
rect 498804 336892 499488 336920
rect 498804 336880 498810 336892
rect 499482 336880 499488 336892
rect 499540 336880 499546 336932
rect 504910 336880 504916 336932
rect 504968 336920 504974 336932
rect 534074 336920 534080 336932
rect 504968 336892 534080 336920
rect 504968 336880 504974 336892
rect 534074 336880 534080 336892
rect 534132 336880 534138 336932
rect 465040 336824 467604 336852
rect 465040 336812 465046 336824
rect 467742 336812 467748 336864
rect 467800 336852 467806 336864
rect 469950 336852 469956 336864
rect 467800 336824 469956 336852
rect 467800 336812 467806 336824
rect 469950 336812 469956 336824
rect 470008 336812 470014 336864
rect 480990 336812 480996 336864
rect 481048 336852 481054 336864
rect 485038 336852 485044 336864
rect 481048 336824 485044 336852
rect 481048 336812 481054 336824
rect 485038 336812 485044 336824
rect 485096 336812 485102 336864
rect 513466 336812 513472 336864
rect 513524 336852 513530 336864
rect 542998 336852 543004 336864
rect 513524 336824 543004 336852
rect 513524 336812 513530 336824
rect 542998 336812 543004 336824
rect 543056 336812 543062 336864
rect 446456 336756 447180 336784
rect 446456 336744 446462 336756
rect 447778 336744 447784 336796
rect 447836 336784 447842 336796
rect 455322 336784 455328 336796
rect 447836 336756 455328 336784
rect 447836 336744 447842 336756
rect 455322 336744 455328 336756
rect 455380 336744 455386 336796
rect 460198 336744 460204 336796
rect 460256 336784 460262 336796
rect 462590 336784 462596 336796
rect 460256 336756 462596 336784
rect 460256 336744 460262 336756
rect 462590 336744 462596 336756
rect 462648 336744 462654 336796
rect 464430 336744 464436 336796
rect 464488 336784 464494 336796
rect 465718 336784 465724 336796
rect 464488 336756 465724 336784
rect 464488 336744 464494 336756
rect 465718 336744 465724 336756
rect 465776 336744 465782 336796
rect 469858 336744 469864 336796
rect 469916 336784 469922 336796
rect 471238 336784 471244 336796
rect 469916 336756 471244 336784
rect 469916 336744 469922 336756
rect 471238 336744 471244 336756
rect 471296 336744 471302 336796
rect 474918 336744 474924 336796
rect 474976 336784 474982 336796
rect 476022 336784 476028 336796
rect 474976 336756 476028 336784
rect 474976 336744 474982 336756
rect 476022 336744 476028 336756
rect 476080 336744 476086 336796
rect 476114 336744 476120 336796
rect 476172 336784 476178 336796
rect 477586 336784 477592 336796
rect 476172 336756 477592 336784
rect 476172 336744 476178 336756
rect 477586 336744 477592 336756
rect 477644 336744 477650 336796
rect 477954 336744 477960 336796
rect 478012 336784 478018 336796
rect 478782 336784 478788 336796
rect 478012 336756 478788 336784
rect 478012 336744 478018 336756
rect 478782 336744 478788 336756
rect 478840 336744 478846 336796
rect 480346 336744 480352 336796
rect 480404 336784 480410 336796
rect 481542 336784 481548 336796
rect 480404 336756 481548 336784
rect 480404 336744 480410 336756
rect 481542 336744 481548 336756
rect 481600 336744 481606 336796
rect 481634 336744 481640 336796
rect 481692 336784 481698 336796
rect 482922 336784 482928 336796
rect 481692 336756 482928 336784
rect 481692 336744 481698 336756
rect 482922 336744 482928 336756
rect 482980 336744 482986 336796
rect 483474 336744 483480 336796
rect 483532 336784 483538 336796
rect 484302 336784 484308 336796
rect 483532 336756 484308 336784
rect 483532 336744 483538 336756
rect 484302 336744 484308 336756
rect 484360 336744 484366 336796
rect 484670 336744 484676 336796
rect 484728 336784 484734 336796
rect 485682 336784 485688 336796
rect 484728 336756 485688 336784
rect 484728 336744 484734 336756
rect 485682 336744 485688 336756
rect 485740 336744 485746 336796
rect 503438 336744 503444 336796
rect 503496 336784 503502 336796
rect 524417 336787 524475 336793
rect 524417 336784 524429 336787
rect 503496 336756 524429 336784
rect 503496 336744 503502 336756
rect 524417 336753 524429 336756
rect 524463 336753 524475 336787
rect 524417 336747 524475 336753
rect 524506 336744 524512 336796
rect 524564 336784 524570 336796
rect 525610 336784 525616 336796
rect 524564 336756 525616 336784
rect 524564 336744 524570 336756
rect 525610 336744 525616 336756
rect 525668 336744 525674 336796
rect 526346 336744 526352 336796
rect 526404 336784 526410 336796
rect 526404 336756 527496 336784
rect 526404 336744 526410 336756
rect 382642 336716 382648 336728
rect 367143 336688 377168 336716
rect 382476 336688 382648 336716
rect 367143 336685 367155 336688
rect 367097 336679 367155 336685
rect 382476 336660 382504 336688
rect 382642 336676 382648 336688
rect 382700 336676 382706 336728
rect 527468 336716 527496 336756
rect 527542 336744 527548 336796
rect 527600 336784 527606 336796
rect 528462 336784 528468 336796
rect 527600 336756 528468 336784
rect 527600 336744 527606 336756
rect 528462 336744 528468 336756
rect 528520 336744 528526 336796
rect 528738 336744 528744 336796
rect 528796 336784 528802 336796
rect 529842 336784 529848 336796
rect 528796 336756 529848 336784
rect 528796 336744 528802 336756
rect 529842 336744 529848 336756
rect 529900 336744 529906 336796
rect 531501 336787 531559 336793
rect 531501 336784 531513 336787
rect 529952 336756 531513 336784
rect 529952 336716 529980 336756
rect 531501 336753 531513 336756
rect 531547 336753 531559 336787
rect 531501 336747 531559 336753
rect 527468 336688 529980 336716
rect 382458 336608 382464 336660
rect 382516 336608 382522 336660
rect 230658 335588 230664 335640
rect 230716 335628 230722 335640
rect 231486 335628 231492 335640
rect 230716 335600 231492 335628
rect 230716 335588 230722 335600
rect 231486 335588 231492 335600
rect 231544 335588 231550 335640
rect 237466 335588 237472 335640
rect 237524 335628 237530 335640
rect 238294 335628 238300 335640
rect 237524 335600 238300 335628
rect 237524 335588 237530 335600
rect 238294 335588 238300 335600
rect 238352 335588 238358 335640
rect 241514 335588 241520 335640
rect 241572 335628 241578 335640
rect 241974 335628 241980 335640
rect 241572 335600 241980 335628
rect 241572 335588 241578 335600
rect 241974 335588 241980 335600
rect 242032 335588 242038 335640
rect 243078 335588 243084 335640
rect 243136 335628 243142 335640
rect 243814 335628 243820 335640
rect 243136 335600 243820 335628
rect 243136 335588 243142 335600
rect 243814 335588 243820 335600
rect 243872 335588 243878 335640
rect 245654 335588 245660 335640
rect 245712 335628 245718 335640
rect 246206 335628 246212 335640
rect 245712 335600 246212 335628
rect 245712 335588 245718 335600
rect 246206 335588 246212 335600
rect 246264 335588 246270 335640
rect 248414 335588 248420 335640
rect 248472 335628 248478 335640
rect 249150 335628 249156 335640
rect 248472 335600 249156 335628
rect 248472 335588 248478 335600
rect 249150 335588 249156 335600
rect 249208 335588 249214 335640
rect 302326 335588 302332 335640
rect 302384 335628 302390 335640
rect 303062 335628 303068 335640
rect 302384 335600 303068 335628
rect 302384 335588 302390 335600
rect 303062 335588 303068 335600
rect 303120 335588 303126 335640
rect 303614 335588 303620 335640
rect 303672 335628 303678 335640
rect 304350 335628 304356 335640
rect 303672 335600 304356 335628
rect 303672 335588 303678 335600
rect 304350 335588 304356 335600
rect 304408 335588 304414 335640
rect 307846 335588 307852 335640
rect 307904 335628 307910 335640
rect 308030 335628 308036 335640
rect 307904 335600 308036 335628
rect 307904 335588 307910 335600
rect 308030 335588 308036 335600
rect 308088 335588 308094 335640
rect 310698 335588 310704 335640
rect 310756 335628 310762 335640
rect 311158 335628 311164 335640
rect 310756 335600 311164 335628
rect 310756 335588 310762 335600
rect 311158 335588 311164 335600
rect 311216 335588 311222 335640
rect 323118 335588 323124 335640
rect 323176 335628 323182 335640
rect 323854 335628 323860 335640
rect 323176 335600 323860 335628
rect 323176 335588 323182 335600
rect 323854 335588 323860 335600
rect 323912 335588 323918 335640
rect 325694 335588 325700 335640
rect 325752 335628 325758 335640
rect 326430 335628 326436 335640
rect 325752 335600 326436 335628
rect 325752 335588 325758 335600
rect 326430 335588 326436 335600
rect 326488 335588 326494 335640
rect 328638 335588 328644 335640
rect 328696 335628 328702 335640
rect 329374 335628 329380 335640
rect 328696 335600 329380 335628
rect 328696 335588 328702 335600
rect 329374 335588 329380 335600
rect 329432 335588 329438 335640
rect 335354 335588 335360 335640
rect 335412 335628 335418 335640
rect 336182 335628 336188 335640
rect 335412 335600 336188 335628
rect 335412 335588 335418 335600
rect 336182 335588 336188 335600
rect 336240 335588 336246 335640
rect 340874 335588 340880 335640
rect 340932 335628 340938 335640
rect 341702 335628 341708 335640
rect 340932 335600 341708 335628
rect 340932 335588 340938 335600
rect 341702 335588 341708 335600
rect 341760 335588 341766 335640
rect 345014 335588 345020 335640
rect 345072 335628 345078 335640
rect 345934 335628 345940 335640
rect 345072 335600 345940 335628
rect 345072 335588 345078 335600
rect 345934 335588 345940 335600
rect 345992 335588 345998 335640
rect 349154 335588 349160 335640
rect 349212 335628 349218 335640
rect 349614 335628 349620 335640
rect 349212 335600 349620 335628
rect 349212 335588 349218 335600
rect 349614 335588 349620 335600
rect 349672 335588 349678 335640
rect 350534 335588 350540 335640
rect 350592 335628 350598 335640
rect 351454 335628 351460 335640
rect 350592 335600 351460 335628
rect 350592 335588 350598 335600
rect 351454 335588 351460 335600
rect 351512 335588 351518 335640
rect 354674 335588 354680 335640
rect 354732 335628 354738 335640
rect 355134 335628 355140 335640
rect 354732 335600 355140 335628
rect 354732 335588 354738 335600
rect 355134 335588 355140 335600
rect 355192 335588 355198 335640
rect 357618 335588 357624 335640
rect 357676 335628 357682 335640
rect 358262 335628 358268 335640
rect 357676 335600 358268 335628
rect 357676 335588 357682 335600
rect 358262 335588 358268 335600
rect 358320 335588 358326 335640
rect 360194 335588 360200 335640
rect 360252 335628 360258 335640
rect 360654 335628 360660 335640
rect 360252 335600 360660 335628
rect 360252 335588 360258 335600
rect 360654 335588 360660 335600
rect 360712 335588 360718 335640
rect 361666 335588 361672 335640
rect 361724 335628 361730 335640
rect 362494 335628 362500 335640
rect 361724 335600 362500 335628
rect 361724 335588 361730 335600
rect 362494 335588 362500 335600
rect 362552 335588 362558 335640
rect 362954 335588 362960 335640
rect 363012 335628 363018 335640
rect 363782 335628 363788 335640
rect 363012 335600 363788 335628
rect 363012 335588 363018 335600
rect 363782 335588 363788 335600
rect 363840 335588 363846 335640
rect 377030 335628 377036 335640
rect 376991 335600 377036 335628
rect 377030 335588 377036 335600
rect 377088 335588 377094 335640
rect 378226 335588 378232 335640
rect 378284 335628 378290 335640
rect 379054 335628 379060 335640
rect 378284 335600 379060 335628
rect 378284 335588 378290 335600
rect 379054 335588 379060 335600
rect 379112 335588 379118 335640
rect 405918 335588 405924 335640
rect 405976 335628 405982 335640
rect 406654 335628 406660 335640
rect 405976 335600 406660 335628
rect 405976 335588 405982 335600
rect 406654 335588 406660 335600
rect 406712 335588 406718 335640
rect 422294 335588 422300 335640
rect 422352 335628 422358 335640
rect 423214 335628 423220 335640
rect 422352 335600 423220 335628
rect 422352 335588 422358 335600
rect 423214 335588 423220 335600
rect 423272 335588 423278 335640
rect 430574 335588 430580 335640
rect 430632 335628 430638 335640
rect 431126 335628 431132 335640
rect 430632 335600 431132 335628
rect 430632 335588 430638 335600
rect 431126 335588 431132 335600
rect 431184 335588 431190 335640
rect 334066 335384 334072 335436
rect 334124 335424 334130 335436
rect 334124 335396 334204 335424
rect 334124 335384 334130 335396
rect 318978 335316 318984 335368
rect 319036 335356 319042 335368
rect 319622 335356 319628 335368
rect 319036 335328 319628 335356
rect 319036 335316 319042 335328
rect 319622 335316 319628 335328
rect 319680 335316 319686 335368
rect 294049 335291 294107 335297
rect 294049 335257 294061 335291
rect 294095 335288 294107 335291
rect 294506 335288 294512 335300
rect 294095 335260 294512 335288
rect 294095 335257 294107 335260
rect 294049 335251 294107 335257
rect 294506 335248 294512 335260
rect 294564 335248 294570 335300
rect 334176 335232 334204 335396
rect 356514 335288 356520 335300
rect 356475 335260 356520 335288
rect 356514 335248 356520 335260
rect 356572 335248 356578 335300
rect 334158 335180 334164 335232
rect 334216 335180 334222 335232
rect 252738 334568 252744 334620
rect 252796 334608 252802 334620
rect 253290 334608 253296 334620
rect 252796 334580 253296 334608
rect 252796 334568 252802 334580
rect 253290 334568 253296 334580
rect 253348 334568 253354 334620
rect 296806 334432 296812 334484
rect 296864 334472 296870 334484
rect 297542 334472 297548 334484
rect 296864 334444 297548 334472
rect 296864 334432 296870 334444
rect 297542 334432 297548 334444
rect 297600 334432 297606 334484
rect 427998 334296 428004 334348
rect 428056 334336 428062 334348
rect 428458 334336 428464 334348
rect 428056 334308 428464 334336
rect 428056 334296 428062 334308
rect 428458 334296 428464 334308
rect 428516 334296 428522 334348
rect 299474 333888 299480 333940
rect 299532 333928 299538 333940
rect 300118 333928 300124 333940
rect 299532 333900 300124 333928
rect 299532 333888 299538 333900
rect 300118 333888 300124 333900
rect 300176 333888 300182 333940
rect 259638 333276 259644 333328
rect 259696 333316 259702 333328
rect 260282 333316 260288 333328
rect 259696 333288 260288 333316
rect 259696 333276 259702 333288
rect 260282 333276 260288 333288
rect 260340 333276 260346 333328
rect 352006 333276 352012 333328
rect 352064 333316 352070 333328
rect 352650 333316 352656 333328
rect 352064 333288 352656 333316
rect 352064 333276 352070 333288
rect 352650 333276 352656 333288
rect 352708 333276 352714 333328
rect 466546 333276 466552 333328
rect 466604 333316 466610 333328
rect 467098 333316 467104 333328
rect 466604 333288 467104 333316
rect 466604 333276 466610 333288
rect 467098 333276 467104 333288
rect 467156 333276 467162 333328
rect 339494 333208 339500 333260
rect 339552 333248 339558 333260
rect 340414 333248 340420 333260
rect 339552 333220 340420 333248
rect 339552 333208 339558 333220
rect 340414 333208 340420 333220
rect 340472 333208 340478 333260
rect 343634 332188 343640 332240
rect 343692 332228 343698 332240
rect 344094 332228 344100 332240
rect 343692 332200 344100 332228
rect 343692 332188 343698 332200
rect 344094 332188 344100 332200
rect 344152 332188 344158 332240
rect 306374 331916 306380 331968
rect 306432 331956 306438 331968
rect 306742 331956 306748 331968
rect 306432 331928 306748 331956
rect 306432 331916 306438 331928
rect 306742 331916 306748 331928
rect 306800 331916 306806 331968
rect 324406 331848 324412 331900
rect 324464 331888 324470 331900
rect 325050 331888 325056 331900
rect 324464 331860 325056 331888
rect 324464 331848 324470 331860
rect 325050 331848 325056 331860
rect 325108 331848 325114 331900
rect 327258 331848 327264 331900
rect 327316 331888 327322 331900
rect 327442 331888 327448 331900
rect 327316 331860 327448 331888
rect 327316 331848 327322 331860
rect 327442 331848 327448 331860
rect 327500 331848 327506 331900
rect 333974 331576 333980 331628
rect 334032 331616 334038 331628
rect 334250 331616 334256 331628
rect 334032 331588 334256 331616
rect 334032 331576 334038 331588
rect 334250 331576 334256 331588
rect 334308 331576 334314 331628
rect 295794 331276 295800 331288
rect 295628 331248 295800 331276
rect 295628 331220 295656 331248
rect 295794 331236 295800 331248
rect 295852 331236 295858 331288
rect 295610 331168 295616 331220
rect 295668 331168 295674 331220
rect 305178 331168 305184 331220
rect 305236 331168 305242 331220
rect 416774 331168 416780 331220
rect 416832 331208 416838 331220
rect 416958 331208 416964 331220
rect 416832 331180 416964 331208
rect 416832 331168 416838 331180
rect 416958 331168 416964 331180
rect 417016 331168 417022 331220
rect 422294 331168 422300 331220
rect 422352 331208 422358 331220
rect 422478 331208 422484 331220
rect 422352 331180 422484 331208
rect 422352 331168 422358 331180
rect 422478 331168 422484 331180
rect 422536 331168 422542 331220
rect 305196 331140 305224 331168
rect 305270 331140 305276 331152
rect 305196 331112 305276 331140
rect 305270 331100 305276 331112
rect 305328 331100 305334 331152
rect 381170 331140 381176 331152
rect 381131 331112 381176 331140
rect 381170 331100 381176 331112
rect 381228 331100 381234 331152
rect 254210 330420 254216 330472
rect 254268 330460 254274 330472
rect 254762 330460 254768 330472
rect 254268 330432 254768 330460
rect 254268 330420 254274 330432
rect 254762 330420 254768 330432
rect 254820 330420 254826 330472
rect 371510 328556 371516 328568
rect 371344 328528 371516 328556
rect 371344 328500 371372 328528
rect 371510 328516 371516 328528
rect 371568 328516 371574 328568
rect 236270 328448 236276 328500
rect 236328 328488 236334 328500
rect 236914 328488 236920 328500
rect 236328 328460 236920 328488
rect 236328 328448 236334 328460
rect 236914 328448 236920 328460
rect 236972 328448 236978 328500
rect 241790 328448 241796 328500
rect 241848 328488 241854 328500
rect 242342 328488 242348 328500
rect 241848 328460 242348 328488
rect 241848 328448 241854 328460
rect 242342 328448 242348 328460
rect 242400 328448 242406 328500
rect 265250 328448 265256 328500
rect 265308 328488 265314 328500
rect 265618 328488 265624 328500
rect 265308 328460 265624 328488
rect 265308 328448 265314 328460
rect 265618 328448 265624 328460
rect 265676 328448 265682 328500
rect 267090 328448 267096 328500
rect 267148 328488 267154 328500
rect 267553 328491 267611 328497
rect 267553 328488 267565 328491
rect 267148 328460 267565 328488
rect 267148 328448 267154 328460
rect 267553 328457 267565 328460
rect 267599 328457 267611 328491
rect 267553 328451 267611 328457
rect 270770 328448 270776 328500
rect 270828 328488 270834 328500
rect 271138 328488 271144 328500
rect 270828 328460 271144 328488
rect 270828 328448 270834 328460
rect 271138 328448 271144 328460
rect 271196 328448 271202 328500
rect 309410 328448 309416 328500
rect 309468 328488 309474 328500
rect 309686 328488 309692 328500
rect 309468 328460 309692 328488
rect 309468 328448 309474 328460
rect 309686 328448 309692 328460
rect 309744 328448 309750 328500
rect 330018 328448 330024 328500
rect 330076 328488 330082 328500
rect 330570 328488 330576 328500
rect 330076 328460 330576 328488
rect 330076 328448 330082 328460
rect 330570 328448 330576 328460
rect 330628 328448 330634 328500
rect 331490 328448 331496 328500
rect 331548 328488 331554 328500
rect 331674 328488 331680 328500
rect 331548 328460 331680 328488
rect 331548 328448 331554 328460
rect 331674 328448 331680 328460
rect 331732 328448 331738 328500
rect 334434 328448 334440 328500
rect 334492 328488 334498 328500
rect 334802 328488 334808 328500
rect 334492 328460 334808 328488
rect 334492 328448 334498 328460
rect 334802 328448 334808 328460
rect 334860 328448 334866 328500
rect 336918 328448 336924 328500
rect 336976 328488 336982 328500
rect 337194 328488 337200 328500
rect 336976 328460 337200 328488
rect 336976 328448 336982 328460
rect 337194 328448 337200 328460
rect 337252 328448 337258 328500
rect 342622 328448 342628 328500
rect 342680 328488 342686 328500
rect 342990 328488 342996 328500
rect 342680 328460 342996 328488
rect 342680 328448 342686 328460
rect 342990 328448 342996 328460
rect 343048 328448 343054 328500
rect 353570 328448 353576 328500
rect 353628 328488 353634 328500
rect 353938 328488 353944 328500
rect 353628 328460 353944 328488
rect 353628 328448 353634 328460
rect 353938 328448 353944 328460
rect 353996 328448 354002 328500
rect 359090 328448 359096 328500
rect 359148 328488 359154 328500
rect 359458 328488 359464 328500
rect 359148 328460 359464 328488
rect 359148 328448 359154 328460
rect 359458 328448 359464 328460
rect 359516 328448 359522 328500
rect 364610 328448 364616 328500
rect 364668 328488 364674 328500
rect 364794 328488 364800 328500
rect 364668 328460 364800 328488
rect 364668 328448 364674 328460
rect 364794 328448 364800 328460
rect 364852 328448 364858 328500
rect 367278 328448 367284 328500
rect 367336 328488 367342 328500
rect 367830 328488 367836 328500
rect 367336 328460 367836 328488
rect 367336 328448 367342 328460
rect 367830 328448 367836 328460
rect 367888 328448 367894 328500
rect 370130 328448 370136 328500
rect 370188 328488 370194 328500
rect 370314 328488 370320 328500
rect 370188 328460 370320 328488
rect 370188 328448 370194 328460
rect 370314 328448 370320 328460
rect 370372 328448 370378 328500
rect 371326 328448 371332 328500
rect 371384 328448 371390 328500
rect 381078 328448 381084 328500
rect 381136 328488 381142 328500
rect 381173 328491 381231 328497
rect 381173 328488 381185 328491
rect 381136 328460 381185 328488
rect 381136 328448 381142 328460
rect 381173 328457 381185 328460
rect 381219 328457 381231 328491
rect 381173 328451 381231 328457
rect 386690 328448 386696 328500
rect 386748 328488 386754 328500
rect 386874 328488 386880 328500
rect 386748 328460 386880 328488
rect 386748 328448 386754 328460
rect 386874 328448 386880 328460
rect 386932 328448 386938 328500
rect 232222 328380 232228 328432
rect 232280 328420 232286 328432
rect 232314 328420 232320 328432
rect 232280 328392 232320 328420
rect 232280 328380 232286 328392
rect 232314 328380 232320 328392
rect 232372 328380 232378 328432
rect 392302 328420 392308 328432
rect 392263 328392 392308 328420
rect 392302 328380 392308 328392
rect 392360 328380 392366 328432
rect 393222 328420 393228 328432
rect 393183 328392 393228 328420
rect 393222 328380 393228 328392
rect 393280 328380 393286 328432
rect 397822 328420 397828 328432
rect 397783 328392 397828 328420
rect 397822 328380 397828 328392
rect 397880 328380 397886 328432
rect 400306 328380 400312 328432
rect 400364 328420 400370 328432
rect 400582 328420 400588 328432
rect 400364 328392 400588 328420
rect 400364 328380 400370 328392
rect 400582 328380 400588 328392
rect 400640 328380 400646 328432
rect 416869 328423 416927 328429
rect 416869 328389 416881 328423
rect 416915 328420 416927 328423
rect 416958 328420 416964 328432
rect 416915 328392 416964 328420
rect 416915 328389 416927 328392
rect 416869 328383 416927 328389
rect 416958 328380 416964 328392
rect 417016 328380 417022 328432
rect 422389 328423 422447 328429
rect 422389 328389 422401 328423
rect 422435 328420 422447 328423
rect 422478 328420 422484 328432
rect 422435 328392 422484 328420
rect 422435 328389 422447 328392
rect 422389 328383 422447 328389
rect 422478 328380 422484 328392
rect 422536 328380 422542 328432
rect 427909 328423 427967 328429
rect 427909 328389 427921 328423
rect 427955 328420 427967 328423
rect 427998 328420 428004 328432
rect 427955 328392 428004 328420
rect 427955 328389 427967 328392
rect 427909 328383 427967 328389
rect 427998 328380 428004 328392
rect 428056 328380 428062 328432
rect 433702 328420 433708 328432
rect 433663 328392 433708 328420
rect 433702 328380 433708 328392
rect 433760 328380 433766 328432
rect 472069 328423 472127 328429
rect 472069 328389 472081 328423
rect 472115 328420 472127 328423
rect 472158 328420 472164 328432
rect 472115 328392 472164 328420
rect 472115 328389 472127 328392
rect 472069 328383 472127 328389
rect 472158 328380 472164 328392
rect 472216 328380 472222 328432
rect 377030 327128 377036 327140
rect 376991 327100 377036 327128
rect 377030 327088 377036 327100
rect 377088 327088 377094 327140
rect 477310 327088 477316 327140
rect 477368 327128 477374 327140
rect 480346 327128 480352 327140
rect 477368 327100 480352 327128
rect 477368 327088 477374 327100
rect 480346 327088 480352 327100
rect 480404 327088 480410 327140
rect 281626 327020 281632 327072
rect 281684 327060 281690 327072
rect 281994 327060 282000 327072
rect 281684 327032 282000 327060
rect 281684 327020 281690 327032
rect 281994 327020 282000 327032
rect 282052 327020 282058 327072
rect 292758 327060 292764 327072
rect 292719 327032 292764 327060
rect 292758 327020 292764 327032
rect 292816 327020 292822 327072
rect 357529 327063 357587 327069
rect 357529 327029 357541 327063
rect 357575 327060 357587 327063
rect 357618 327060 357624 327072
rect 357575 327032 357624 327060
rect 357575 327029 357587 327032
rect 357529 327023 357587 327029
rect 357618 327020 357624 327032
rect 357676 327020 357682 327072
rect 382458 327060 382464 327072
rect 382419 327032 382464 327060
rect 382458 327020 382464 327032
rect 382516 327020 382522 327072
rect 400306 327060 400312 327072
rect 400267 327032 400312 327060
rect 400306 327020 400312 327032
rect 400364 327020 400370 327072
rect 294046 325700 294052 325712
rect 294007 325672 294052 325700
rect 294046 325660 294052 325672
rect 294104 325660 294110 325712
rect 321646 325660 321652 325712
rect 321704 325700 321710 325712
rect 322106 325700 322112 325712
rect 321704 325672 322112 325700
rect 321704 325660 321710 325672
rect 322106 325660 322112 325672
rect 322164 325660 322170 325712
rect 451366 325660 451372 325712
rect 451424 325700 451430 325712
rect 451550 325700 451556 325712
rect 451424 325672 451556 325700
rect 451424 325660 451430 325672
rect 451550 325660 451556 325672
rect 451608 325660 451614 325712
rect 348050 324300 348056 324352
rect 348108 324340 348114 324352
rect 348234 324340 348240 324352
rect 348108 324312 348240 324340
rect 348108 324300 348114 324312
rect 348234 324300 348240 324312
rect 348292 324300 348298 324352
rect 232314 324272 232320 324284
rect 232275 324244 232320 324272
rect 232314 324232 232320 324244
rect 232372 324232 232378 324284
rect 277302 323552 277308 323604
rect 277360 323592 277366 323604
rect 277578 323592 277584 323604
rect 277360 323564 277584 323592
rect 277360 323552 277366 323564
rect 277578 323552 277584 323564
rect 277636 323552 277642 323604
rect 530670 322872 530676 322924
rect 530728 322912 530734 322924
rect 579614 322912 579620 322924
rect 530728 322884 579620 322912
rect 530728 322872 530734 322884
rect 579614 322872 579620 322884
rect 579672 322872 579678 322924
rect 249978 321688 249984 321700
rect 249939 321660 249984 321688
rect 249978 321648 249984 321660
rect 250036 321648 250042 321700
rect 261018 321648 261024 321700
rect 261076 321648 261082 321700
rect 259638 321620 259644 321632
rect 259599 321592 259644 321620
rect 259638 321580 259644 321592
rect 259696 321580 259702 321632
rect 261036 321564 261064 321648
rect 327258 321580 327264 321632
rect 327316 321580 327322 321632
rect 348050 321620 348056 321632
rect 347976 321592 348056 321620
rect 261018 321512 261024 321564
rect 261076 321512 261082 321564
rect 327276 321496 327304 321580
rect 347976 321564 348004 321592
rect 348050 321580 348056 321592
rect 348108 321580 348114 321632
rect 359090 321620 359096 321632
rect 359016 321592 359096 321620
rect 359016 321564 359044 321592
rect 359090 321580 359096 321592
rect 359148 321580 359154 321632
rect 387978 321580 387984 321632
rect 388036 321580 388042 321632
rect 408678 321580 408684 321632
rect 408736 321580 408742 321632
rect 466546 321620 466552 321632
rect 466507 321592 466552 321620
rect 466546 321580 466552 321592
rect 466604 321580 466610 321632
rect 347958 321512 347964 321564
rect 348016 321512 348022 321564
rect 358998 321512 359004 321564
rect 359056 321512 359062 321564
rect 327258 321444 327264 321496
rect 327316 321444 327322 321496
rect 387996 321416 388024 321580
rect 408696 321484 408724 321580
rect 408770 321484 408776 321496
rect 408696 321456 408776 321484
rect 408770 321444 408776 321456
rect 408828 321444 408834 321496
rect 388070 321416 388076 321428
rect 387996 321388 388076 321416
rect 388070 321376 388076 321388
rect 388128 321376 388134 321428
rect 252738 318900 252744 318912
rect 252572 318872 252744 318900
rect 252572 318844 252600 318872
rect 252738 318860 252744 318872
rect 252796 318860 252802 318912
rect 233418 318792 233424 318844
rect 233476 318832 233482 318844
rect 233510 318832 233516 318844
rect 233476 318804 233516 318832
rect 233476 318792 233482 318804
rect 233510 318792 233516 318804
rect 233568 318792 233574 318844
rect 236270 318792 236276 318844
rect 236328 318832 236334 318844
rect 236362 318832 236368 318844
rect 236328 318804 236368 318832
rect 236328 318792 236334 318804
rect 236362 318792 236368 318804
rect 236420 318792 236426 318844
rect 252554 318792 252560 318844
rect 252612 318792 252618 318844
rect 259638 318832 259644 318844
rect 259599 318804 259644 318832
rect 259638 318792 259644 318804
rect 259696 318792 259702 318844
rect 375558 318792 375564 318844
rect 375616 318832 375622 318844
rect 375742 318832 375748 318844
rect 375616 318804 375748 318832
rect 375616 318792 375622 318804
rect 375742 318792 375748 318804
rect 375800 318792 375806 318844
rect 376938 318792 376944 318844
rect 376996 318832 377002 318844
rect 377030 318832 377036 318844
rect 376996 318804 377036 318832
rect 376996 318792 377002 318804
rect 377030 318792 377036 318804
rect 377088 318792 377094 318844
rect 392305 318835 392363 318841
rect 392305 318801 392317 318835
rect 392351 318832 392363 318835
rect 392394 318832 392400 318844
rect 392351 318804 392400 318832
rect 392351 318801 392363 318804
rect 392305 318795 392363 318801
rect 392394 318792 392400 318804
rect 392452 318792 392458 318844
rect 393222 318832 393228 318844
rect 393183 318804 393228 318832
rect 393222 318792 393228 318804
rect 393280 318792 393286 318844
rect 397825 318835 397883 318841
rect 397825 318801 397837 318835
rect 397871 318832 397883 318835
rect 397914 318832 397920 318844
rect 397871 318804 397920 318832
rect 397871 318801 397883 318804
rect 397825 318795 397883 318801
rect 397914 318792 397920 318804
rect 397972 318792 397978 318844
rect 400309 318835 400367 318841
rect 400309 318801 400321 318835
rect 400355 318832 400367 318835
rect 400490 318832 400496 318844
rect 400355 318804 400496 318832
rect 400355 318801 400367 318804
rect 400309 318795 400367 318801
rect 400490 318792 400496 318804
rect 400548 318792 400554 318844
rect 416866 318832 416872 318844
rect 416827 318804 416872 318832
rect 416866 318792 416872 318804
rect 416924 318792 416930 318844
rect 422386 318832 422392 318844
rect 422347 318804 422392 318832
rect 422386 318792 422392 318804
rect 422444 318792 422450 318844
rect 427906 318832 427912 318844
rect 427867 318804 427912 318832
rect 427906 318792 427912 318804
rect 427964 318792 427970 318844
rect 433705 318835 433763 318841
rect 433705 318801 433717 318835
rect 433751 318832 433763 318835
rect 433794 318832 433800 318844
rect 433751 318804 433800 318832
rect 433751 318801 433763 318804
rect 433705 318795 433763 318801
rect 433794 318792 433800 318804
rect 433852 318792 433858 318844
rect 466546 318832 466552 318844
rect 466507 318804 466552 318832
rect 466546 318792 466552 318804
rect 466604 318792 466610 318844
rect 472066 318832 472072 318844
rect 472027 318804 472072 318832
rect 472066 318792 472072 318804
rect 472124 318792 472130 318844
rect 283006 318724 283012 318776
rect 283064 318764 283070 318776
rect 283098 318764 283104 318776
rect 283064 318736 283104 318764
rect 283064 318724 283070 318736
rect 283098 318724 283104 318736
rect 283156 318724 283162 318776
rect 288618 318764 288624 318776
rect 288579 318736 288624 318764
rect 288618 318724 288624 318736
rect 288676 318724 288682 318776
rect 365806 318724 365812 318776
rect 365864 318764 365870 318776
rect 365898 318764 365904 318776
rect 365864 318736 365904 318764
rect 365864 318724 365870 318736
rect 365898 318724 365904 318736
rect 365956 318724 365962 318776
rect 371326 318724 371332 318776
rect 371384 318764 371390 318776
rect 371418 318764 371424 318776
rect 371384 318736 371424 318764
rect 371384 318724 371390 318736
rect 371418 318724 371424 318736
rect 371476 318724 371482 318776
rect 386690 318764 386696 318776
rect 386651 318736 386696 318764
rect 386690 318724 386696 318736
rect 386748 318724 386754 318776
rect 382458 317540 382464 317552
rect 382419 317512 382464 317540
rect 382458 317500 382464 317512
rect 382516 317500 382522 317552
rect 249978 317472 249984 317484
rect 249939 317444 249984 317472
rect 249978 317432 249984 317444
rect 250036 317432 250042 317484
rect 292758 317472 292764 317484
rect 292719 317444 292764 317472
rect 292758 317432 292764 317444
rect 292816 317432 292822 317484
rect 334434 317432 334440 317484
rect 334492 317472 334498 317484
rect 334526 317472 334532 317484
rect 334492 317444 334532 317472
rect 334492 317432 334498 317444
rect 334526 317432 334532 317444
rect 334584 317432 334590 317484
rect 356514 317472 356520 317484
rect 356475 317444 356520 317472
rect 356514 317432 356520 317444
rect 356572 317432 356578 317484
rect 357526 317472 357532 317484
rect 357487 317444 357532 317472
rect 357526 317432 357532 317444
rect 357584 317432 357590 317484
rect 255406 317364 255412 317416
rect 255464 317364 255470 317416
rect 281626 317404 281632 317416
rect 281587 317376 281632 317404
rect 281626 317364 281632 317376
rect 281684 317364 281690 317416
rect 283006 317404 283012 317416
rect 282967 317376 283012 317404
rect 283006 317364 283012 317376
rect 283064 317364 283070 317416
rect 327258 317364 327264 317416
rect 327316 317364 327322 317416
rect 332686 317364 332692 317416
rect 332744 317404 332750 317416
rect 332870 317404 332876 317416
rect 332744 317376 332876 317404
rect 332744 317364 332750 317376
rect 332870 317364 332876 317376
rect 332928 317364 332934 317416
rect 365806 317364 365812 317416
rect 365864 317404 365870 317416
rect 365898 317404 365904 317416
rect 365864 317376 365904 317404
rect 365864 317364 365870 317376
rect 365898 317364 365904 317376
rect 365956 317364 365962 317416
rect 371326 317404 371332 317416
rect 371287 317376 371332 317404
rect 371326 317364 371332 317376
rect 371384 317364 371390 317416
rect 376938 317404 376944 317416
rect 376899 317376 376944 317404
rect 376938 317364 376944 317376
rect 376996 317364 377002 317416
rect 381078 317364 381084 317416
rect 381136 317404 381142 317416
rect 381354 317404 381360 317416
rect 381136 317376 381360 317404
rect 381136 317364 381142 317376
rect 381354 317364 381360 317376
rect 381412 317364 381418 317416
rect 382458 317404 382464 317416
rect 382419 317376 382464 317404
rect 382458 317364 382464 317376
rect 382516 317364 382522 317416
rect 480346 317404 480352 317416
rect 480307 317376 480352 317404
rect 480346 317364 480352 317376
rect 480404 317364 480410 317416
rect 255424 317336 255452 317364
rect 255682 317336 255688 317348
rect 255424 317308 255688 317336
rect 255682 317296 255688 317308
rect 255740 317296 255746 317348
rect 327276 317280 327304 317364
rect 327258 317228 327264 317280
rect 327316 317228 327322 317280
rect 451550 316072 451556 316124
rect 451608 316112 451614 316124
rect 451734 316112 451740 316124
rect 451608 316084 451740 316112
rect 451608 316072 451614 316084
rect 451734 316072 451740 316084
rect 451792 316072 451798 316124
rect 294138 316004 294144 316056
rect 294196 316044 294202 316056
rect 294322 316044 294328 316056
rect 294196 316016 294328 316044
rect 294196 316004 294202 316016
rect 294322 316004 294328 316016
rect 294380 316004 294386 316056
rect 321462 316004 321468 316056
rect 321520 316044 321526 316056
rect 321738 316044 321744 316056
rect 321520 316016 321744 316044
rect 321520 316004 321526 316016
rect 321738 316004 321744 316016
rect 321796 316004 321802 316056
rect 352098 316004 352104 316056
rect 352156 316044 352162 316056
rect 352282 316044 352288 316056
rect 352156 316016 352288 316044
rect 352156 316004 352162 316016
rect 352282 316004 352288 316016
rect 352340 316004 352346 316056
rect 255501 315979 255559 315985
rect 255501 315945 255513 315979
rect 255547 315976 255559 315979
rect 255682 315976 255688 315988
rect 255547 315948 255688 315976
rect 255547 315945 255559 315948
rect 255501 315939 255559 315945
rect 255682 315936 255688 315948
rect 255740 315936 255746 315988
rect 400490 315976 400496 315988
rect 400451 315948 400496 315976
rect 400490 315936 400496 315948
rect 400548 315936 400554 315988
rect 408770 315976 408776 315988
rect 408731 315948 408776 315976
rect 408770 315936 408776 315948
rect 408828 315936 408834 315988
rect 451550 315976 451556 315988
rect 451511 315948 451556 315976
rect 451550 315936 451556 315948
rect 451608 315936 451614 315988
rect 232317 314687 232375 314693
rect 232317 314653 232329 314687
rect 232363 314684 232375 314687
rect 232406 314684 232412 314696
rect 232363 314656 232412 314684
rect 232363 314653 232375 314656
rect 232317 314647 232375 314653
rect 232406 314644 232412 314656
rect 232464 314644 232470 314696
rect 232314 313256 232320 313268
rect 232275 313228 232320 313256
rect 232314 313216 232320 313228
rect 232372 313216 232378 313268
rect 249886 312536 249892 312588
rect 249944 312576 249950 312588
rect 250070 312576 250076 312588
rect 249944 312548 250076 312576
rect 249944 312536 249950 312548
rect 250070 312536 250076 312548
rect 250128 312536 250134 312588
rect 277578 311964 277584 311976
rect 277539 311936 277584 311964
rect 277578 311924 277584 311936
rect 277636 311924 277642 311976
rect 294138 311924 294144 311976
rect 294196 311924 294202 311976
rect 294156 311840 294184 311924
rect 397546 311856 397552 311908
rect 397604 311896 397610 311908
rect 397914 311896 397920 311908
rect 397604 311868 397920 311896
rect 397604 311856 397610 311868
rect 397914 311856 397920 311868
rect 397972 311856 397978 311908
rect 433426 311856 433432 311908
rect 433484 311896 433490 311908
rect 433794 311896 433800 311908
rect 433484 311868 433800 311896
rect 433484 311856 433490 311868
rect 433794 311856 433800 311868
rect 433852 311856 433858 311908
rect 294138 311788 294144 311840
rect 294196 311788 294202 311840
rect 318886 311788 318892 311840
rect 318944 311828 318950 311840
rect 319070 311828 319076 311840
rect 318944 311800 319076 311828
rect 318944 311788 318950 311800
rect 319070 311788 319076 311800
rect 319128 311788 319134 311840
rect 346578 311828 346584 311840
rect 346539 311800 346584 311828
rect 346578 311788 346584 311800
rect 346636 311788 346642 311840
rect 416774 311788 416780 311840
rect 416832 311828 416838 311840
rect 416958 311828 416964 311840
rect 416832 311800 416964 311828
rect 416832 311788 416838 311800
rect 416958 311788 416964 311800
rect 417016 311788 417022 311840
rect 422294 311788 422300 311840
rect 422352 311828 422358 311840
rect 422478 311828 422484 311840
rect 422352 311800 422484 311828
rect 422352 311788 422358 311800
rect 422478 311788 422484 311800
rect 422536 311788 422542 311840
rect 427814 311788 427820 311840
rect 427872 311828 427878 311840
rect 427998 311828 428004 311840
rect 427872 311800 428004 311828
rect 427872 311788 427878 311800
rect 427998 311788 428004 311800
rect 428056 311788 428062 311840
rect 466454 311788 466460 311840
rect 466512 311828 466518 311840
rect 466638 311828 466644 311840
rect 466512 311800 466644 311828
rect 466512 311788 466518 311800
rect 466638 311788 466644 311800
rect 466696 311788 466702 311840
rect 471974 311788 471980 311840
rect 472032 311828 472038 311840
rect 472158 311828 472164 311840
rect 472032 311800 472164 311828
rect 472032 311788 472038 311800
rect 472158 311788 472164 311800
rect 472216 311788 472222 311840
rect 321462 311176 321468 311228
rect 321520 311216 321526 311228
rect 321738 311216 321744 311228
rect 321520 311188 321744 311216
rect 321520 311176 321526 311188
rect 321738 311176 321744 311188
rect 321796 311176 321802 311228
rect 392026 310904 392032 310956
rect 392084 310944 392090 310956
rect 392486 310944 392492 310956
rect 392084 310916 392492 310944
rect 392084 310904 392090 310916
rect 392486 310904 392492 310916
rect 392544 310904 392550 310956
rect 342622 309244 342628 309256
rect 342456 309216 342628 309244
rect 342456 309188 342484 309216
rect 342622 309204 342628 309216
rect 342680 309204 342686 309256
rect 252554 309136 252560 309188
rect 252612 309176 252618 309188
rect 252738 309176 252744 309188
rect 252612 309148 252744 309176
rect 252612 309136 252618 309148
rect 252738 309136 252744 309148
rect 252796 309136 252802 309188
rect 267090 309176 267096 309188
rect 267051 309148 267096 309176
rect 267090 309136 267096 309148
rect 267148 309136 267154 309188
rect 288618 309176 288624 309188
rect 288579 309148 288624 309176
rect 288618 309136 288624 309148
rect 288676 309136 288682 309188
rect 305178 309136 305184 309188
rect 305236 309176 305242 309188
rect 305270 309176 305276 309188
rect 305236 309148 305276 309176
rect 305236 309136 305242 309148
rect 305270 309136 305276 309148
rect 305328 309136 305334 309188
rect 336826 309136 336832 309188
rect 336884 309176 336890 309188
rect 336918 309176 336924 309188
rect 336884 309148 336924 309176
rect 336884 309136 336890 309148
rect 336918 309136 336924 309148
rect 336976 309136 336982 309188
rect 342438 309136 342444 309188
rect 342496 309136 342502 309188
rect 346578 309176 346584 309188
rect 346539 309148 346584 309176
rect 346578 309136 346584 309148
rect 346636 309136 346642 309188
rect 353478 309136 353484 309188
rect 353536 309176 353542 309188
rect 353570 309176 353576 309188
rect 353536 309148 353576 309176
rect 353536 309136 353542 309148
rect 353570 309136 353576 309148
rect 353628 309136 353634 309188
rect 364518 309136 364524 309188
rect 364576 309176 364582 309188
rect 364610 309176 364616 309188
rect 364576 309148 364616 309176
rect 364576 309136 364582 309148
rect 364610 309136 364616 309148
rect 364668 309136 364674 309188
rect 367370 309136 367376 309188
rect 367428 309176 367434 309188
rect 367462 309176 367468 309188
rect 367428 309148 367468 309176
rect 367428 309136 367434 309148
rect 367462 309136 367468 309148
rect 367520 309136 367526 309188
rect 386690 309176 386696 309188
rect 386651 309148 386696 309176
rect 386690 309136 386696 309148
rect 386748 309136 386754 309188
rect 270678 309108 270684 309120
rect 270639 309080 270684 309108
rect 270678 309068 270684 309080
rect 270736 309068 270742 309120
rect 309318 309108 309324 309120
rect 309279 309080 309324 309108
rect 309318 309068 309324 309080
rect 309376 309068 309382 309120
rect 318981 309111 319039 309117
rect 318981 309077 318993 309111
rect 319027 309108 319039 309111
rect 319070 309108 319076 309120
rect 319027 309080 319076 309108
rect 319027 309077 319039 309080
rect 318981 309071 319039 309077
rect 319070 309068 319076 309080
rect 319128 309068 319134 309120
rect 371326 309108 371332 309120
rect 371287 309080 371332 309108
rect 371326 309068 371332 309080
rect 371384 309068 371390 309120
rect 416869 309111 416927 309117
rect 416869 309077 416881 309111
rect 416915 309108 416927 309111
rect 416958 309108 416964 309120
rect 416915 309080 416964 309108
rect 416915 309077 416927 309080
rect 416869 309071 416927 309077
rect 416958 309068 416964 309080
rect 417016 309068 417022 309120
rect 422478 309108 422484 309120
rect 422439 309080 422484 309108
rect 422478 309068 422484 309080
rect 422536 309068 422542 309120
rect 427998 309108 428004 309120
rect 427959 309080 428004 309108
rect 427998 309068 428004 309080
rect 428056 309068 428062 309120
rect 433426 309108 433432 309120
rect 433387 309080 433432 309108
rect 433426 309068 433432 309080
rect 433484 309068 433490 309120
rect 466549 309111 466607 309117
rect 466549 309077 466561 309111
rect 466595 309108 466607 309111
rect 466638 309108 466644 309120
rect 466595 309080 466644 309108
rect 466595 309077 466607 309080
rect 466549 309071 466607 309077
rect 466638 309068 466644 309080
rect 466696 309068 466702 309120
rect 472069 309111 472127 309117
rect 472069 309077 472081 309111
rect 472115 309108 472127 309111
rect 472158 309108 472164 309120
rect 472115 309080 472164 309108
rect 472115 309077 472127 309080
rect 472069 309071 472127 309077
rect 472158 309068 472164 309080
rect 472216 309068 472222 309120
rect 277486 309000 277492 309052
rect 277544 309040 277550 309052
rect 277581 309043 277639 309049
rect 277581 309040 277593 309043
rect 277544 309012 277593 309040
rect 277544 309000 277550 309012
rect 277581 309009 277593 309012
rect 277627 309009 277639 309043
rect 342438 309040 342444 309052
rect 342399 309012 342444 309040
rect 277581 309003 277639 309009
rect 342438 309000 342444 309012
rect 342496 309000 342502 309052
rect 2774 308796 2780 308848
rect 2832 308836 2838 308848
rect 4982 308836 4988 308848
rect 2832 308808 4988 308836
rect 2832 308796 2838 308808
rect 4982 308796 4988 308808
rect 5040 308796 5046 308848
rect 287146 307844 287152 307896
rect 287204 307884 287210 307896
rect 287330 307884 287336 307896
rect 287204 307856 287336 307884
rect 287204 307844 287210 307856
rect 287330 307844 287336 307856
rect 287388 307844 287394 307896
rect 261018 307776 261024 307828
rect 261076 307816 261082 307828
rect 261110 307816 261116 307828
rect 261076 307788 261116 307816
rect 261076 307776 261082 307788
rect 261110 307776 261116 307788
rect 261168 307776 261174 307828
rect 267090 307816 267096 307828
rect 267051 307788 267096 307816
rect 267090 307776 267096 307788
rect 267148 307776 267154 307828
rect 281626 307816 281632 307828
rect 281587 307788 281632 307816
rect 281626 307776 281632 307788
rect 281684 307776 281690 307828
rect 283006 307816 283012 307828
rect 282967 307788 283012 307816
rect 283006 307776 283012 307788
rect 283064 307776 283070 307828
rect 376938 307816 376944 307828
rect 376899 307788 376944 307816
rect 376938 307776 376944 307788
rect 376996 307776 377002 307828
rect 382458 307816 382464 307828
rect 382419 307788 382464 307816
rect 382458 307776 382464 307788
rect 382516 307776 382522 307828
rect 480346 307816 480352 307828
rect 480307 307788 480352 307816
rect 480346 307776 480352 307788
rect 480404 307776 480410 307828
rect 242989 307751 243047 307757
rect 242989 307717 243001 307751
rect 243035 307748 243047 307751
rect 243078 307748 243084 307760
rect 243035 307720 243084 307748
rect 243035 307717 243047 307720
rect 242989 307711 243047 307717
rect 243078 307708 243084 307720
rect 243136 307708 243142 307760
rect 277578 307748 277584 307760
rect 277539 307720 277584 307748
rect 277578 307708 277584 307720
rect 277636 307708 277642 307760
rect 287241 307751 287299 307757
rect 287241 307717 287253 307751
rect 287287 307748 287299 307751
rect 287330 307748 287336 307760
rect 287287 307720 287336 307748
rect 287287 307717 287299 307720
rect 287241 307711 287299 307717
rect 287330 307708 287336 307720
rect 287388 307708 287394 307760
rect 295518 307748 295524 307760
rect 295479 307720 295524 307748
rect 295518 307708 295524 307720
rect 295576 307708 295582 307760
rect 364518 307748 364524 307760
rect 364479 307720 364524 307748
rect 364518 307708 364524 307720
rect 364576 307708 364582 307760
rect 332686 306416 332692 306468
rect 332744 306456 332750 306468
rect 332870 306456 332876 306468
rect 332744 306428 332876 306456
rect 332744 306416 332750 306428
rect 332870 306416 332876 306428
rect 332928 306416 332934 306468
rect 352098 306348 352104 306400
rect 352156 306388 352162 306400
rect 352282 306388 352288 306400
rect 352156 306360 352288 306388
rect 352156 306348 352162 306360
rect 352282 306348 352288 306360
rect 352340 306348 352346 306400
rect 357526 306348 357532 306400
rect 357584 306388 357590 306400
rect 357710 306388 357716 306400
rect 357584 306360 357716 306388
rect 357584 306348 357590 306360
rect 357710 306348 357716 306360
rect 357768 306348 357774 306400
rect 236362 304920 236368 304972
rect 236420 304960 236426 304972
rect 236546 304960 236552 304972
rect 236420 304932 236552 304960
rect 236420 304920 236426 304932
rect 236546 304920 236552 304932
rect 236604 304920 236610 304972
rect 281626 302268 281632 302320
rect 281684 302268 281690 302320
rect 283006 302268 283012 302320
rect 283064 302268 283070 302320
rect 298278 302268 298284 302320
rect 298336 302268 298342 302320
rect 233326 302200 233332 302252
rect 233384 302240 233390 302252
rect 233510 302240 233516 302252
rect 233384 302212 233516 302240
rect 233384 302200 233390 302212
rect 233510 302200 233516 302212
rect 233568 302200 233574 302252
rect 281644 302104 281672 302268
rect 281810 302104 281816 302116
rect 281644 302076 281816 302104
rect 281810 302064 281816 302076
rect 281868 302064 281874 302116
rect 283024 302104 283052 302268
rect 283098 302104 283104 302116
rect 283024 302076 283104 302104
rect 283098 302064 283104 302076
rect 283156 302064 283162 302116
rect 298296 302104 298324 302268
rect 298370 302104 298376 302116
rect 298296 302076 298376 302104
rect 298370 302064 298376 302076
rect 298428 302064 298434 302116
rect 408770 302104 408776 302116
rect 408731 302076 408776 302104
rect 408770 302064 408776 302076
rect 408828 302064 408834 302116
rect 451550 302104 451556 302116
rect 451511 302076 451556 302104
rect 451550 302064 451556 302076
rect 451608 302064 451614 302116
rect 422478 299928 422484 299940
rect 422439 299900 422484 299928
rect 422478 299888 422484 299900
rect 422536 299888 422542 299940
rect 342441 299591 342499 299597
rect 342441 299557 342453 299591
rect 342487 299588 342499 299591
rect 342530 299588 342536 299600
rect 342487 299560 342536 299588
rect 342487 299557 342499 299560
rect 342441 299551 342499 299557
rect 342530 299548 342536 299560
rect 342588 299548 342594 299600
rect 347958 299548 347964 299600
rect 348016 299548 348022 299600
rect 353478 299548 353484 299600
rect 353536 299548 353542 299600
rect 265158 299480 265164 299532
rect 265216 299520 265222 299532
rect 265250 299520 265256 299532
rect 265216 299492 265256 299520
rect 265216 299480 265222 299492
rect 265250 299480 265256 299492
rect 265308 299480 265314 299532
rect 270681 299523 270739 299529
rect 270681 299489 270693 299523
rect 270727 299520 270739 299523
rect 270770 299520 270776 299532
rect 270727 299492 270776 299520
rect 270727 299489 270739 299492
rect 270681 299483 270739 299489
rect 270770 299480 270776 299492
rect 270828 299480 270834 299532
rect 309321 299523 309379 299529
rect 309321 299489 309333 299523
rect 309367 299520 309379 299523
rect 309410 299520 309416 299532
rect 309367 299492 309416 299520
rect 309367 299489 309379 299492
rect 309321 299483 309379 299489
rect 309410 299480 309416 299492
rect 309468 299480 309474 299532
rect 318978 299520 318984 299532
rect 318939 299492 318984 299520
rect 318978 299480 318984 299492
rect 319036 299480 319042 299532
rect 241790 299452 241796 299464
rect 241751 299424 241796 299452
rect 241790 299412 241796 299424
rect 241848 299412 241854 299464
rect 249978 299452 249984 299464
rect 249939 299424 249984 299452
rect 249978 299412 249984 299424
rect 250036 299412 250042 299464
rect 281629 299455 281687 299461
rect 281629 299421 281641 299455
rect 281675 299452 281687 299455
rect 281810 299452 281816 299464
rect 281675 299424 281816 299452
rect 281675 299421 281687 299424
rect 281629 299415 281687 299421
rect 281810 299412 281816 299424
rect 281868 299412 281874 299464
rect 283098 299452 283104 299464
rect 283059 299424 283104 299452
rect 283098 299412 283104 299424
rect 283156 299412 283162 299464
rect 288618 299452 288624 299464
rect 288579 299424 288624 299452
rect 288618 299412 288624 299424
rect 288676 299412 288682 299464
rect 305178 299452 305184 299464
rect 305139 299424 305184 299452
rect 305178 299412 305184 299424
rect 305236 299412 305242 299464
rect 310698 299452 310704 299464
rect 310659 299424 310704 299452
rect 310698 299412 310704 299424
rect 310756 299412 310762 299464
rect 331398 299412 331404 299464
rect 331456 299452 331462 299464
rect 331490 299452 331496 299464
rect 331456 299424 331496 299452
rect 331456 299412 331462 299424
rect 331490 299412 331496 299424
rect 331548 299412 331554 299464
rect 346578 299452 346584 299464
rect 346539 299424 346584 299452
rect 346578 299412 346584 299424
rect 346636 299412 346642 299464
rect 347976 299396 348004 299548
rect 353496 299396 353524 299548
rect 416866 299520 416872 299532
rect 416827 299492 416872 299520
rect 416866 299480 416872 299492
rect 416924 299480 416930 299532
rect 427998 299520 428004 299532
rect 427959 299492 428004 299520
rect 427998 299480 428004 299492
rect 428056 299480 428062 299532
rect 433429 299523 433487 299529
rect 433429 299489 433441 299523
rect 433475 299520 433487 299523
rect 433702 299520 433708 299532
rect 433475 299492 433708 299520
rect 433475 299489 433487 299492
rect 433429 299483 433487 299489
rect 433702 299480 433708 299492
rect 433760 299480 433766 299532
rect 466546 299520 466552 299532
rect 466507 299492 466552 299520
rect 466546 299480 466552 299492
rect 466604 299480 466610 299532
rect 472066 299520 472072 299532
rect 472027 299492 472072 299520
rect 472066 299480 472072 299492
rect 472124 299480 472130 299532
rect 370038 299412 370044 299464
rect 370096 299452 370102 299464
rect 370130 299452 370136 299464
rect 370096 299424 370136 299452
rect 370096 299412 370102 299424
rect 370130 299412 370136 299424
rect 370188 299412 370194 299464
rect 376938 299452 376944 299464
rect 376899 299424 376944 299452
rect 376938 299412 376944 299424
rect 376996 299412 377002 299464
rect 400490 299452 400496 299464
rect 400451 299424 400496 299452
rect 400490 299412 400496 299424
rect 400548 299412 400554 299464
rect 530578 299412 530584 299464
rect 530636 299452 530642 299464
rect 579706 299452 579712 299464
rect 530636 299424 579712 299452
rect 530636 299412 530642 299424
rect 579706 299412 579712 299424
rect 579764 299412 579770 299464
rect 347958 299344 347964 299396
rect 348016 299344 348022 299396
rect 353478 299344 353484 299396
rect 353536 299344 353542 299396
rect 242986 298228 242992 298240
rect 242947 298200 242992 298228
rect 242986 298188 242992 298200
rect 243044 298188 243050 298240
rect 277578 298228 277584 298240
rect 277539 298200 277584 298228
rect 277578 298188 277584 298200
rect 277636 298188 277642 298240
rect 295521 298231 295579 298237
rect 295521 298197 295533 298231
rect 295567 298228 295579 298231
rect 295567 298200 295656 298228
rect 295567 298197 295579 298200
rect 295521 298191 295579 298197
rect 255498 298160 255504 298172
rect 255459 298132 255504 298160
rect 255498 298120 255504 298132
rect 255556 298120 255562 298172
rect 261018 298120 261024 298172
rect 261076 298160 261082 298172
rect 261202 298160 261208 298172
rect 261076 298132 261208 298160
rect 261076 298120 261082 298132
rect 261202 298120 261208 298132
rect 261260 298120 261266 298172
rect 287238 298160 287244 298172
rect 287199 298132 287244 298160
rect 287238 298120 287244 298132
rect 287296 298120 287302 298172
rect 242986 298092 242992 298104
rect 242947 298064 242992 298092
rect 242986 298052 242992 298064
rect 243044 298052 243050 298104
rect 265161 298095 265219 298101
rect 265161 298061 265173 298095
rect 265207 298092 265219 298095
rect 265250 298092 265256 298104
rect 265207 298064 265256 298092
rect 265207 298061 265219 298064
rect 265161 298055 265219 298061
rect 265250 298052 265256 298064
rect 265308 298052 265314 298104
rect 267001 298095 267059 298101
rect 267001 298061 267013 298095
rect 267047 298092 267059 298095
rect 267090 298092 267096 298104
rect 267047 298064 267096 298092
rect 267047 298061 267059 298064
rect 267001 298055 267059 298061
rect 267090 298052 267096 298064
rect 267148 298052 267154 298104
rect 270770 298052 270776 298104
rect 270828 298092 270834 298104
rect 270862 298092 270868 298104
rect 270828 298064 270868 298092
rect 270828 298052 270834 298064
rect 270862 298052 270868 298064
rect 270920 298052 270926 298104
rect 277578 298092 277584 298104
rect 277539 298064 277584 298092
rect 277578 298052 277584 298064
rect 277636 298052 277642 298104
rect 292669 298095 292727 298101
rect 292669 298061 292681 298095
rect 292715 298092 292727 298095
rect 292758 298092 292764 298104
rect 292715 298064 292764 298092
rect 292715 298061 292727 298064
rect 292669 298055 292727 298061
rect 292758 298052 292764 298064
rect 292816 298052 292822 298104
rect 295628 298101 295656 298200
rect 334250 298160 334256 298172
rect 334211 298132 334256 298160
rect 334250 298120 334256 298132
rect 334308 298120 334314 298172
rect 364521 298163 364579 298169
rect 364521 298129 364533 298163
rect 364567 298160 364579 298163
rect 364610 298160 364616 298172
rect 364567 298132 364616 298160
rect 364567 298129 364579 298132
rect 364521 298123 364579 298129
rect 364610 298120 364616 298132
rect 364668 298120 364674 298172
rect 295613 298095 295671 298101
rect 295613 298061 295625 298095
rect 295659 298061 295671 298095
rect 347958 298092 347964 298104
rect 347919 298064 347964 298092
rect 295613 298055 295671 298061
rect 347958 298052 347964 298064
rect 348016 298052 348022 298104
rect 352098 298092 352104 298104
rect 352059 298064 352104 298092
rect 352098 298052 352104 298064
rect 352156 298052 352162 298104
rect 353478 298052 353484 298104
rect 353536 298092 353542 298104
rect 353570 298092 353576 298104
rect 353536 298064 353576 298092
rect 353536 298052 353542 298064
rect 353570 298052 353576 298064
rect 353628 298052 353634 298104
rect 370038 298092 370044 298104
rect 369999 298064 370044 298092
rect 370038 298052 370044 298064
rect 370096 298052 370102 298104
rect 375466 298092 375472 298104
rect 375427 298064 375472 298092
rect 375466 298052 375472 298064
rect 375524 298052 375530 298104
rect 397730 298092 397736 298104
rect 397691 298064 397736 298092
rect 397730 298052 397736 298064
rect 397788 298052 397794 298104
rect 480346 298092 480352 298104
rect 480307 298064 480352 298092
rect 480346 298052 480352 298064
rect 480404 298052 480410 298104
rect 382458 297984 382464 298036
rect 382516 298024 382522 298036
rect 382550 298024 382556 298036
rect 382516 297996 382556 298024
rect 382516 297984 382522 297996
rect 382550 297984 382556 297996
rect 382608 297984 382614 298036
rect 332778 296692 332784 296744
rect 332836 296732 332842 296744
rect 332962 296732 332968 296744
rect 332836 296704 332968 296732
rect 332836 296692 332842 296704
rect 332962 296692 332968 296704
rect 333020 296692 333026 296744
rect 334250 296732 334256 296744
rect 334211 296704 334256 296732
rect 334250 296692 334256 296704
rect 334308 296692 334314 296744
rect 298370 296664 298376 296676
rect 298331 296636 298376 296664
rect 298370 296624 298376 296636
rect 298428 296624 298434 296676
rect 236270 295264 236276 295316
rect 236328 295304 236334 295316
rect 236454 295304 236460 295316
rect 236328 295276 236460 295304
rect 236328 295264 236334 295276
rect 236454 295264 236460 295276
rect 236512 295264 236518 295316
rect 3326 294924 3332 294976
rect 3384 294964 3390 294976
rect 7742 294964 7748 294976
rect 3384 294936 7748 294964
rect 3384 294924 3390 294936
rect 7742 294924 7748 294936
rect 7800 294924 7806 294976
rect 232314 294896 232320 294908
rect 232275 294868 232320 294896
rect 232314 294856 232320 294868
rect 232372 294856 232378 294908
rect 232314 293904 232320 293956
rect 232372 293944 232378 293956
rect 232406 293944 232412 293956
rect 232372 293916 232412 293944
rect 232372 293904 232378 293916
rect 232406 293904 232412 293916
rect 232464 293904 232470 293956
rect 295613 293267 295671 293273
rect 295613 293233 295625 293267
rect 295659 293264 295671 293267
rect 295702 293264 295708 293276
rect 295659 293236 295708 293264
rect 295659 293233 295671 293236
rect 295613 293227 295671 293233
rect 295702 293224 295708 293236
rect 295760 293224 295766 293276
rect 255498 292612 255504 292664
rect 255556 292612 255562 292664
rect 321738 292612 321744 292664
rect 321796 292612 321802 292664
rect 327258 292612 327264 292664
rect 327316 292612 327322 292664
rect 330018 292612 330024 292664
rect 330076 292612 330082 292664
rect 367370 292612 367376 292664
rect 367428 292612 367434 292664
rect 408770 292652 408776 292664
rect 408696 292624 408776 292652
rect 255516 292528 255544 292612
rect 321756 292528 321784 292612
rect 327276 292528 327304 292612
rect 330036 292528 330064 292612
rect 367388 292528 367416 292612
rect 392210 292584 392216 292596
rect 392136 292556 392216 292584
rect 392136 292528 392164 292556
rect 392210 292544 392216 292556
rect 392268 292544 392274 292596
rect 408696 292528 408724 292624
rect 408770 292612 408776 292624
rect 408828 292612 408834 292664
rect 451550 292652 451556 292664
rect 451476 292624 451556 292652
rect 451476 292528 451504 292624
rect 451550 292612 451556 292624
rect 451608 292612 451614 292664
rect 232406 292516 232412 292528
rect 232367 292488 232412 292516
rect 232406 292476 232412 292488
rect 232464 292476 232470 292528
rect 236454 292516 236460 292528
rect 236415 292488 236460 292516
rect 236454 292476 236460 292488
rect 236512 292476 236518 292528
rect 244458 292476 244464 292528
rect 244516 292476 244522 292528
rect 255498 292476 255504 292528
rect 255556 292476 255562 292528
rect 321738 292476 321744 292528
rect 321796 292476 321802 292528
rect 327258 292476 327264 292528
rect 327316 292476 327322 292528
rect 330018 292476 330024 292528
rect 330076 292476 330082 292528
rect 367370 292476 367376 292528
rect 367428 292476 367434 292528
rect 392118 292476 392124 292528
rect 392176 292476 392182 292528
rect 408678 292476 408684 292528
rect 408736 292476 408742 292528
rect 451458 292476 451464 292528
rect 451516 292476 451522 292528
rect 466454 292476 466460 292528
rect 466512 292516 466518 292528
rect 466638 292516 466644 292528
rect 466512 292488 466644 292516
rect 466512 292476 466518 292488
rect 466638 292476 466644 292488
rect 466696 292476 466702 292528
rect 471974 292476 471980 292528
rect 472032 292516 472038 292528
rect 472158 292516 472164 292528
rect 472032 292488 472164 292516
rect 472032 292476 472038 292488
rect 472158 292476 472164 292488
rect 472216 292476 472222 292528
rect 244476 292392 244504 292476
rect 244458 292340 244464 292392
rect 244516 292340 244522 292392
rect 364518 291360 364524 291372
rect 364479 291332 364524 291360
rect 364518 291320 364524 291332
rect 364576 291320 364582 291372
rect 241790 289864 241796 289876
rect 241751 289836 241796 289864
rect 241790 289824 241796 289836
rect 241848 289824 241854 289876
rect 249978 289864 249984 289876
rect 249939 289836 249984 289864
rect 249978 289824 249984 289836
rect 250036 289824 250042 289876
rect 281626 289864 281632 289876
rect 281587 289836 281632 289864
rect 281626 289824 281632 289836
rect 281684 289824 281690 289876
rect 283098 289864 283104 289876
rect 283059 289836 283104 289864
rect 283098 289824 283104 289836
rect 283156 289824 283162 289876
rect 288618 289864 288624 289876
rect 288579 289836 288624 289864
rect 288618 289824 288624 289836
rect 288676 289824 288682 289876
rect 305178 289864 305184 289876
rect 305139 289836 305184 289864
rect 305178 289824 305184 289836
rect 305236 289824 305242 289876
rect 309318 289824 309324 289876
rect 309376 289864 309382 289876
rect 309594 289864 309600 289876
rect 309376 289836 309600 289864
rect 309376 289824 309382 289836
rect 309594 289824 309600 289836
rect 309652 289824 309658 289876
rect 310698 289864 310704 289876
rect 310659 289836 310704 289864
rect 310698 289824 310704 289836
rect 310756 289824 310762 289876
rect 324498 289824 324504 289876
rect 324556 289864 324562 289876
rect 324682 289864 324688 289876
rect 324556 289836 324688 289864
rect 324556 289824 324562 289836
rect 324682 289824 324688 289836
rect 324740 289824 324746 289876
rect 346578 289864 346584 289876
rect 346539 289836 346584 289864
rect 346578 289824 346584 289836
rect 346636 289824 346642 289876
rect 376938 289864 376944 289876
rect 376899 289836 376944 289864
rect 376938 289824 376944 289836
rect 376996 289824 377002 289876
rect 381078 289824 381084 289876
rect 381136 289864 381142 289876
rect 381354 289864 381360 289876
rect 381136 289836 381360 289864
rect 381136 289824 381142 289836
rect 381354 289824 381360 289836
rect 381412 289824 381418 289876
rect 252738 289796 252744 289808
rect 252699 289768 252744 289796
rect 252738 289756 252744 289768
rect 252796 289756 252802 289808
rect 254118 289796 254124 289808
rect 254079 289768 254124 289796
rect 254118 289756 254124 289768
rect 254176 289756 254182 289808
rect 259638 289796 259644 289808
rect 259599 289768 259644 289796
rect 259638 289756 259644 289768
rect 259696 289756 259702 289808
rect 334250 289796 334256 289808
rect 334211 289768 334256 289796
rect 334250 289756 334256 289768
rect 334308 289756 334314 289808
rect 356422 289756 356428 289808
rect 356480 289756 356486 289808
rect 375466 289796 375472 289808
rect 375427 289768 375472 289796
rect 375466 289756 375472 289768
rect 375524 289756 375530 289808
rect 309318 289728 309324 289740
rect 309279 289700 309324 289728
rect 309318 289688 309324 289700
rect 309376 289688 309382 289740
rect 356440 289728 356468 289756
rect 356514 289728 356520 289740
rect 356440 289700 356520 289728
rect 356514 289688 356520 289700
rect 356572 289688 356578 289740
rect 265158 288436 265164 288448
rect 265119 288408 265164 288436
rect 265158 288396 265164 288408
rect 265216 288396 265222 288448
rect 292666 288436 292672 288448
rect 292627 288408 292672 288436
rect 292666 288396 292672 288408
rect 292724 288396 292730 288448
rect 347961 288439 348019 288445
rect 347961 288405 347973 288439
rect 348007 288436 348019 288439
rect 348050 288436 348056 288448
rect 348007 288408 348056 288436
rect 348007 288405 348019 288408
rect 347961 288399 348019 288405
rect 348050 288396 348056 288408
rect 348108 288396 348114 288448
rect 370038 288436 370044 288448
rect 369999 288408 370044 288436
rect 370038 288396 370044 288408
rect 370096 288396 370102 288448
rect 397730 288436 397736 288448
rect 397691 288408 397736 288436
rect 397730 288396 397736 288408
rect 397788 288396 397794 288448
rect 480346 288436 480352 288448
rect 480307 288408 480352 288436
rect 480346 288396 480352 288408
rect 480404 288396 480410 288448
rect 408678 288368 408684 288380
rect 408639 288340 408684 288368
rect 408678 288328 408684 288340
rect 408736 288328 408742 288380
rect 352098 287960 352104 287972
rect 352059 287932 352104 287960
rect 352098 287920 352104 287932
rect 352156 287920 352162 287972
rect 298373 287079 298431 287085
rect 298373 287045 298385 287079
rect 298419 287076 298431 287079
rect 298462 287076 298468 287088
rect 298419 287048 298468 287076
rect 298419 287045 298431 287048
rect 298373 287039 298431 287045
rect 298462 287036 298468 287048
rect 298520 287036 298526 287088
rect 386598 287076 386604 287088
rect 386559 287048 386604 287076
rect 386598 287036 386604 287048
rect 386656 287036 386662 287088
rect 364521 284971 364579 284977
rect 364521 284937 364533 284971
rect 364567 284968 364579 284971
rect 364610 284968 364616 284980
rect 364567 284940 364616 284968
rect 364567 284937 364579 284940
rect 364521 284931 364579 284937
rect 364610 284928 364616 284940
rect 364668 284928 364674 284980
rect 236454 284356 236460 284368
rect 236415 284328 236460 284356
rect 236454 284316 236460 284328
rect 236512 284316 236518 284368
rect 232406 282928 232412 282940
rect 232367 282900 232412 282928
rect 232406 282888 232412 282900
rect 232464 282888 232470 282940
rect 233326 282888 233332 282940
rect 233384 282928 233390 282940
rect 233510 282928 233516 282940
rect 233384 282900 233516 282928
rect 233384 282888 233390 282900
rect 233510 282888 233516 282900
rect 233568 282888 233574 282940
rect 342530 282928 342536 282940
rect 342491 282900 342536 282928
rect 342530 282888 342536 282900
rect 342588 282888 342594 282940
rect 370038 282888 370044 282940
rect 370096 282888 370102 282940
rect 381078 282888 381084 282940
rect 381136 282888 381142 282940
rect 422294 282888 422300 282940
rect 422352 282928 422358 282940
rect 422478 282928 422484 282940
rect 422352 282900 422484 282928
rect 422352 282888 422358 282900
rect 422478 282888 422484 282900
rect 422536 282888 422542 282940
rect 427814 282888 427820 282940
rect 427872 282928 427878 282940
rect 427998 282928 428004 282940
rect 427872 282900 428004 282928
rect 427872 282888 427878 282900
rect 427998 282888 428004 282900
rect 428056 282888 428062 282940
rect 334253 282795 334311 282801
rect 334253 282761 334265 282795
rect 334299 282792 334311 282795
rect 334434 282792 334440 282804
rect 334299 282764 334440 282792
rect 334299 282761 334311 282764
rect 334253 282755 334311 282761
rect 334434 282752 334440 282764
rect 334492 282752 334498 282804
rect 370056 282792 370084 282888
rect 375466 282820 375472 282872
rect 375524 282820 375530 282872
rect 370130 282792 370136 282804
rect 370056 282764 370136 282792
rect 370130 282752 370136 282764
rect 370188 282752 370194 282804
rect 375484 282792 375512 282820
rect 375650 282792 375656 282804
rect 375484 282764 375656 282792
rect 375650 282752 375656 282764
rect 375708 282752 375714 282804
rect 381096 282792 381124 282888
rect 400490 282820 400496 282872
rect 400548 282820 400554 282872
rect 381170 282792 381176 282804
rect 381096 282764 381176 282792
rect 381170 282752 381176 282764
rect 381228 282752 381234 282804
rect 400508 282736 400536 282820
rect 400490 282684 400496 282736
rect 400548 282684 400554 282736
rect 342530 280276 342536 280288
rect 342491 280248 342536 280276
rect 342530 280236 342536 280248
rect 342588 280236 342594 280288
rect 242989 280211 243047 280217
rect 242989 280177 243001 280211
rect 243035 280208 243047 280211
rect 243170 280208 243176 280220
rect 243035 280180 243176 280208
rect 243035 280177 243047 280180
rect 242989 280171 243047 280177
rect 243170 280168 243176 280180
rect 243228 280168 243234 280220
rect 252738 280208 252744 280220
rect 252699 280180 252744 280208
rect 252738 280168 252744 280180
rect 252796 280168 252802 280220
rect 265066 280168 265072 280220
rect 265124 280208 265130 280220
rect 265250 280208 265256 280220
rect 265124 280180 265256 280208
rect 265124 280168 265130 280180
rect 265250 280168 265256 280180
rect 265308 280168 265314 280220
rect 266998 280208 267004 280220
rect 266959 280180 267004 280208
rect 266998 280168 267004 280180
rect 267056 280168 267062 280220
rect 277581 280211 277639 280217
rect 277581 280177 277593 280211
rect 277627 280208 277639 280211
rect 277670 280208 277676 280220
rect 277627 280180 277676 280208
rect 277627 280177 277639 280180
rect 277581 280171 277639 280177
rect 277670 280168 277676 280180
rect 277728 280168 277734 280220
rect 281718 280168 281724 280220
rect 281776 280208 281782 280220
rect 281902 280208 281908 280220
rect 281776 280180 281908 280208
rect 281776 280168 281782 280180
rect 281902 280168 281908 280180
rect 281960 280168 281966 280220
rect 292666 280168 292672 280220
rect 292724 280208 292730 280220
rect 292758 280208 292764 280220
rect 292724 280180 292764 280208
rect 292724 280168 292730 280180
rect 292758 280168 292764 280180
rect 292816 280168 292822 280220
rect 309321 280211 309379 280217
rect 309321 280177 309333 280211
rect 309367 280208 309379 280211
rect 309410 280208 309416 280220
rect 309367 280180 309416 280208
rect 309367 280177 309379 280180
rect 309321 280171 309379 280177
rect 309410 280168 309416 280180
rect 309468 280168 309474 280220
rect 324406 280168 324412 280220
rect 324464 280208 324470 280220
rect 324682 280208 324688 280220
rect 324464 280180 324688 280208
rect 324464 280168 324470 280180
rect 324682 280168 324688 280180
rect 324740 280168 324746 280220
rect 397454 280168 397460 280220
rect 397512 280168 397518 280220
rect 3142 280100 3148 280152
rect 3200 280140 3206 280152
rect 6270 280140 6276 280152
rect 3200 280112 6276 280140
rect 3200 280100 3206 280112
rect 6270 280100 6276 280112
rect 6328 280100 6334 280152
rect 241790 280140 241796 280152
rect 241751 280112 241796 280140
rect 241790 280100 241796 280112
rect 241848 280100 241854 280152
rect 270586 280100 270592 280152
rect 270644 280140 270650 280152
rect 270862 280140 270868 280152
rect 270644 280112 270868 280140
rect 270644 280100 270650 280112
rect 270862 280100 270868 280112
rect 270920 280100 270926 280152
rect 288618 280140 288624 280152
rect 288579 280112 288624 280140
rect 288618 280100 288624 280112
rect 288676 280100 288682 280152
rect 295426 280100 295432 280152
rect 295484 280140 295490 280152
rect 295702 280140 295708 280152
rect 295484 280112 295708 280140
rect 295484 280100 295490 280112
rect 295702 280100 295708 280112
rect 295760 280100 295766 280152
rect 298462 280140 298468 280152
rect 298296 280112 298468 280140
rect 298296 280084 298324 280112
rect 298462 280100 298468 280112
rect 298520 280100 298526 280152
rect 305178 280140 305184 280152
rect 305139 280112 305184 280140
rect 305178 280100 305184 280112
rect 305236 280100 305242 280152
rect 310698 280140 310704 280152
rect 310659 280112 310704 280140
rect 310698 280100 310704 280112
rect 310756 280100 310762 280152
rect 318978 280100 318984 280152
rect 319036 280140 319042 280152
rect 319070 280140 319076 280152
rect 319036 280112 319076 280140
rect 319036 280100 319042 280112
rect 319070 280100 319076 280112
rect 319128 280100 319134 280152
rect 321738 280140 321744 280152
rect 321699 280112 321744 280140
rect 321738 280100 321744 280112
rect 321796 280100 321802 280152
rect 327258 280140 327264 280152
rect 327219 280112 327264 280140
rect 327258 280100 327264 280112
rect 327316 280100 327322 280152
rect 331398 280100 331404 280152
rect 331456 280140 331462 280152
rect 331490 280140 331496 280152
rect 331456 280112 331496 280140
rect 331456 280100 331462 280112
rect 331490 280100 331496 280112
rect 331548 280100 331554 280152
rect 334345 280143 334403 280149
rect 334345 280109 334357 280143
rect 334391 280140 334403 280143
rect 334434 280140 334440 280152
rect 334391 280112 334440 280140
rect 334391 280109 334403 280112
rect 334345 280103 334403 280109
rect 334434 280100 334440 280112
rect 334492 280100 334498 280152
rect 346578 280140 346584 280152
rect 346539 280112 346584 280140
rect 346578 280100 346584 280112
rect 346636 280100 346642 280152
rect 348050 280100 348056 280152
rect 348108 280140 348114 280152
rect 348142 280140 348148 280152
rect 348108 280112 348148 280140
rect 348108 280100 348114 280112
rect 348142 280100 348148 280112
rect 348200 280100 348206 280152
rect 352098 280100 352104 280152
rect 352156 280140 352162 280152
rect 352282 280140 352288 280152
rect 352156 280112 352288 280140
rect 352156 280100 352162 280112
rect 352282 280100 352288 280112
rect 352340 280100 352346 280152
rect 353478 280100 353484 280152
rect 353536 280140 353542 280152
rect 353570 280140 353576 280152
rect 353536 280112 353576 280140
rect 353536 280100 353542 280112
rect 353570 280100 353576 280112
rect 353628 280100 353634 280152
rect 358998 280100 359004 280152
rect 359056 280140 359062 280152
rect 359090 280140 359096 280152
rect 359056 280112 359096 280140
rect 359056 280100 359062 280112
rect 359090 280100 359096 280112
rect 359148 280100 359154 280152
rect 364518 280100 364524 280152
rect 364576 280140 364582 280152
rect 364610 280140 364616 280152
rect 364576 280112 364616 280140
rect 364576 280100 364582 280112
rect 364610 280100 364616 280112
rect 364668 280100 364674 280152
rect 365898 280100 365904 280152
rect 365956 280140 365962 280152
rect 365990 280140 365996 280152
rect 365956 280112 365996 280140
rect 365956 280100 365962 280112
rect 365990 280100 365996 280112
rect 366048 280100 366054 280152
rect 369762 280100 369768 280152
rect 369820 280140 369826 280152
rect 370130 280140 370136 280152
rect 369820 280112 370136 280140
rect 369820 280100 369826 280112
rect 370130 280100 370136 280112
rect 370188 280100 370194 280152
rect 371418 280100 371424 280152
rect 371476 280140 371482 280152
rect 371510 280140 371516 280152
rect 371476 280112 371516 280140
rect 371476 280100 371482 280112
rect 371510 280100 371516 280112
rect 371568 280100 371574 280152
rect 375190 280100 375196 280152
rect 375248 280140 375254 280152
rect 375650 280140 375656 280152
rect 375248 280112 375656 280140
rect 375248 280100 375254 280112
rect 375650 280100 375656 280112
rect 375708 280100 375714 280152
rect 382458 280140 382464 280152
rect 382419 280112 382464 280140
rect 382458 280100 382464 280112
rect 382516 280100 382522 280152
rect 397472 280084 397500 280168
rect 416866 280140 416872 280152
rect 416827 280112 416872 280140
rect 416866 280100 416872 280112
rect 416924 280100 416930 280152
rect 433610 280140 433616 280152
rect 433571 280112 433616 280140
rect 433610 280100 433616 280112
rect 433668 280100 433674 280152
rect 466546 280140 466552 280152
rect 466507 280112 466552 280140
rect 466546 280100 466552 280112
rect 466604 280100 466610 280152
rect 472066 280140 472072 280152
rect 472027 280112 472072 280140
rect 472066 280100 472072 280112
rect 472124 280100 472130 280152
rect 298278 280032 298284 280084
rect 298336 280032 298342 280084
rect 381081 280075 381139 280081
rect 381081 280041 381093 280075
rect 381127 280072 381139 280075
rect 381170 280072 381176 280084
rect 381127 280044 381176 280072
rect 381127 280041 381139 280044
rect 381081 280035 381139 280041
rect 381170 280032 381176 280044
rect 381228 280032 381234 280084
rect 397454 280032 397460 280084
rect 397512 280032 397518 280084
rect 357618 278740 357624 278792
rect 357676 278780 357682 278792
rect 357802 278780 357808 278792
rect 357676 278752 357808 278780
rect 357676 278740 357682 278752
rect 357802 278740 357808 278752
rect 357860 278740 357866 278792
rect 386601 278783 386659 278789
rect 386601 278749 386613 278783
rect 386647 278780 386659 278783
rect 386690 278780 386696 278792
rect 386647 278752 386696 278780
rect 386647 278749 386659 278752
rect 386601 278743 386659 278749
rect 386690 278740 386696 278752
rect 386748 278740 386754 278792
rect 397638 278740 397644 278792
rect 397696 278780 397702 278792
rect 397730 278780 397736 278792
rect 397696 278752 397736 278780
rect 397696 278740 397702 278752
rect 397730 278740 397736 278752
rect 397788 278740 397794 278792
rect 408681 278783 408739 278789
rect 408681 278749 408693 278783
rect 408727 278780 408739 278783
rect 408770 278780 408776 278792
rect 408727 278752 408776 278780
rect 408727 278749 408739 278752
rect 408681 278743 408739 278749
rect 408770 278740 408776 278752
rect 408828 278740 408834 278792
rect 451274 278740 451280 278792
rect 451332 278780 451338 278792
rect 451550 278780 451556 278792
rect 451332 278752 451556 278780
rect 451332 278740 451338 278752
rect 451550 278740 451556 278752
rect 451608 278740 451614 278792
rect 270586 278712 270592 278724
rect 270547 278684 270592 278712
rect 270586 278672 270592 278684
rect 270644 278672 270650 278724
rect 397638 278576 397644 278588
rect 397599 278548 397644 278576
rect 397638 278536 397644 278548
rect 397696 278536 397702 278588
rect 254121 277423 254179 277429
rect 254121 277389 254133 277423
rect 254167 277420 254179 277423
rect 254210 277420 254216 277432
rect 254167 277392 254216 277420
rect 254167 277389 254179 277392
rect 254121 277383 254179 277389
rect 254210 277380 254216 277392
rect 254268 277380 254274 277432
rect 259641 277423 259699 277429
rect 259641 277389 259653 277423
rect 259687 277420 259699 277423
rect 259730 277420 259736 277432
rect 259687 277392 259736 277420
rect 259687 277389 259699 277392
rect 259641 277383 259699 277389
rect 259730 277380 259736 277392
rect 259788 277380 259794 277432
rect 356422 277380 356428 277432
rect 356480 277420 356486 277432
rect 356698 277420 356704 277432
rect 356480 277392 356704 277420
rect 356480 277380 356486 277392
rect 356698 277380 356704 277392
rect 356756 277380 356762 277432
rect 545666 274932 545672 274984
rect 545724 274972 545730 274984
rect 550542 274972 550548 274984
rect 545724 274944 550548 274972
rect 545724 274932 545730 274944
rect 550542 274932 550548 274944
rect 550600 274932 550606 274984
rect 369762 274796 369768 274848
rect 369820 274836 369826 274848
rect 370130 274836 370136 274848
rect 369820 274808 370136 274836
rect 369820 274796 369826 274808
rect 370130 274796 370136 274808
rect 370188 274796 370194 274848
rect 295426 273952 295432 273964
rect 295387 273924 295432 273952
rect 295426 273912 295432 273924
rect 295484 273912 295490 273964
rect 451550 273748 451556 273760
rect 451511 273720 451556 273748
rect 451550 273708 451556 273720
rect 451608 273708 451614 273760
rect 232130 273300 232136 273352
rect 232188 273340 232194 273352
rect 232406 273340 232412 273352
rect 232188 273312 232412 273340
rect 232188 273300 232194 273312
rect 232406 273300 232412 273312
rect 232464 273300 232470 273352
rect 330018 273300 330024 273352
rect 330076 273300 330082 273352
rect 356422 273340 356428 273352
rect 356383 273312 356428 273340
rect 356422 273300 356428 273312
rect 356480 273300 356486 273352
rect 357618 273300 357624 273352
rect 357676 273300 357682 273352
rect 367370 273300 367376 273352
rect 367428 273300 367434 273352
rect 408770 273340 408776 273352
rect 408696 273312 408776 273340
rect 236270 273232 236276 273284
rect 236328 273232 236334 273284
rect 236181 273139 236239 273145
rect 236181 273105 236193 273139
rect 236227 273136 236239 273139
rect 236288 273136 236316 273232
rect 330036 273216 330064 273300
rect 357636 273216 357664 273300
rect 367388 273216 367416 273300
rect 386598 273272 386604 273284
rect 386559 273244 386604 273272
rect 386598 273232 386604 273244
rect 386656 273232 386662 273284
rect 408696 273216 408724 273312
rect 408770 273300 408776 273312
rect 408828 273300 408834 273352
rect 244458 273164 244464 273216
rect 244516 273164 244522 273216
rect 272058 273164 272064 273216
rect 272116 273164 272122 273216
rect 283098 273164 283104 273216
rect 283156 273164 283162 273216
rect 294138 273164 294144 273216
rect 294196 273164 294202 273216
rect 330018 273164 330024 273216
rect 330076 273164 330082 273216
rect 334342 273204 334348 273216
rect 334303 273176 334348 273204
rect 334342 273164 334348 273176
rect 334400 273164 334406 273216
rect 357618 273164 357624 273216
rect 357676 273164 357682 273216
rect 367370 273164 367376 273216
rect 367428 273164 367434 273216
rect 376938 273164 376944 273216
rect 376996 273164 377002 273216
rect 400398 273164 400404 273216
rect 400456 273204 400462 273216
rect 400582 273204 400588 273216
rect 400456 273176 400588 273204
rect 400456 273164 400462 273176
rect 400582 273164 400588 273176
rect 400640 273164 400646 273216
rect 408678 273164 408684 273216
rect 408736 273164 408742 273216
rect 236227 273108 236316 273136
rect 236227 273105 236239 273108
rect 236181 273099 236239 273105
rect 244476 273080 244504 273164
rect 272076 273080 272104 273164
rect 283116 273080 283144 273164
rect 294156 273080 294184 273164
rect 376956 273080 376984 273164
rect 244458 273028 244464 273080
rect 244516 273028 244522 273080
rect 249978 273028 249984 273080
rect 250036 273028 250042 273080
rect 272058 273028 272064 273080
rect 272116 273028 272122 273080
rect 283098 273028 283104 273080
rect 283156 273028 283162 273080
rect 294138 273028 294144 273080
rect 294196 273028 294202 273080
rect 376938 273028 376944 273080
rect 376996 273028 377002 273080
rect 249996 272944 250024 273028
rect 249978 272892 249984 272944
rect 250036 272892 250042 272944
rect 321738 272184 321744 272196
rect 321699 272156 321744 272184
rect 321738 272144 321744 272156
rect 321796 272144 321802 272196
rect 327258 272184 327264 272196
rect 327219 272156 327264 272184
rect 327258 272144 327264 272156
rect 327316 272144 327322 272196
rect 232130 271844 232136 271856
rect 232091 271816 232136 271844
rect 232130 271804 232136 271816
rect 232188 271804 232194 271856
rect 241790 270552 241796 270564
rect 241751 270524 241796 270552
rect 241790 270512 241796 270524
rect 241848 270512 241854 270564
rect 288618 270552 288624 270564
rect 288579 270524 288624 270552
rect 288618 270512 288624 270524
rect 288676 270512 288682 270564
rect 305178 270552 305184 270564
rect 305139 270524 305184 270552
rect 305178 270512 305184 270524
rect 305236 270512 305242 270564
rect 309318 270512 309324 270564
rect 309376 270552 309382 270564
rect 309594 270552 309600 270564
rect 309376 270524 309600 270552
rect 309376 270512 309382 270524
rect 309594 270512 309600 270524
rect 309652 270512 309658 270564
rect 310698 270552 310704 270564
rect 310659 270524 310704 270552
rect 310698 270512 310704 270524
rect 310756 270512 310762 270564
rect 346578 270552 346584 270564
rect 346539 270524 346584 270552
rect 346578 270512 346584 270524
rect 346636 270512 346642 270564
rect 381078 270552 381084 270564
rect 381039 270524 381084 270552
rect 381078 270512 381084 270524
rect 381136 270512 381142 270564
rect 382458 270552 382464 270564
rect 382419 270524 382464 270552
rect 382458 270512 382464 270524
rect 382516 270512 382522 270564
rect 416869 270555 416927 270561
rect 416869 270521 416881 270555
rect 416915 270552 416927 270555
rect 416958 270552 416964 270564
rect 416915 270524 416964 270552
rect 416915 270521 416927 270524
rect 416869 270515 416927 270521
rect 416958 270512 416964 270524
rect 417016 270512 417022 270564
rect 433613 270555 433671 270561
rect 433613 270521 433625 270555
rect 433659 270552 433671 270555
rect 433702 270552 433708 270564
rect 433659 270524 433708 270552
rect 433659 270521 433671 270524
rect 433613 270515 433671 270521
rect 433702 270512 433708 270524
rect 433760 270512 433766 270564
rect 466549 270555 466607 270561
rect 466549 270521 466561 270555
rect 466595 270552 466607 270555
rect 466638 270552 466644 270564
rect 466595 270524 466644 270552
rect 466595 270521 466607 270524
rect 466549 270515 466607 270521
rect 466638 270512 466644 270524
rect 466696 270512 466702 270564
rect 472069 270555 472127 270561
rect 472069 270521 472081 270555
rect 472115 270552 472127 270555
rect 472158 270552 472164 270564
rect 472115 270524 472164 270552
rect 472115 270521 472127 270524
rect 472069 270515 472127 270521
rect 472158 270512 472164 270524
rect 472216 270512 472222 270564
rect 243078 270484 243084 270496
rect 243039 270456 243084 270484
rect 243078 270444 243084 270456
rect 243136 270444 243142 270496
rect 252738 270484 252744 270496
rect 252699 270456 252744 270484
rect 252738 270444 252744 270456
rect 252796 270444 252802 270496
rect 267090 270484 267096 270496
rect 267051 270456 267096 270484
rect 267090 270444 267096 270456
rect 267148 270444 267154 270496
rect 356422 270484 356428 270496
rect 356383 270456 356428 270484
rect 356422 270444 356428 270456
rect 356480 270444 356486 270496
rect 400493 270487 400551 270493
rect 400493 270453 400505 270487
rect 400539 270484 400551 270487
rect 400582 270484 400588 270496
rect 400539 270456 400588 270484
rect 400539 270453 400551 270456
rect 400493 270447 400551 270453
rect 400582 270444 400588 270456
rect 400640 270444 400646 270496
rect 309318 270416 309324 270428
rect 309279 270388 309324 270416
rect 309318 270376 309324 270388
rect 309376 270376 309382 270428
rect 381078 270416 381084 270428
rect 381039 270388 381084 270416
rect 381078 270376 381084 270388
rect 381136 270376 381142 270428
rect 386598 269192 386604 269204
rect 386559 269164 386604 269192
rect 386598 269152 386604 269164
rect 386656 269152 386662 269204
rect 287238 269084 287244 269136
rect 287296 269124 287302 269136
rect 287422 269124 287428 269136
rect 287296 269096 287428 269124
rect 287296 269084 287302 269096
rect 287422 269084 287428 269096
rect 287480 269084 287486 269136
rect 393222 269084 393228 269136
rect 393280 269124 393286 269136
rect 393406 269124 393412 269136
rect 393280 269096 393412 269124
rect 393280 269084 393286 269096
rect 393406 269084 393412 269096
rect 393464 269084 393470 269136
rect 397641 269127 397699 269133
rect 397641 269093 397653 269127
rect 397687 269124 397699 269127
rect 397914 269124 397920 269136
rect 397687 269096 397920 269124
rect 397687 269093 397699 269096
rect 397641 269087 397699 269093
rect 397914 269084 397920 269096
rect 397972 269084 397978 269136
rect 480162 269084 480168 269136
rect 480220 269124 480226 269136
rect 480346 269124 480352 269136
rect 480220 269096 480352 269124
rect 480220 269084 480226 269096
rect 480346 269084 480352 269096
rect 480404 269084 480410 269136
rect 281810 269056 281816 269068
rect 281771 269028 281816 269056
rect 281810 269016 281816 269028
rect 281868 269016 281874 269068
rect 292666 269056 292672 269068
rect 292627 269028 292672 269056
rect 292666 269016 292672 269028
rect 292724 269016 292730 269068
rect 375190 269016 375196 269068
rect 375248 269056 375254 269068
rect 375650 269056 375656 269068
rect 375248 269028 375656 269056
rect 375248 269016 375254 269028
rect 375650 269016 375656 269028
rect 375708 269016 375714 269068
rect 347866 267724 347872 267776
rect 347924 267764 347930 267776
rect 348234 267764 348240 267776
rect 347924 267736 348240 267764
rect 347924 267724 347930 267736
rect 348234 267724 348240 267736
rect 348292 267724 348298 267776
rect 386509 264299 386567 264305
rect 386509 264265 386521 264299
rect 386555 264296 386567 264299
rect 386598 264296 386604 264308
rect 386555 264268 386604 264296
rect 386555 264265 386567 264268
rect 386509 264259 386567 264265
rect 386598 264256 386604 264268
rect 386656 264256 386662 264308
rect 392029 264299 392087 264305
rect 392029 264265 392041 264299
rect 392075 264296 392087 264299
rect 392210 264296 392216 264308
rect 392075 264268 392216 264296
rect 392075 264265 392087 264268
rect 392029 264259 392087 264265
rect 392210 264256 392216 264268
rect 392268 264256 392274 264308
rect 236181 263687 236239 263693
rect 236181 263653 236193 263687
rect 236227 263684 236239 263687
rect 236227 263656 236316 263684
rect 236227 263653 236239 263656
rect 236181 263647 236239 263653
rect 233326 263576 233332 263628
rect 233384 263616 233390 263628
rect 233510 263616 233516 263628
rect 233384 263588 233516 263616
rect 233384 263576 233390 263588
rect 233510 263576 233516 263588
rect 233568 263576 233574 263628
rect 235994 263508 236000 263560
rect 236052 263548 236058 263560
rect 236288 263548 236316 263656
rect 356422 263644 356428 263696
rect 356480 263644 356486 263696
rect 324406 263616 324412 263628
rect 324367 263588 324412 263616
rect 324406 263576 324412 263588
rect 324464 263576 324470 263628
rect 334342 263576 334348 263628
rect 334400 263576 334406 263628
rect 342530 263616 342536 263628
rect 342491 263588 342536 263616
rect 342530 263576 342536 263588
rect 342588 263576 342594 263628
rect 353478 263576 353484 263628
rect 353536 263576 353542 263628
rect 236052 263520 236316 263548
rect 236052 263508 236058 263520
rect 331306 263508 331312 263560
rect 331364 263548 331370 263560
rect 331364 263520 331536 263548
rect 331364 263508 331370 263520
rect 331508 263492 331536 263520
rect 295429 263483 295487 263489
rect 295429 263449 295441 263483
rect 295475 263480 295487 263483
rect 295610 263480 295616 263492
rect 295475 263452 295616 263480
rect 295475 263449 295487 263452
rect 295429 263443 295487 263449
rect 295610 263440 295616 263452
rect 295668 263440 295674 263492
rect 331490 263440 331496 263492
rect 331548 263440 331554 263492
rect 334360 263480 334388 263576
rect 334434 263480 334440 263492
rect 334360 263452 334440 263480
rect 334434 263440 334440 263452
rect 334492 263440 334498 263492
rect 353496 263480 353524 263576
rect 356440 263548 356468 263644
rect 408678 263576 408684 263628
rect 408736 263576 408742 263628
rect 422294 263576 422300 263628
rect 422352 263616 422358 263628
rect 422478 263616 422484 263628
rect 422352 263588 422484 263616
rect 422352 263576 422358 263588
rect 422478 263576 422484 263588
rect 422536 263576 422542 263628
rect 427814 263576 427820 263628
rect 427872 263616 427878 263628
rect 427998 263616 428004 263628
rect 427872 263588 428004 263616
rect 427872 263576 427878 263588
rect 427998 263576 428004 263588
rect 428056 263576 428062 263628
rect 356514 263548 356520 263560
rect 356440 263520 356520 263548
rect 356514 263508 356520 263520
rect 356572 263508 356578 263560
rect 353570 263480 353576 263492
rect 353496 263452 353576 263480
rect 353570 263440 353576 263452
rect 353628 263440 353634 263492
rect 408696 263480 408724 263576
rect 408770 263480 408776 263492
rect 408696 263452 408776 263480
rect 408770 263440 408776 263452
rect 408828 263440 408834 263492
rect 451550 263480 451556 263492
rect 451511 263452 451556 263480
rect 451550 263440 451556 263452
rect 451608 263440 451614 263492
rect 232133 262259 232191 262265
rect 232133 262225 232145 262259
rect 232179 262256 232191 262259
rect 232314 262256 232320 262268
rect 232179 262228 232320 262256
rect 232179 262225 232191 262228
rect 232133 262219 232191 262225
rect 232314 262216 232320 262228
rect 232372 262216 232378 262268
rect 243081 260899 243139 260905
rect 243081 260865 243093 260899
rect 243127 260896 243139 260899
rect 243170 260896 243176 260908
rect 243127 260868 243176 260896
rect 243127 260865 243139 260868
rect 243081 260859 243139 260865
rect 243170 260856 243176 260868
rect 243228 260856 243234 260908
rect 252738 260896 252744 260908
rect 252699 260868 252744 260896
rect 252738 260856 252744 260868
rect 252796 260856 252802 260908
rect 267090 260896 267096 260908
rect 267051 260868 267096 260896
rect 267090 260856 267096 260868
rect 267148 260856 267154 260908
rect 270589 260899 270647 260905
rect 270589 260865 270601 260899
rect 270635 260896 270647 260899
rect 270770 260896 270776 260908
rect 270635 260868 270776 260896
rect 270635 260865 270647 260868
rect 270589 260859 270647 260865
rect 270770 260856 270776 260868
rect 270828 260856 270834 260908
rect 309321 260899 309379 260905
rect 309321 260865 309333 260899
rect 309367 260896 309379 260899
rect 309410 260896 309416 260908
rect 309367 260868 309416 260896
rect 309367 260865 309379 260868
rect 309321 260859 309379 260865
rect 309410 260856 309416 260868
rect 309468 260856 309474 260908
rect 324406 260896 324412 260908
rect 324367 260868 324412 260896
rect 324406 260856 324412 260868
rect 324464 260856 324470 260908
rect 342530 260896 342536 260908
rect 342491 260868 342536 260896
rect 342530 260856 342536 260868
rect 342588 260856 342594 260908
rect 359090 260856 359096 260908
rect 359148 260896 359154 260908
rect 359182 260896 359188 260908
rect 359148 260868 359188 260896
rect 359148 260856 359154 260868
rect 359182 260856 359188 260868
rect 359240 260856 359246 260908
rect 381081 260899 381139 260905
rect 381081 260865 381093 260899
rect 381127 260896 381139 260899
rect 381170 260896 381176 260908
rect 381127 260868 381176 260896
rect 381127 260865 381139 260868
rect 381081 260859 381139 260865
rect 381170 260856 381176 260868
rect 381228 260856 381234 260908
rect 397638 260856 397644 260908
rect 397696 260896 397702 260908
rect 397914 260896 397920 260908
rect 397696 260868 397920 260896
rect 397696 260856 397702 260868
rect 397914 260856 397920 260868
rect 397972 260856 397978 260908
rect 400490 260896 400496 260908
rect 400451 260868 400496 260896
rect 400490 260856 400496 260868
rect 400548 260856 400554 260908
rect 241790 260828 241796 260840
rect 241751 260800 241796 260828
rect 241790 260788 241796 260800
rect 241848 260788 241854 260840
rect 265250 260828 265256 260840
rect 265211 260800 265256 260828
rect 265250 260788 265256 260800
rect 265308 260788 265314 260840
rect 272058 260828 272064 260840
rect 272019 260800 272064 260828
rect 272058 260788 272064 260800
rect 272116 260788 272122 260840
rect 277578 260788 277584 260840
rect 277636 260828 277642 260840
rect 277670 260828 277676 260840
rect 277636 260800 277676 260828
rect 277636 260788 277642 260800
rect 277670 260788 277676 260800
rect 277728 260788 277734 260840
rect 288618 260828 288624 260840
rect 288579 260800 288624 260828
rect 288618 260788 288624 260800
rect 288676 260788 288682 260840
rect 294138 260828 294144 260840
rect 294099 260800 294144 260828
rect 294138 260788 294144 260800
rect 294196 260788 294202 260840
rect 295521 260831 295579 260837
rect 295521 260797 295533 260831
rect 295567 260828 295579 260831
rect 295610 260828 295616 260840
rect 295567 260800 295616 260828
rect 295567 260797 295579 260800
rect 295521 260791 295579 260797
rect 295610 260788 295616 260800
rect 295668 260788 295674 260840
rect 305178 260828 305184 260840
rect 305139 260800 305184 260828
rect 305178 260788 305184 260800
rect 305236 260788 305242 260840
rect 310698 260828 310704 260840
rect 310659 260800 310704 260828
rect 310698 260788 310704 260800
rect 310756 260788 310762 260840
rect 318978 260788 318984 260840
rect 319036 260828 319042 260840
rect 319070 260828 319076 260840
rect 319036 260800 319076 260828
rect 319036 260788 319042 260800
rect 319070 260788 319076 260800
rect 319128 260788 319134 260840
rect 321738 260828 321744 260840
rect 321699 260800 321744 260828
rect 321738 260788 321744 260800
rect 321796 260788 321802 260840
rect 327258 260828 327264 260840
rect 327219 260800 327264 260828
rect 327258 260788 327264 260800
rect 327316 260788 327322 260840
rect 331122 260788 331128 260840
rect 331180 260828 331186 260840
rect 331490 260828 331496 260840
rect 331180 260800 331496 260828
rect 331180 260788 331186 260800
rect 331490 260788 331496 260800
rect 331548 260788 331554 260840
rect 334345 260831 334403 260837
rect 334345 260797 334357 260831
rect 334391 260828 334403 260831
rect 334434 260828 334440 260840
rect 334391 260800 334440 260828
rect 334391 260797 334403 260800
rect 334345 260791 334403 260797
rect 334434 260788 334440 260800
rect 334492 260788 334498 260840
rect 346578 260828 346584 260840
rect 346539 260800 346584 260828
rect 346578 260788 346584 260800
rect 346636 260788 346642 260840
rect 382458 260828 382464 260840
rect 382419 260800 382464 260828
rect 382458 260788 382464 260800
rect 382516 260788 382522 260840
rect 416866 260828 416872 260840
rect 416827 260800 416872 260828
rect 416866 260788 416872 260800
rect 416924 260788 416930 260840
rect 433610 260828 433616 260840
rect 433571 260800 433616 260828
rect 433610 260788 433616 260800
rect 433668 260788 433674 260840
rect 466546 260828 466552 260840
rect 466507 260800 466552 260828
rect 466546 260788 466552 260800
rect 466604 260788 466610 260840
rect 472066 260828 472072 260840
rect 472027 260800 472072 260828
rect 472066 260788 472072 260800
rect 472124 260788 472130 260840
rect 292669 260763 292727 260769
rect 292669 260729 292681 260763
rect 292715 260760 292727 260763
rect 292758 260760 292764 260772
rect 292715 260732 292764 260760
rect 292715 260729 292727 260732
rect 292669 260723 292727 260729
rect 292758 260720 292764 260732
rect 292816 260720 292822 260772
rect 309321 260763 309379 260769
rect 309321 260729 309333 260763
rect 309367 260760 309379 260763
rect 309410 260760 309416 260772
rect 309367 260732 309416 260760
rect 309367 260729 309379 260732
rect 309321 260723 309379 260729
rect 309410 260720 309416 260732
rect 309468 260720 309474 260772
rect 342441 260763 342499 260769
rect 342441 260729 342453 260763
rect 342487 260760 342499 260763
rect 342530 260760 342536 260772
rect 342487 260732 342536 260760
rect 342487 260729 342499 260732
rect 342441 260723 342499 260729
rect 342530 260720 342536 260732
rect 342588 260720 342594 260772
rect 281813 259471 281871 259477
rect 281813 259437 281825 259471
rect 281859 259468 281871 259471
rect 281994 259468 282000 259480
rect 281859 259440 282000 259468
rect 281859 259437 281871 259440
rect 281813 259431 281871 259437
rect 281994 259428 282000 259440
rect 282052 259428 282058 259480
rect 351822 259428 351828 259480
rect 351880 259468 351886 259480
rect 352006 259468 352012 259480
rect 351880 259440 352012 259468
rect 351880 259428 351886 259440
rect 352006 259428 352012 259440
rect 352064 259428 352070 259480
rect 386506 259468 386512 259480
rect 386467 259440 386512 259468
rect 386506 259428 386512 259440
rect 386564 259428 386570 259480
rect 392026 259468 392032 259480
rect 391987 259440 392032 259468
rect 392026 259428 392032 259440
rect 392084 259428 392090 259480
rect 393222 259428 393228 259480
rect 393280 259468 393286 259480
rect 393406 259468 393412 259480
rect 393280 259440 393412 259468
rect 393280 259428 393286 259440
rect 393406 259428 393412 259440
rect 393464 259428 393470 259480
rect 451550 259400 451556 259412
rect 451511 259372 451556 259400
rect 451550 259360 451556 259372
rect 451608 259360 451614 259412
rect 356422 258000 356428 258052
rect 356480 258040 356486 258052
rect 356606 258040 356612 258052
rect 356480 258012 356612 258040
rect 356480 258000 356486 258012
rect 356606 258000 356612 258012
rect 356664 258000 356670 258052
rect 408770 258000 408776 258052
rect 408828 258040 408834 258052
rect 408954 258040 408960 258052
rect 408828 258012 408960 258040
rect 408828 258000 408834 258012
rect 408954 258000 408960 258012
rect 409012 258000 409018 258052
rect 254121 254031 254179 254037
rect 254121 253997 254133 254031
rect 254167 254028 254179 254031
rect 254210 254028 254216 254040
rect 254167 254000 254216 254028
rect 254167 253997 254179 254000
rect 254121 253991 254179 253997
rect 254210 253988 254216 254000
rect 254268 253988 254274 254040
rect 259641 254031 259699 254037
rect 259641 253997 259653 254031
rect 259687 254028 259699 254031
rect 259730 254028 259736 254040
rect 259687 254000 259736 254028
rect 259687 253997 259699 254000
rect 259641 253991 259699 253997
rect 259730 253988 259736 254000
rect 259788 253988 259794 254040
rect 261018 253988 261024 254040
rect 261076 253988 261082 254040
rect 330018 253988 330024 254040
rect 330076 253988 330082 254040
rect 370041 254031 370099 254037
rect 370041 253997 370053 254031
rect 370087 254028 370099 254031
rect 370130 254028 370136 254040
rect 370087 254000 370136 254028
rect 370087 253997 370099 254000
rect 370041 253991 370099 253997
rect 370130 253988 370136 254000
rect 370188 253988 370194 254040
rect 375561 254031 375619 254037
rect 375561 253997 375573 254031
rect 375607 254028 375619 254031
rect 375650 254028 375656 254040
rect 375607 254000 375656 254028
rect 375607 253997 375619 254000
rect 375561 253991 375619 253997
rect 375650 253988 375656 254000
rect 375708 253988 375714 254040
rect 232130 253920 232136 253972
rect 232188 253960 232194 253972
rect 232314 253960 232320 253972
rect 232188 253932 232320 253960
rect 232188 253920 232194 253932
rect 232314 253920 232320 253932
rect 232372 253920 232378 253972
rect 261036 253904 261064 253988
rect 330036 253904 330064 253988
rect 397549 253963 397607 253969
rect 397549 253929 397561 253963
rect 397595 253960 397607 253963
rect 397730 253960 397736 253972
rect 397595 253932 397736 253960
rect 397595 253929 397607 253932
rect 397549 253923 397607 253929
rect 397730 253920 397736 253932
rect 397788 253920 397794 253972
rect 236270 253892 236276 253904
rect 236231 253864 236276 253892
rect 236270 253852 236276 253864
rect 236328 253852 236334 253904
rect 244458 253852 244464 253904
rect 244516 253852 244522 253904
rect 261018 253852 261024 253904
rect 261076 253852 261082 253904
rect 283098 253852 283104 253904
rect 283156 253852 283162 253904
rect 330018 253852 330024 253904
rect 330076 253852 330082 253904
rect 376938 253852 376944 253904
rect 376996 253852 377002 253904
rect 387978 253852 387984 253904
rect 388036 253852 388042 253904
rect 400398 253852 400404 253904
rect 400456 253892 400462 253904
rect 400582 253892 400588 253904
rect 400456 253864 400588 253892
rect 400456 253852 400462 253864
rect 400582 253852 400588 253864
rect 400640 253852 400646 253904
rect 244476 253768 244504 253852
rect 283116 253768 283144 253852
rect 376956 253768 376984 253852
rect 387996 253768 388024 253852
rect 244458 253716 244464 253768
rect 244516 253716 244522 253768
rect 249978 253716 249984 253768
rect 250036 253716 250042 253768
rect 267090 253716 267096 253768
rect 267148 253716 267154 253768
rect 283098 253716 283104 253768
rect 283156 253716 283162 253768
rect 376938 253716 376944 253768
rect 376996 253716 377002 253768
rect 387978 253716 387984 253768
rect 388036 253716 388042 253768
rect 249996 253632 250024 253716
rect 267108 253688 267136 253716
rect 267182 253688 267188 253700
rect 267108 253660 267188 253688
rect 267182 253648 267188 253660
rect 267240 253648 267246 253700
rect 249978 253580 249984 253632
rect 250036 253580 250042 253632
rect 334342 251308 334348 251320
rect 334303 251280 334348 251308
rect 334342 251268 334348 251280
rect 334400 251268 334406 251320
rect 381262 251308 381268 251320
rect 381096 251280 381268 251308
rect 381096 251252 381124 251280
rect 381262 251268 381268 251280
rect 381320 251268 381326 251320
rect 393222 251308 393228 251320
rect 393148 251280 393228 251308
rect 241790 251240 241796 251252
rect 241751 251212 241796 251240
rect 241790 251200 241796 251212
rect 241848 251200 241854 251252
rect 265250 251240 265256 251252
rect 265211 251212 265256 251240
rect 265250 251200 265256 251212
rect 265308 251200 265314 251252
rect 270678 251200 270684 251252
rect 270736 251240 270742 251252
rect 270954 251240 270960 251252
rect 270736 251212 270960 251240
rect 270736 251200 270742 251212
rect 270954 251200 270960 251212
rect 271012 251200 271018 251252
rect 272058 251240 272064 251252
rect 272019 251212 272064 251240
rect 272058 251200 272064 251212
rect 272116 251200 272122 251252
rect 288618 251240 288624 251252
rect 288579 251212 288624 251240
rect 288618 251200 288624 251212
rect 288676 251200 288682 251252
rect 294138 251240 294144 251252
rect 294099 251212 294144 251240
rect 294138 251200 294144 251212
rect 294196 251200 294202 251252
rect 295518 251240 295524 251252
rect 295479 251212 295524 251240
rect 295518 251200 295524 251212
rect 295576 251200 295582 251252
rect 305178 251240 305184 251252
rect 305139 251212 305184 251240
rect 305178 251200 305184 251212
rect 305236 251200 305242 251252
rect 309318 251240 309324 251252
rect 309279 251212 309324 251240
rect 309318 251200 309324 251212
rect 309376 251200 309382 251252
rect 310698 251240 310704 251252
rect 310659 251212 310704 251240
rect 310698 251200 310704 251212
rect 310756 251200 310762 251252
rect 321738 251240 321744 251252
rect 321699 251212 321744 251240
rect 321738 251200 321744 251212
rect 321796 251200 321802 251252
rect 327258 251240 327264 251252
rect 327219 251212 327264 251240
rect 327258 251200 327264 251212
rect 327316 251200 327322 251252
rect 342438 251240 342444 251252
rect 342399 251212 342444 251240
rect 342438 251200 342444 251212
rect 342496 251200 342502 251252
rect 346578 251240 346584 251252
rect 346539 251212 346584 251240
rect 346578 251200 346584 251212
rect 346636 251200 346642 251252
rect 352006 251200 352012 251252
rect 352064 251240 352070 251252
rect 352098 251240 352104 251252
rect 352064 251212 352104 251240
rect 352064 251200 352070 251212
rect 352098 251200 352104 251212
rect 352156 251200 352162 251252
rect 381078 251200 381084 251252
rect 381136 251200 381142 251252
rect 382458 251240 382464 251252
rect 382419 251212 382464 251240
rect 382458 251200 382464 251212
rect 382516 251200 382522 251252
rect 292758 251172 292764 251184
rect 292719 251144 292764 251172
rect 292758 251132 292764 251144
rect 292816 251132 292822 251184
rect 298278 251132 298284 251184
rect 298336 251172 298342 251184
rect 298554 251172 298560 251184
rect 298336 251144 298560 251172
rect 298336 251132 298342 251144
rect 298554 251132 298560 251144
rect 298612 251132 298618 251184
rect 334342 251172 334348 251184
rect 334303 251144 334348 251172
rect 334342 251132 334348 251144
rect 334400 251132 334406 251184
rect 353570 251172 353576 251184
rect 353531 251144 353576 251172
rect 353570 251132 353576 251144
rect 353628 251132 353634 251184
rect 386506 251132 386512 251184
rect 386564 251172 386570 251184
rect 386874 251172 386880 251184
rect 386564 251144 386880 251172
rect 386564 251132 386570 251144
rect 386874 251132 386880 251144
rect 386932 251132 386938 251184
rect 393148 251116 393176 251280
rect 393222 251268 393228 251280
rect 393280 251268 393286 251320
rect 416869 251243 416927 251249
rect 416869 251209 416881 251243
rect 416915 251240 416927 251243
rect 416958 251240 416964 251252
rect 416915 251212 416964 251240
rect 416915 251209 416927 251212
rect 416869 251203 416927 251209
rect 416958 251200 416964 251212
rect 417016 251200 417022 251252
rect 433613 251243 433671 251249
rect 433613 251209 433625 251243
rect 433659 251240 433671 251243
rect 433702 251240 433708 251252
rect 433659 251212 433708 251240
rect 433659 251209 433671 251212
rect 433613 251203 433671 251209
rect 433702 251200 433708 251212
rect 433760 251200 433766 251252
rect 466549 251243 466607 251249
rect 466549 251209 466561 251243
rect 466595 251240 466607 251243
rect 466638 251240 466644 251252
rect 466595 251212 466644 251240
rect 466595 251209 466607 251212
rect 466549 251203 466607 251209
rect 466638 251200 466644 251212
rect 466696 251200 466702 251252
rect 472069 251243 472127 251249
rect 472069 251209 472081 251243
rect 472115 251240 472127 251243
rect 472158 251240 472164 251252
rect 472115 251212 472164 251240
rect 472115 251209 472127 251212
rect 472069 251203 472127 251209
rect 472158 251200 472164 251212
rect 472216 251200 472222 251252
rect 400493 251175 400551 251181
rect 400493 251141 400505 251175
rect 400539 251172 400551 251175
rect 400582 251172 400588 251184
rect 400539 251144 400588 251172
rect 400539 251141 400551 251144
rect 400493 251135 400551 251141
rect 400582 251132 400588 251144
rect 400640 251132 400646 251184
rect 407666 251132 407672 251184
rect 407724 251172 407730 251184
rect 407758 251172 407764 251184
rect 407724 251144 407764 251172
rect 407724 251132 407730 251144
rect 407758 251132 407764 251144
rect 407816 251132 407822 251184
rect 393130 251064 393136 251116
rect 393188 251064 393194 251116
rect 348050 250084 348056 250096
rect 348011 250056 348056 250084
rect 348050 250044 348056 250056
rect 348108 250044 348114 250096
rect 359090 249948 359096 249960
rect 359016 249920 359096 249948
rect 359016 249892 359044 249920
rect 359090 249908 359096 249920
rect 359148 249908 359154 249960
rect 287146 249840 287152 249892
rect 287204 249880 287210 249892
rect 287330 249880 287336 249892
rect 287204 249852 287336 249880
rect 287204 249840 287210 249852
rect 287330 249840 287336 249852
rect 287388 249840 287394 249892
rect 358998 249840 359004 249892
rect 359056 249840 359062 249892
rect 364518 249840 364524 249892
rect 364576 249880 364582 249892
rect 364610 249880 364616 249892
rect 364576 249852 364616 249880
rect 364576 249840 364582 249852
rect 364610 249840 364616 249852
rect 364668 249840 364674 249892
rect 397546 249812 397552 249824
rect 397507 249784 397552 249812
rect 397546 249772 397552 249784
rect 397604 249772 397610 249824
rect 480162 249772 480168 249824
rect 480220 249812 480226 249824
rect 480346 249812 480352 249824
rect 480220 249784 480352 249812
rect 480220 249772 480226 249784
rect 480346 249772 480352 249784
rect 480404 249772 480410 249824
rect 254118 248520 254124 248532
rect 254079 248492 254124 248520
rect 254118 248480 254124 248492
rect 254176 248480 254182 248532
rect 259638 248520 259644 248532
rect 259599 248492 259644 248520
rect 259638 248480 259644 248492
rect 259696 248480 259702 248532
rect 370038 248520 370044 248532
rect 369999 248492 370044 248520
rect 370038 248480 370044 248492
rect 370096 248480 370102 248532
rect 375558 248520 375564 248532
rect 375519 248492 375564 248520
rect 375558 248480 375564 248492
rect 375616 248480 375622 248532
rect 254118 248384 254124 248396
rect 254079 248356 254124 248384
rect 254118 248344 254124 248356
rect 254176 248344 254182 248396
rect 259362 248344 259368 248396
rect 259420 248384 259426 248396
rect 259638 248384 259644 248396
rect 259420 248356 259644 248384
rect 259420 248344 259426 248356
rect 259638 248344 259644 248356
rect 259696 248344 259702 248396
rect 281994 248344 282000 248396
rect 282052 248384 282058 248396
rect 282178 248384 282184 248396
rect 282052 248356 282184 248384
rect 282052 248344 282058 248356
rect 282178 248344 282184 248356
rect 282236 248344 282242 248396
rect 356330 248344 356336 248396
rect 356388 248384 356394 248396
rect 356422 248384 356428 248396
rect 356388 248356 356428 248384
rect 356388 248344 356394 248356
rect 356422 248344 356428 248356
rect 356480 248344 356486 248396
rect 370038 248344 370044 248396
rect 370096 248384 370102 248396
rect 370314 248384 370320 248396
rect 370096 248356 370320 248384
rect 370096 248344 370102 248356
rect 370314 248344 370320 248356
rect 370372 248344 370378 248396
rect 375558 248384 375564 248396
rect 375519 248356 375564 248384
rect 375558 248344 375564 248356
rect 375616 248344 375622 248396
rect 397546 244984 397552 244996
rect 397507 244956 397552 244984
rect 397546 244944 397552 244956
rect 397604 244944 397610 244996
rect 236273 244375 236331 244381
rect 236273 244341 236285 244375
rect 236319 244341 236331 244375
rect 236273 244335 236331 244341
rect 233326 244264 233332 244316
rect 233384 244304 233390 244316
rect 233510 244304 233516 244316
rect 233384 244276 233516 244304
rect 233384 244264 233390 244276
rect 233510 244264 233516 244276
rect 233568 244264 233574 244316
rect 231946 244196 231952 244248
rect 232004 244236 232010 244248
rect 232130 244236 232136 244248
rect 232004 244208 232136 244236
rect 232004 244196 232010 244208
rect 232130 244196 232136 244208
rect 232188 244196 232194 244248
rect 236288 244245 236316 244335
rect 265158 244332 265164 244384
rect 265216 244332 265222 244384
rect 243078 244264 243084 244316
rect 243136 244264 243142 244316
rect 236273 244239 236331 244245
rect 236273 244205 236285 244239
rect 236319 244205 236331 244239
rect 236273 244199 236331 244205
rect 243096 244168 243124 244264
rect 254118 244236 254124 244248
rect 254079 244208 254124 244236
rect 254118 244196 254124 244208
rect 254176 244196 254182 244248
rect 265176 244180 265204 244332
rect 270678 244264 270684 244316
rect 270736 244264 270742 244316
rect 324406 244304 324412 244316
rect 324367 244276 324412 244304
rect 324406 244264 324412 244276
rect 324464 244264 324470 244316
rect 364518 244264 364524 244316
rect 364576 244264 364582 244316
rect 381078 244264 381084 244316
rect 381136 244264 381142 244316
rect 422294 244264 422300 244316
rect 422352 244304 422358 244316
rect 422478 244304 422484 244316
rect 422352 244276 422484 244304
rect 422352 244264 422358 244276
rect 422478 244264 422484 244276
rect 422536 244264 422542 244316
rect 427814 244264 427820 244316
rect 427872 244304 427878 244316
rect 427998 244304 428004 244316
rect 427872 244276 428004 244304
rect 427872 244264 427878 244276
rect 427998 244264 428004 244276
rect 428056 244264 428062 244316
rect 243170 244168 243176 244180
rect 243096 244140 243176 244168
rect 243170 244128 243176 244140
rect 243228 244128 243234 244180
rect 265158 244128 265164 244180
rect 265216 244128 265222 244180
rect 270696 244168 270724 244264
rect 270770 244168 270776 244180
rect 270696 244140 270776 244168
rect 270770 244128 270776 244140
rect 270828 244128 270834 244180
rect 334342 244168 334348 244180
rect 334303 244140 334348 244168
rect 334342 244128 334348 244140
rect 334400 244128 334406 244180
rect 364536 244168 364564 244264
rect 364610 244168 364616 244180
rect 364536 244140 364616 244168
rect 364610 244128 364616 244140
rect 364668 244128 364674 244180
rect 381096 244168 381124 244264
rect 381170 244168 381176 244180
rect 381096 244140 381176 244168
rect 381170 244128 381176 244140
rect 381228 244128 381234 244180
rect 451550 244168 451556 244180
rect 451511 244140 451556 244168
rect 451550 244128 451556 244140
rect 451608 244128 451614 244180
rect 375558 242808 375564 242820
rect 375519 242780 375564 242808
rect 375558 242768 375564 242780
rect 375616 242768 375622 242820
rect 324406 241584 324412 241596
rect 324367 241556 324412 241584
rect 324406 241544 324412 241556
rect 324464 241544 324470 241596
rect 266814 241476 266820 241528
rect 266872 241516 266878 241528
rect 266906 241516 266912 241528
rect 266872 241488 266912 241516
rect 266872 241476 266878 241488
rect 266906 241476 266912 241488
rect 266964 241476 266970 241528
rect 295702 241476 295708 241528
rect 295760 241516 295766 241528
rect 295794 241516 295800 241528
rect 295760 241488 295800 241516
rect 295760 241476 295766 241488
rect 295794 241476 295800 241488
rect 295852 241476 295858 241528
rect 309502 241476 309508 241528
rect 309560 241516 309566 241528
rect 309594 241516 309600 241528
rect 309560 241488 309600 241516
rect 309560 241476 309566 241488
rect 309594 241476 309600 241488
rect 309652 241476 309658 241528
rect 331122 241476 331128 241528
rect 331180 241516 331186 241528
rect 331490 241516 331496 241528
rect 331180 241488 331496 241516
rect 331180 241476 331186 241488
rect 331490 241476 331496 241488
rect 331548 241476 331554 241528
rect 348050 241516 348056 241528
rect 348011 241488 348056 241516
rect 348050 241476 348056 241488
rect 348108 241476 348114 241528
rect 353570 241516 353576 241528
rect 353531 241488 353576 241516
rect 353570 241476 353576 241488
rect 353628 241476 353634 241528
rect 392026 241476 392032 241528
rect 392084 241516 392090 241528
rect 392118 241516 392124 241528
rect 392084 241488 392124 241516
rect 392084 241476 392090 241488
rect 392118 241476 392124 241488
rect 392176 241476 392182 241528
rect 400490 241516 400496 241528
rect 400451 241488 400496 241516
rect 400490 241476 400496 241488
rect 400548 241476 400554 241528
rect 324406 241408 324412 241460
rect 324464 241448 324470 241460
rect 324498 241448 324504 241460
rect 324464 241420 324504 241448
rect 324464 241408 324470 241420
rect 324498 241408 324504 241420
rect 324556 241408 324562 241460
rect 466546 241408 466552 241460
rect 466604 241448 466610 241460
rect 466638 241448 466644 241460
rect 466604 241420 466644 241448
rect 466604 241408 466610 241420
rect 466638 241408 466644 241420
rect 466696 241408 466702 241460
rect 287238 240116 287244 240168
rect 287296 240156 287302 240168
rect 287422 240156 287428 240168
rect 287296 240128 287428 240156
rect 287296 240116 287302 240128
rect 287422 240116 287428 240128
rect 287480 240116 287486 240168
rect 292758 240156 292764 240168
rect 292719 240128 292764 240156
rect 292758 240116 292764 240128
rect 292816 240116 292822 240168
rect 359090 240116 359096 240168
rect 359148 240156 359154 240168
rect 359274 240156 359280 240168
rect 359148 240128 359280 240156
rect 359148 240116 359154 240128
rect 359274 240116 359280 240128
rect 359332 240116 359338 240168
rect 392946 240116 392952 240168
rect 393004 240156 393010 240168
rect 393222 240156 393228 240168
rect 393004 240128 393228 240156
rect 393004 240116 393010 240128
rect 393222 240116 393228 240128
rect 393280 240116 393286 240168
rect 397549 240159 397607 240165
rect 397549 240125 397561 240159
rect 397595 240156 397607 240159
rect 397638 240156 397644 240168
rect 397595 240128 397644 240156
rect 397595 240125 397607 240128
rect 397549 240119 397607 240125
rect 397638 240116 397644 240128
rect 397696 240116 397702 240168
rect 407482 240116 407488 240168
rect 407540 240156 407546 240168
rect 407758 240156 407764 240168
rect 407540 240128 407764 240156
rect 407540 240116 407546 240128
rect 407758 240116 407764 240128
rect 407816 240116 407822 240168
rect 292758 240020 292764 240032
rect 292719 239992 292764 240020
rect 292758 239980 292764 239992
rect 292816 239980 292822 240032
rect 356514 238620 356520 238672
rect 356572 238660 356578 238672
rect 356606 238660 356612 238672
rect 356572 238632 356612 238660
rect 356572 238620 356578 238632
rect 356606 238620 356612 238632
rect 356664 238620 356670 238672
rect 2774 237124 2780 237176
rect 2832 237164 2838 237176
rect 4890 237164 4896 237176
rect 2832 237136 4896 237164
rect 2832 237124 2838 237136
rect 4890 237124 4896 237136
rect 4948 237124 4954 237176
rect 281902 234716 281908 234728
rect 281828 234688 281908 234716
rect 236270 234648 236276 234660
rect 236231 234620 236276 234648
rect 236270 234608 236276 234620
rect 236328 234608 236334 234660
rect 255590 234648 255596 234660
rect 255516 234620 255596 234648
rect 255516 234592 255544 234620
rect 255590 234608 255596 234620
rect 255648 234608 255654 234660
rect 261110 234648 261116 234660
rect 261036 234620 261116 234648
rect 261036 234592 261064 234620
rect 261110 234608 261116 234620
rect 261168 234608 261174 234660
rect 281828 234592 281856 234688
rect 281902 234676 281908 234688
rect 281960 234676 281966 234728
rect 397638 234676 397644 234728
rect 397696 234676 397702 234728
rect 451550 234716 451556 234728
rect 451476 234688 451556 234716
rect 321830 234648 321836 234660
rect 321756 234620 321836 234648
rect 321756 234592 321784 234620
rect 321830 234608 321836 234620
rect 321888 234608 321894 234660
rect 330110 234648 330116 234660
rect 330036 234620 330116 234648
rect 330036 234592 330064 234620
rect 330110 234608 330116 234620
rect 330168 234608 330174 234660
rect 357710 234648 357716 234660
rect 357636 234620 357716 234648
rect 357636 234592 357664 234620
rect 357710 234608 357716 234620
rect 357768 234608 357774 234660
rect 367462 234648 367468 234660
rect 367388 234620 367468 234648
rect 367388 234592 367416 234620
rect 367462 234608 367468 234620
rect 367520 234608 367526 234660
rect 381170 234648 381176 234660
rect 381096 234620 381176 234648
rect 381096 234592 381124 234620
rect 381170 234608 381176 234620
rect 381228 234608 381234 234660
rect 397656 234592 397684 234676
rect 451476 234592 451504 234688
rect 451550 234676 451556 234688
rect 451608 234676 451614 234728
rect 255498 234540 255504 234592
rect 255556 234540 255562 234592
rect 261018 234540 261024 234592
rect 261076 234540 261082 234592
rect 281810 234540 281816 234592
rect 281868 234540 281874 234592
rect 309318 234540 309324 234592
rect 309376 234580 309382 234592
rect 309594 234580 309600 234592
rect 309376 234552 309600 234580
rect 309376 234540 309382 234552
rect 309594 234540 309600 234552
rect 309652 234540 309658 234592
rect 321738 234540 321744 234592
rect 321796 234540 321802 234592
rect 330018 234540 330024 234592
rect 330076 234540 330082 234592
rect 357618 234540 357624 234592
rect 357676 234540 357682 234592
rect 367370 234540 367376 234592
rect 367428 234540 367434 234592
rect 376938 234540 376944 234592
rect 376996 234540 377002 234592
rect 381078 234540 381084 234592
rect 381136 234540 381142 234592
rect 387978 234540 387984 234592
rect 388036 234540 388042 234592
rect 397638 234540 397644 234592
rect 397696 234540 397702 234592
rect 400398 234540 400404 234592
rect 400456 234580 400462 234592
rect 400582 234580 400588 234592
rect 400456 234552 400588 234580
rect 400456 234540 400462 234552
rect 400582 234540 400588 234552
rect 400640 234540 400646 234592
rect 451458 234540 451464 234592
rect 451516 234540 451522 234592
rect 351822 234472 351828 234524
rect 351880 234512 351886 234524
rect 352098 234512 352104 234524
rect 351880 234484 352104 234512
rect 351880 234472 351886 234484
rect 352098 234472 352104 234484
rect 352156 234472 352162 234524
rect 376956 234456 376984 234540
rect 387996 234456 388024 234540
rect 376938 234404 376944 234456
rect 376996 234404 377002 234456
rect 387978 234404 387984 234456
rect 388036 234404 388042 234456
rect 359090 233860 359096 233912
rect 359148 233900 359154 233912
rect 359274 233900 359280 233912
rect 359148 233872 359280 233900
rect 359148 233860 359154 233872
rect 359274 233860 359280 233872
rect 359332 233860 359338 233912
rect 369762 233860 369768 233912
rect 369820 233900 369826 233912
rect 370314 233900 370320 233912
rect 369820 233872 370320 233900
rect 369820 233860 369826 233872
rect 370314 233860 370320 233872
rect 370372 233860 370378 233912
rect 265158 231956 265164 232008
rect 265216 231996 265222 232008
rect 265216 231968 265296 231996
rect 265216 231956 265222 231968
rect 265268 231872 265296 231968
rect 334342 231956 334348 232008
rect 334400 231996 334406 232008
rect 334400 231968 334480 231996
rect 334400 231956 334406 231968
rect 334452 231872 334480 231968
rect 265250 231820 265256 231872
rect 265308 231820 265314 231872
rect 271874 231820 271880 231872
rect 271932 231860 271938 231872
rect 272058 231860 272064 231872
rect 271932 231832 272064 231860
rect 271932 231820 271938 231832
rect 272058 231820 272064 231832
rect 272116 231820 272122 231872
rect 277578 231820 277584 231872
rect 277636 231860 277642 231872
rect 277670 231860 277676 231872
rect 277636 231832 277676 231860
rect 277636 231820 277642 231832
rect 277670 231820 277676 231832
rect 277728 231820 277734 231872
rect 293954 231820 293960 231872
rect 294012 231860 294018 231872
rect 294138 231860 294144 231872
rect 294012 231832 294144 231860
rect 294012 231820 294018 231832
rect 294138 231820 294144 231832
rect 294196 231820 294202 231872
rect 295518 231820 295524 231872
rect 295576 231860 295582 231872
rect 295794 231860 295800 231872
rect 295576 231832 295800 231860
rect 295576 231820 295582 231832
rect 295794 231820 295800 231832
rect 295852 231820 295858 231872
rect 298278 231820 298284 231872
rect 298336 231860 298342 231872
rect 298554 231860 298560 231872
rect 298336 231832 298560 231860
rect 298336 231820 298342 231832
rect 298554 231820 298560 231832
rect 298612 231820 298618 231872
rect 305178 231820 305184 231872
rect 305236 231860 305242 231872
rect 305362 231860 305368 231872
rect 305236 231832 305368 231860
rect 305236 231820 305242 231832
rect 305362 231820 305368 231832
rect 305420 231820 305426 231872
rect 310698 231820 310704 231872
rect 310756 231860 310762 231872
rect 310882 231860 310888 231872
rect 310756 231832 310888 231860
rect 310756 231820 310762 231832
rect 310882 231820 310888 231832
rect 310940 231820 310946 231872
rect 318978 231820 318984 231872
rect 319036 231860 319042 231872
rect 319070 231860 319076 231872
rect 319036 231832 319076 231860
rect 319036 231820 319042 231832
rect 319070 231820 319076 231832
rect 319128 231820 319134 231872
rect 331309 231863 331367 231869
rect 331309 231829 331321 231863
rect 331355 231860 331367 231863
rect 331490 231860 331496 231872
rect 331355 231832 331496 231860
rect 331355 231829 331367 231832
rect 331309 231823 331367 231829
rect 331490 231820 331496 231832
rect 331548 231820 331554 231872
rect 334434 231820 334440 231872
rect 334492 231820 334498 231872
rect 346578 231820 346584 231872
rect 346636 231860 346642 231872
rect 346762 231860 346768 231872
rect 346636 231832 346768 231860
rect 346636 231820 346642 231832
rect 346762 231820 346768 231832
rect 346820 231820 346826 231872
rect 364610 231820 364616 231872
rect 364668 231820 364674 231872
rect 382274 231820 382280 231872
rect 382332 231860 382338 231872
rect 382458 231860 382464 231872
rect 382332 231832 382464 231860
rect 382332 231820 382338 231832
rect 382458 231820 382464 231832
rect 382516 231820 382522 231872
rect 386598 231820 386604 231872
rect 386656 231860 386662 231872
rect 386874 231860 386880 231872
rect 386656 231832 386880 231860
rect 386656 231820 386662 231832
rect 386874 231820 386880 231832
rect 386932 231820 386938 231872
rect 416958 231820 416964 231872
rect 417016 231860 417022 231872
rect 417142 231860 417148 231872
rect 417016 231832 417148 231860
rect 417016 231820 417022 231832
rect 417142 231820 417148 231832
rect 417200 231820 417206 231872
rect 433426 231820 433432 231872
rect 433484 231860 433490 231872
rect 433702 231860 433708 231872
rect 433484 231832 433708 231860
rect 433484 231820 433490 231832
rect 433702 231820 433708 231832
rect 433760 231820 433766 231872
rect 472158 231820 472164 231872
rect 472216 231860 472222 231872
rect 472342 231860 472348 231872
rect 472216 231832 472348 231860
rect 472216 231820 472222 231832
rect 472342 231820 472348 231832
rect 472400 231820 472406 231872
rect 259638 231792 259644 231804
rect 259599 231764 259644 231792
rect 259638 231752 259644 231764
rect 259696 231752 259702 231804
rect 309318 231792 309324 231804
rect 309279 231764 309324 231792
rect 309318 231752 309324 231764
rect 309376 231752 309382 231804
rect 364518 231752 364524 231804
rect 364576 231792 364582 231804
rect 364628 231792 364656 231820
rect 364576 231764 364656 231792
rect 364576 231752 364582 231764
rect 347958 230528 347964 230580
rect 348016 230568 348022 230580
rect 348050 230568 348056 230580
rect 348016 230540 348056 230568
rect 348016 230528 348022 230540
rect 348050 230528 348056 230540
rect 348108 230528 348114 230580
rect 353478 230528 353484 230580
rect 353536 230568 353542 230580
rect 353570 230568 353576 230580
rect 353536 230540 353576 230568
rect 353536 230528 353542 230540
rect 353570 230528 353576 230540
rect 353628 230528 353634 230580
rect 242710 230460 242716 230512
rect 242768 230500 242774 230512
rect 242802 230500 242808 230512
rect 242768 230472 242808 230500
rect 242768 230460 242774 230472
rect 242802 230460 242808 230472
rect 242860 230460 242866 230512
rect 270586 230460 270592 230512
rect 270644 230500 270650 230512
rect 270678 230500 270684 230512
rect 270644 230472 270684 230500
rect 270644 230460 270650 230472
rect 270678 230460 270684 230472
rect 270736 230460 270742 230512
rect 292758 230500 292764 230512
rect 292719 230472 292764 230500
rect 292758 230460 292764 230472
rect 292816 230460 292822 230512
rect 480162 230460 480168 230512
rect 480220 230500 480226 230512
rect 480346 230500 480352 230512
rect 480220 230472 480352 230500
rect 480220 230460 480226 230472
rect 480346 230460 480352 230472
rect 480404 230460 480410 230512
rect 281721 229075 281779 229081
rect 281721 229041 281733 229075
rect 281767 229072 281779 229075
rect 281810 229072 281816 229084
rect 281767 229044 281816 229072
rect 281767 229041 281779 229044
rect 281721 229035 281779 229041
rect 281810 229032 281816 229044
rect 281868 229032 281874 229084
rect 332870 229032 332876 229084
rect 332928 229072 332934 229084
rect 333054 229072 333060 229084
rect 332928 229044 333060 229072
rect 332928 229032 332934 229044
rect 333054 229032 333060 229044
rect 333112 229032 333118 229084
rect 331306 227780 331312 227792
rect 331267 227752 331312 227780
rect 331306 227740 331312 227752
rect 331364 227740 331370 227792
rect 236270 225088 236276 225140
rect 236328 225088 236334 225140
rect 236288 225004 236316 225088
rect 233326 224952 233332 225004
rect 233384 224992 233390 225004
rect 233510 224992 233516 225004
rect 233384 224964 233516 224992
rect 233384 224952 233390 224964
rect 233510 224952 233516 224964
rect 233568 224952 233574 225004
rect 236270 224952 236276 225004
rect 236328 224952 236334 225004
rect 270770 224992 270776 225004
rect 270696 224964 270776 224992
rect 270696 224936 270724 224964
rect 270770 224952 270776 224964
rect 270828 224952 270834 225004
rect 347958 224952 347964 225004
rect 348016 224952 348022 225004
rect 353478 224952 353484 225004
rect 353536 224952 353542 225004
rect 381078 224952 381084 225004
rect 381136 224952 381142 225004
rect 422294 224952 422300 225004
rect 422352 224992 422358 225004
rect 422478 224992 422484 225004
rect 422352 224964 422484 224992
rect 422352 224952 422358 224964
rect 422478 224952 422484 224964
rect 422536 224952 422542 225004
rect 427814 224952 427820 225004
rect 427872 224992 427878 225004
rect 427998 224992 428004 225004
rect 427872 224964 428004 224992
rect 427872 224952 427878 224964
rect 427998 224952 428004 224964
rect 428056 224952 428062 225004
rect 451277 224995 451335 225001
rect 451277 224961 451289 224995
rect 451323 224992 451335 224995
rect 451366 224992 451372 225004
rect 451323 224964 451372 224992
rect 451323 224961 451335 224964
rect 451277 224955 451335 224961
rect 451366 224952 451372 224964
rect 451424 224952 451430 225004
rect 270678 224884 270684 224936
rect 270736 224884 270742 224936
rect 236270 224856 236276 224868
rect 236231 224828 236276 224856
rect 236270 224816 236276 224828
rect 236328 224816 236334 224868
rect 347976 224856 348004 224952
rect 348050 224856 348056 224868
rect 347976 224828 348056 224856
rect 348050 224816 348056 224828
rect 348108 224816 348114 224868
rect 353496 224856 353524 224952
rect 353570 224856 353576 224868
rect 353496 224828 353576 224856
rect 353570 224816 353576 224828
rect 353628 224816 353634 224868
rect 381096 224856 381124 224952
rect 408678 224884 408684 224936
rect 408736 224924 408742 224936
rect 408862 224924 408868 224936
rect 408736 224896 408868 224924
rect 408736 224884 408742 224896
rect 408862 224884 408868 224896
rect 408920 224884 408926 224936
rect 381170 224856 381176 224868
rect 381096 224828 381176 224856
rect 381170 224816 381176 224828
rect 381228 224816 381234 224868
rect 242802 222164 242808 222216
rect 242860 222204 242866 222216
rect 243170 222204 243176 222216
rect 242860 222176 243176 222204
rect 242860 222164 242866 222176
rect 243170 222164 243176 222176
rect 243228 222164 243234 222216
rect 252738 222164 252744 222216
rect 252796 222204 252802 222216
rect 252922 222204 252928 222216
rect 252796 222176 252928 222204
rect 252796 222164 252802 222176
rect 252922 222164 252928 222176
rect 252980 222164 252986 222216
rect 259641 222207 259699 222213
rect 259641 222173 259653 222207
rect 259687 222204 259699 222207
rect 259730 222204 259736 222216
rect 259687 222176 259736 222204
rect 259687 222173 259699 222176
rect 259641 222167 259699 222173
rect 259730 222164 259736 222176
rect 259788 222164 259794 222216
rect 295518 222164 295524 222216
rect 295576 222204 295582 222216
rect 295794 222204 295800 222216
rect 295576 222176 295800 222204
rect 295576 222164 295582 222176
rect 295794 222164 295800 222176
rect 295852 222164 295858 222216
rect 298278 222164 298284 222216
rect 298336 222204 298342 222216
rect 298554 222204 298560 222216
rect 298336 222176 298560 222204
rect 298336 222164 298342 222176
rect 298554 222164 298560 222176
rect 298612 222164 298618 222216
rect 309321 222207 309379 222213
rect 309321 222173 309333 222207
rect 309367 222204 309379 222207
rect 309502 222204 309508 222216
rect 309367 222176 309508 222204
rect 309367 222173 309379 222176
rect 309321 222167 309379 222173
rect 309502 222164 309508 222176
rect 309560 222164 309566 222216
rect 392118 222164 392124 222216
rect 392176 222204 392182 222216
rect 392302 222204 392308 222216
rect 392176 222176 392308 222204
rect 392176 222164 392182 222176
rect 392302 222164 392308 222176
rect 392360 222164 392366 222216
rect 400398 222164 400404 222216
rect 400456 222204 400462 222216
rect 400490 222204 400496 222216
rect 400456 222176 400496 222204
rect 400456 222164 400462 222176
rect 400490 222164 400496 222176
rect 400548 222164 400554 222216
rect 451274 222204 451280 222216
rect 451235 222176 451280 222204
rect 451274 222164 451280 222176
rect 451332 222164 451338 222216
rect 466546 222096 466552 222148
rect 466604 222136 466610 222148
rect 466638 222136 466644 222148
rect 466604 222108 466644 222136
rect 466604 222096 466610 222108
rect 466638 222096 466644 222108
rect 466696 222096 466702 222148
rect 243078 222068 243084 222080
rect 243039 222040 243084 222068
rect 243078 222028 243084 222040
rect 243136 222028 243142 222080
rect 292758 220912 292764 220924
rect 292684 220884 292764 220912
rect 292684 220856 292712 220884
rect 292758 220872 292764 220884
rect 292816 220872 292822 220924
rect 266722 220804 266728 220856
rect 266780 220844 266786 220856
rect 266906 220844 266912 220856
rect 266780 220816 266912 220844
rect 266780 220804 266786 220816
rect 266906 220804 266912 220816
rect 266964 220804 266970 220856
rect 292666 220804 292672 220856
rect 292724 220804 292730 220856
rect 327258 220804 327264 220856
rect 327316 220844 327322 220856
rect 327442 220844 327448 220856
rect 327316 220816 327448 220844
rect 327316 220804 327322 220816
rect 327442 220804 327448 220816
rect 327500 220804 327506 220856
rect 351822 220804 351828 220856
rect 351880 220844 351886 220856
rect 352006 220844 352012 220856
rect 351880 220816 352012 220844
rect 351880 220804 351886 220816
rect 352006 220804 352012 220816
rect 352064 220804 352070 220856
rect 358906 220804 358912 220856
rect 358964 220844 358970 220856
rect 359090 220844 359096 220856
rect 358964 220816 359096 220844
rect 358964 220804 358970 220816
rect 359090 220804 359096 220816
rect 359148 220804 359154 220856
rect 364426 220804 364432 220856
rect 364484 220844 364490 220856
rect 364702 220844 364708 220856
rect 364484 220816 364708 220844
rect 364484 220804 364490 220816
rect 364702 220804 364708 220816
rect 364760 220804 364766 220856
rect 369762 220804 369768 220856
rect 369820 220844 369826 220856
rect 369946 220844 369952 220856
rect 369820 220816 369952 220844
rect 369820 220804 369826 220816
rect 369946 220804 369952 220816
rect 370004 220804 370010 220856
rect 375466 220804 375472 220856
rect 375524 220844 375530 220856
rect 375558 220844 375564 220856
rect 375524 220816 375564 220844
rect 375524 220804 375530 220816
rect 375558 220804 375564 220816
rect 375616 220804 375622 220856
rect 287238 220668 287244 220720
rect 287296 220708 287302 220720
rect 287330 220708 287336 220720
rect 287296 220680 287336 220708
rect 287296 220668 287302 220680
rect 287330 220668 287336 220680
rect 287388 220668 287394 220720
rect 375466 220668 375472 220720
rect 375524 220708 375530 220720
rect 375834 220708 375840 220720
rect 375524 220680 375840 220708
rect 375524 220668 375530 220680
rect 375834 220668 375840 220680
rect 375892 220668 375898 220720
rect 334342 219416 334348 219428
rect 334303 219388 334348 219416
rect 334342 219376 334348 219388
rect 334400 219376 334406 219428
rect 358906 217948 358912 218000
rect 358964 217988 358970 218000
rect 358998 217988 359004 218000
rect 358964 217960 359004 217988
rect 358964 217948 358970 217960
rect 358998 217948 359004 217960
rect 359056 217948 359062 218000
rect 259730 217444 259736 217456
rect 259656 217416 259736 217444
rect 259656 217388 259684 217416
rect 259730 217404 259736 217416
rect 259788 217404 259794 217456
rect 259638 217336 259644 217388
rect 259696 217336 259702 217388
rect 231854 216588 231860 216640
rect 231912 216628 231918 216640
rect 232038 216628 232044 216640
rect 231912 216600 232044 216628
rect 231912 216588 231918 216600
rect 232038 216588 232044 216600
rect 232096 216588 232102 216640
rect 321738 215976 321744 216028
rect 321796 216016 321802 216028
rect 321922 216016 321928 216028
rect 321796 215988 321928 216016
rect 321796 215976 321802 215988
rect 321922 215976 321928 215988
rect 321980 215976 321986 216028
rect 324498 215976 324504 216028
rect 324556 216016 324562 216028
rect 324682 216016 324688 216028
rect 324556 215988 324688 216016
rect 324556 215976 324562 215988
rect 324682 215976 324688 215988
rect 324740 215976 324746 216028
rect 270678 215404 270684 215416
rect 270639 215376 270684 215404
rect 270678 215364 270684 215376
rect 270736 215364 270742 215416
rect 236270 215336 236276 215348
rect 236231 215308 236276 215336
rect 236270 215296 236276 215308
rect 236328 215296 236334 215348
rect 255590 215336 255596 215348
rect 255516 215308 255596 215336
rect 255516 215280 255544 215308
rect 255590 215296 255596 215308
rect 255648 215296 255654 215348
rect 261110 215336 261116 215348
rect 261036 215308 261116 215336
rect 261036 215280 261064 215308
rect 261110 215296 261116 215308
rect 261168 215296 261174 215348
rect 330110 215336 330116 215348
rect 330036 215308 330116 215336
rect 330036 215280 330064 215308
rect 330110 215296 330116 215308
rect 330168 215296 330174 215348
rect 357710 215336 357716 215348
rect 357636 215308 357716 215336
rect 357636 215280 357664 215308
rect 357710 215296 357716 215308
rect 357768 215296 357774 215348
rect 367462 215336 367468 215348
rect 367388 215308 367468 215336
rect 367388 215280 367416 215308
rect 367462 215296 367468 215308
rect 367520 215296 367526 215348
rect 408770 215336 408776 215348
rect 408731 215308 408776 215336
rect 408770 215296 408776 215308
rect 408828 215296 408834 215348
rect 255498 215228 255504 215280
rect 255556 215228 255562 215280
rect 261018 215228 261024 215280
rect 261076 215228 261082 215280
rect 283098 215228 283104 215280
rect 283156 215228 283162 215280
rect 330018 215228 330024 215280
rect 330076 215228 330082 215280
rect 357618 215228 357624 215280
rect 357676 215228 357682 215280
rect 367370 215228 367376 215280
rect 367428 215228 367434 215280
rect 376938 215228 376944 215280
rect 376996 215228 377002 215280
rect 387978 215228 387984 215280
rect 388036 215228 388042 215280
rect 283116 215144 283144 215228
rect 376956 215144 376984 215228
rect 387996 215144 388024 215228
rect 283098 215092 283104 215144
rect 283156 215092 283162 215144
rect 376938 215092 376944 215144
rect 376996 215092 377002 215144
rect 387978 215092 387984 215144
rect 388036 215092 388042 215144
rect 364334 212780 364340 212832
rect 364392 212820 364398 212832
rect 364392 212792 364437 212820
rect 364392 212780 364398 212792
rect 265158 212644 265164 212696
rect 265216 212684 265222 212696
rect 265216 212656 265296 212684
rect 265216 212644 265222 212656
rect 254210 212616 254216 212628
rect 254136 212588 254216 212616
rect 254136 212560 254164 212588
rect 254210 212576 254216 212588
rect 254268 212576 254274 212628
rect 265268 212560 265296 212656
rect 356514 212616 356520 212628
rect 356440 212588 356520 212616
rect 356440 212560 356468 212588
rect 356514 212576 356520 212588
rect 356572 212576 356578 212628
rect 243081 212551 243139 212557
rect 243081 212517 243093 212551
rect 243127 212548 243139 212551
rect 243170 212548 243176 212560
rect 243127 212520 243176 212548
rect 243127 212517 243139 212520
rect 243081 212511 243139 212517
rect 243170 212508 243176 212520
rect 243228 212508 243234 212560
rect 252738 212508 252744 212560
rect 252796 212548 252802 212560
rect 252830 212548 252836 212560
rect 252796 212520 252836 212548
rect 252796 212508 252802 212520
rect 252830 212508 252836 212520
rect 252888 212508 252894 212560
rect 254118 212508 254124 212560
rect 254176 212508 254182 212560
rect 265250 212508 265256 212560
rect 265308 212508 265314 212560
rect 271874 212508 271880 212560
rect 271932 212548 271938 212560
rect 272058 212548 272064 212560
rect 271932 212520 272064 212548
rect 271932 212508 271938 212520
rect 272058 212508 272064 212520
rect 272116 212508 272122 212560
rect 277578 212508 277584 212560
rect 277636 212548 277642 212560
rect 277670 212548 277676 212560
rect 277636 212520 277676 212548
rect 277636 212508 277642 212520
rect 277670 212508 277676 212520
rect 277728 212508 277734 212560
rect 288434 212508 288440 212560
rect 288492 212548 288498 212560
rect 288618 212548 288624 212560
rect 288492 212520 288624 212548
rect 288492 212508 288498 212520
rect 288618 212508 288624 212520
rect 288676 212508 288682 212560
rect 298278 212508 298284 212560
rect 298336 212548 298342 212560
rect 298554 212548 298560 212560
rect 298336 212520 298560 212548
rect 298336 212508 298342 212520
rect 298554 212508 298560 212520
rect 298612 212508 298618 212560
rect 305178 212508 305184 212560
rect 305236 212548 305242 212560
rect 305362 212548 305368 212560
rect 305236 212520 305368 212548
rect 305236 212508 305242 212520
rect 305362 212508 305368 212520
rect 305420 212508 305426 212560
rect 308122 212508 308128 212560
rect 308180 212548 308186 212560
rect 308306 212548 308312 212560
rect 308180 212520 308312 212548
rect 308180 212508 308186 212520
rect 308306 212508 308312 212520
rect 308364 212508 308370 212560
rect 310698 212508 310704 212560
rect 310756 212548 310762 212560
rect 310882 212548 310888 212560
rect 310756 212520 310888 212548
rect 310756 212508 310762 212520
rect 310882 212508 310888 212520
rect 310940 212508 310946 212560
rect 318978 212508 318984 212560
rect 319036 212548 319042 212560
rect 319070 212548 319076 212560
rect 319036 212520 319076 212548
rect 319036 212508 319042 212520
rect 319070 212508 319076 212520
rect 319128 212508 319134 212560
rect 346578 212508 346584 212560
rect 346636 212548 346642 212560
rect 346762 212548 346768 212560
rect 346636 212520 346768 212548
rect 346636 212508 346642 212520
rect 346762 212508 346768 212520
rect 346820 212508 346826 212560
rect 347958 212508 347964 212560
rect 348016 212548 348022 212560
rect 348142 212548 348148 212560
rect 348016 212520 348148 212548
rect 348016 212508 348022 212520
rect 348142 212508 348148 212520
rect 348200 212508 348206 212560
rect 352006 212508 352012 212560
rect 352064 212548 352070 212560
rect 352098 212548 352104 212560
rect 352064 212520 352104 212548
rect 352064 212508 352070 212520
rect 352098 212508 352104 212520
rect 352156 212508 352162 212560
rect 353478 212508 353484 212560
rect 353536 212548 353542 212560
rect 353662 212548 353668 212560
rect 353536 212520 353668 212548
rect 353536 212508 353542 212520
rect 353662 212508 353668 212520
rect 353720 212508 353726 212560
rect 356422 212508 356428 212560
rect 356480 212508 356486 212560
rect 364153 212551 364211 212557
rect 364153 212517 364165 212551
rect 364199 212548 364211 212551
rect 364426 212548 364432 212560
rect 364199 212520 364432 212548
rect 364199 212517 364211 212520
rect 364153 212511 364211 212517
rect 364426 212508 364432 212520
rect 364484 212508 364490 212560
rect 382274 212508 382280 212560
rect 382332 212548 382338 212560
rect 382458 212548 382464 212560
rect 382332 212520 382464 212548
rect 382332 212508 382338 212520
rect 382458 212508 382464 212520
rect 382516 212508 382522 212560
rect 386598 212508 386604 212560
rect 386656 212548 386662 212560
rect 386874 212548 386880 212560
rect 386656 212520 386880 212548
rect 386656 212508 386662 212520
rect 386874 212508 386880 212520
rect 386932 212508 386938 212560
rect 400306 212508 400312 212560
rect 400364 212548 400370 212560
rect 400582 212548 400588 212560
rect 400364 212520 400588 212548
rect 400364 212508 400370 212520
rect 400582 212508 400588 212520
rect 400640 212508 400646 212560
rect 408770 212548 408776 212560
rect 408731 212520 408776 212548
rect 408770 212508 408776 212520
rect 408828 212508 408834 212560
rect 416958 212508 416964 212560
rect 417016 212548 417022 212560
rect 417142 212548 417148 212560
rect 417016 212520 417148 212548
rect 417016 212508 417022 212520
rect 417142 212508 417148 212520
rect 417200 212508 417206 212560
rect 433426 212508 433432 212560
rect 433484 212548 433490 212560
rect 433702 212548 433708 212560
rect 433484 212520 433708 212548
rect 433484 212508 433490 212520
rect 433702 212508 433708 212520
rect 433760 212508 433766 212560
rect 472158 212508 472164 212560
rect 472216 212548 472222 212560
rect 472342 212548 472348 212560
rect 472216 212520 472348 212548
rect 472216 212508 472222 212520
rect 472342 212508 472348 212520
rect 472400 212508 472406 212560
rect 259638 212480 259644 212492
rect 259599 212452 259644 212480
rect 259638 212440 259644 212452
rect 259696 212440 259702 212492
rect 270678 212480 270684 212492
rect 270639 212452 270684 212480
rect 270678 212440 270684 212452
rect 270736 212440 270742 212492
rect 281721 212483 281779 212489
rect 281721 212449 281733 212483
rect 281767 212480 281779 212483
rect 281810 212480 281816 212492
rect 281767 212452 281816 212480
rect 281767 212449 281779 212452
rect 281721 212443 281779 212449
rect 281810 212440 281816 212452
rect 281868 212440 281874 212492
rect 334345 212483 334403 212489
rect 334345 212449 334357 212483
rect 334391 212480 334403 212483
rect 334434 212480 334440 212492
rect 334391 212452 334440 212480
rect 334391 212449 334403 212452
rect 334345 212443 334403 212449
rect 334434 212440 334440 212452
rect 334492 212440 334498 212492
rect 369946 212480 369952 212492
rect 369907 212452 369952 212480
rect 369946 212440 369952 212452
rect 370004 212440 370010 212492
rect 364334 212372 364340 212424
rect 364392 212412 364398 212424
rect 364392 212384 364437 212412
rect 364392 212372 364398 212384
rect 292666 211148 292672 211200
rect 292724 211188 292730 211200
rect 292758 211188 292764 211200
rect 292724 211160 292764 211188
rect 292724 211148 292730 211160
rect 292758 211148 292764 211160
rect 292816 211148 292822 211200
rect 255314 211080 255320 211132
rect 255372 211120 255378 211132
rect 255498 211120 255504 211132
rect 255372 211092 255504 211120
rect 255372 211080 255378 211092
rect 255498 211080 255504 211092
rect 255556 211080 255562 211132
rect 270678 211120 270684 211132
rect 270639 211092 270684 211120
rect 270678 211080 270684 211092
rect 270736 211080 270742 211132
rect 351822 211080 351828 211132
rect 351880 211120 351886 211132
rect 352006 211120 352012 211132
rect 351880 211092 352012 211120
rect 351880 211080 351886 211092
rect 352006 211080 352012 211092
rect 352064 211080 352070 211132
rect 295518 209760 295524 209772
rect 295479 209732 295524 209760
rect 295518 209720 295524 209732
rect 295576 209720 295582 209772
rect 331122 209720 331128 209772
rect 331180 209760 331186 209772
rect 331306 209760 331312 209772
rect 331180 209732 331312 209760
rect 331180 209720 331186 209732
rect 331306 209720 331312 209732
rect 331364 209720 331370 209772
rect 332686 209720 332692 209772
rect 332744 209760 332750 209772
rect 332870 209760 332876 209772
rect 332744 209732 332876 209760
rect 332744 209720 332750 209732
rect 332870 209720 332876 209732
rect 332928 209720 332934 209772
rect 386598 209720 386604 209772
rect 386656 209760 386662 209772
rect 386782 209760 386788 209772
rect 386656 209732 386788 209760
rect 386656 209720 386662 209732
rect 386782 209720 386788 209732
rect 386840 209720 386846 209772
rect 364150 208400 364156 208412
rect 364111 208372 364156 208400
rect 364150 208360 364156 208372
rect 364208 208360 364214 208412
rect 236362 207000 236368 207052
rect 236420 207040 236426 207052
rect 236420 207012 236684 207040
rect 236420 207000 236426 207012
rect 236656 206916 236684 207012
rect 236638 206864 236644 206916
rect 236696 206864 236702 206916
rect 233326 205640 233332 205692
rect 233384 205680 233390 205692
rect 233510 205680 233516 205692
rect 233384 205652 233516 205680
rect 233384 205640 233390 205652
rect 233510 205640 233516 205652
rect 233568 205640 233574 205692
rect 243170 205680 243176 205692
rect 243131 205652 243176 205680
rect 243170 205640 243176 205652
rect 243228 205640 243234 205692
rect 265250 205680 265256 205692
rect 265211 205652 265256 205680
rect 265250 205640 265256 205652
rect 265308 205640 265314 205692
rect 292758 205640 292764 205692
rect 292816 205640 292822 205692
rect 298278 205640 298284 205692
rect 298336 205640 298342 205692
rect 336826 205680 336832 205692
rect 336787 205652 336832 205680
rect 336826 205640 336832 205652
rect 336884 205640 336890 205692
rect 347958 205640 347964 205692
rect 348016 205640 348022 205692
rect 422294 205640 422300 205692
rect 422352 205680 422358 205692
rect 422478 205680 422484 205692
rect 422352 205652 422484 205680
rect 422352 205640 422358 205652
rect 422478 205640 422484 205652
rect 422536 205640 422542 205692
rect 427814 205640 427820 205692
rect 427872 205680 427878 205692
rect 427998 205680 428004 205692
rect 427872 205652 428004 205680
rect 427872 205640 427878 205652
rect 427998 205640 428004 205652
rect 428056 205640 428062 205692
rect 270678 205612 270684 205624
rect 270639 205584 270684 205612
rect 270678 205572 270684 205584
rect 270736 205572 270742 205624
rect 292776 205544 292804 205640
rect 298296 205612 298324 205640
rect 298370 205612 298376 205624
rect 298296 205584 298376 205612
rect 298370 205572 298376 205584
rect 298428 205572 298434 205624
rect 347976 205612 348004 205640
rect 348050 205612 348056 205624
rect 347976 205584 348056 205612
rect 348050 205572 348056 205584
rect 348108 205572 348114 205624
rect 292850 205544 292856 205556
rect 292776 205516 292856 205544
rect 292850 205504 292856 205516
rect 292908 205504 292914 205556
rect 336734 204348 336740 204400
rect 336792 204388 336798 204400
rect 338114 204388 338120 204400
rect 336792 204360 338120 204388
rect 336792 204348 336798 204360
rect 338114 204348 338120 204360
rect 338172 204348 338178 204400
rect 375190 204348 375196 204400
rect 375248 204388 375254 204400
rect 384942 204388 384948 204400
rect 375248 204360 384948 204388
rect 375248 204348 375254 204360
rect 384942 204348 384948 204360
rect 385000 204348 385006 204400
rect 425054 204348 425060 204400
rect 425112 204388 425118 204400
rect 434530 204388 434536 204400
rect 425112 204360 434536 204388
rect 425112 204348 425118 204360
rect 434530 204348 434536 204360
rect 434588 204348 434594 204400
rect 521654 204348 521660 204400
rect 521712 204388 521718 204400
rect 526438 204388 526444 204400
rect 521712 204360 526444 204388
rect 521712 204348 521718 204360
rect 526438 204348 526444 204360
rect 526496 204348 526502 204400
rect 309318 202920 309324 202972
rect 309376 202960 309382 202972
rect 309410 202960 309416 202972
rect 309376 202932 309416 202960
rect 309376 202920 309382 202932
rect 309410 202920 309416 202932
rect 309468 202920 309474 202972
rect 480257 202963 480315 202969
rect 480257 202929 480269 202963
rect 480303 202960 480315 202963
rect 480346 202960 480352 202972
rect 480303 202932 480352 202960
rect 480303 202929 480315 202932
rect 480257 202923 480315 202929
rect 480346 202920 480352 202932
rect 480404 202920 480410 202972
rect 243170 202892 243176 202904
rect 243131 202864 243176 202892
rect 243170 202852 243176 202864
rect 243228 202852 243234 202904
rect 259641 202895 259699 202901
rect 259641 202861 259653 202895
rect 259687 202892 259699 202895
rect 259730 202892 259736 202904
rect 259687 202864 259736 202892
rect 259687 202861 259699 202864
rect 259641 202855 259699 202861
rect 259730 202852 259736 202864
rect 259788 202852 259794 202904
rect 265250 202892 265256 202904
rect 265211 202864 265256 202892
rect 265250 202852 265256 202864
rect 265308 202852 265314 202904
rect 281718 202852 281724 202904
rect 281776 202892 281782 202904
rect 281902 202892 281908 202904
rect 281776 202864 281908 202892
rect 281776 202852 281782 202864
rect 281902 202852 281908 202864
rect 281960 202852 281966 202904
rect 327258 202852 327264 202904
rect 327316 202892 327322 202904
rect 327350 202892 327356 202904
rect 327316 202864 327356 202892
rect 327316 202852 327322 202864
rect 327350 202852 327356 202864
rect 327408 202852 327414 202904
rect 336826 202892 336832 202904
rect 336787 202864 336832 202892
rect 336826 202852 336832 202864
rect 336884 202852 336890 202904
rect 364150 202852 364156 202904
rect 364208 202892 364214 202904
rect 364610 202892 364616 202904
rect 364208 202864 364616 202892
rect 364208 202852 364214 202864
rect 364610 202852 364616 202864
rect 364668 202852 364674 202904
rect 369946 202892 369952 202904
rect 369907 202864 369952 202892
rect 369946 202852 369952 202864
rect 370004 202852 370010 202904
rect 295518 202824 295524 202836
rect 295479 202796 295524 202824
rect 295518 202784 295524 202796
rect 295576 202784 295582 202836
rect 318978 202784 318984 202836
rect 319036 202824 319042 202836
rect 319070 202824 319076 202836
rect 319036 202796 319076 202824
rect 319036 202784 319042 202796
rect 319070 202784 319076 202796
rect 319128 202784 319134 202836
rect 400490 202784 400496 202836
rect 400548 202824 400554 202836
rect 400582 202824 400588 202836
rect 400548 202796 400588 202824
rect 400548 202784 400554 202796
rect 400582 202784 400588 202796
rect 400640 202784 400646 202836
rect 243078 202756 243084 202768
rect 243039 202728 243084 202756
rect 243078 202716 243084 202728
rect 243136 202716 243142 202768
rect 480254 201532 480260 201544
rect 480215 201504 480260 201532
rect 480254 201492 480260 201504
rect 480312 201492 480318 201544
rect 255498 201424 255504 201476
rect 255556 201464 255562 201476
rect 255590 201464 255596 201476
rect 255556 201436 255596 201464
rect 255556 201424 255562 201436
rect 255590 201424 255596 201436
rect 255648 201424 255654 201476
rect 281902 201464 281908 201476
rect 281863 201436 281908 201464
rect 281902 201424 281908 201436
rect 281960 201424 281966 201476
rect 287330 201424 287336 201476
rect 287388 201464 287394 201476
rect 309321 201467 309379 201473
rect 287388 201436 287468 201464
rect 287388 201424 287394 201436
rect 287440 201408 287468 201436
rect 309321 201433 309333 201467
rect 309367 201464 309379 201467
rect 309410 201464 309416 201476
rect 309367 201436 309416 201464
rect 309367 201433 309379 201436
rect 309321 201427 309379 201433
rect 309410 201424 309416 201436
rect 309468 201424 309474 201476
rect 321738 201424 321744 201476
rect 321796 201464 321802 201476
rect 321922 201464 321928 201476
rect 321796 201436 321928 201464
rect 321796 201424 321802 201436
rect 321922 201424 321928 201436
rect 321980 201424 321986 201476
rect 324498 201424 324504 201476
rect 324556 201464 324562 201476
rect 324682 201464 324688 201476
rect 324556 201436 324688 201464
rect 324556 201424 324562 201436
rect 324682 201424 324688 201436
rect 324740 201424 324746 201476
rect 352098 201464 352104 201476
rect 352059 201436 352104 201464
rect 352098 201424 352104 201436
rect 352156 201424 352162 201476
rect 369946 201464 369952 201476
rect 369907 201436 369952 201464
rect 369946 201424 369952 201436
rect 370004 201424 370010 201476
rect 287422 201356 287428 201408
rect 287480 201356 287486 201408
rect 255498 200104 255504 200116
rect 255459 200076 255504 200104
rect 255498 200064 255504 200076
rect 255556 200064 255562 200116
rect 294138 200064 294144 200116
rect 294196 200104 294202 200116
rect 294230 200104 294236 200116
rect 294196 200076 294236 200104
rect 294196 200064 294202 200076
rect 294230 200064 294236 200076
rect 294288 200064 294294 200116
rect 295518 200064 295524 200116
rect 295576 200104 295582 200116
rect 295705 200107 295763 200113
rect 295705 200104 295717 200107
rect 295576 200076 295717 200104
rect 295576 200064 295582 200076
rect 295705 200073 295717 200076
rect 295751 200073 295763 200107
rect 295705 200067 295763 200073
rect 386598 200064 386604 200116
rect 386656 200104 386662 200116
rect 386874 200104 386880 200116
rect 386656 200076 386880 200104
rect 386656 200064 386662 200076
rect 386874 200064 386880 200076
rect 386932 200064 386938 200116
rect 332778 198676 332784 198688
rect 332739 198648 332784 198676
rect 332778 198636 332784 198648
rect 332836 198636 332842 198688
rect 386598 198676 386604 198688
rect 386559 198648 386604 198676
rect 386598 198636 386604 198648
rect 386656 198636 386662 198688
rect 236454 198568 236460 198620
rect 236512 198608 236518 198620
rect 236638 198608 236644 198620
rect 236512 198580 236644 198608
rect 236512 198568 236518 198580
rect 236638 198568 236644 198580
rect 236696 198568 236702 198620
rect 259730 198132 259736 198144
rect 259656 198104 259736 198132
rect 259656 198076 259684 198104
rect 259730 198092 259736 198104
rect 259788 198092 259794 198144
rect 259638 198024 259644 198076
rect 259696 198024 259702 198076
rect 359090 197276 359096 197328
rect 359148 197316 359154 197328
rect 359185 197319 359243 197325
rect 359185 197316 359197 197319
rect 359148 197288 359197 197316
rect 359148 197276 359154 197288
rect 359185 197285 359197 197288
rect 359231 197285 359243 197319
rect 359185 197279 359243 197285
rect 342714 196596 342720 196648
rect 342772 196636 342778 196648
rect 342898 196636 342904 196648
rect 342772 196608 342904 196636
rect 342772 196596 342778 196608
rect 342898 196596 342904 196608
rect 342956 196596 342962 196648
rect 365714 196596 365720 196648
rect 365772 196636 365778 196648
rect 365898 196636 365904 196648
rect 365772 196608 365904 196636
rect 365772 196596 365778 196608
rect 365898 196596 365904 196608
rect 365956 196596 365962 196648
rect 270589 196095 270647 196101
rect 270589 196061 270601 196095
rect 270635 196092 270647 196095
rect 270770 196092 270776 196104
rect 270635 196064 270776 196092
rect 270635 196061 270647 196064
rect 270589 196055 270647 196061
rect 270770 196052 270776 196064
rect 270828 196052 270834 196104
rect 364610 196052 364616 196104
rect 364668 196092 364674 196104
rect 364794 196092 364800 196104
rect 364668 196064 364800 196092
rect 364668 196052 364674 196064
rect 364794 196052 364800 196064
rect 364852 196052 364858 196104
rect 375561 196095 375619 196101
rect 375561 196061 375573 196095
rect 375607 196092 375619 196095
rect 375650 196092 375656 196104
rect 375607 196064 375656 196092
rect 375607 196061 375619 196064
rect 375561 196055 375619 196061
rect 375650 196052 375656 196064
rect 375708 196052 375714 196104
rect 433702 196092 433708 196104
rect 433663 196064 433708 196092
rect 433702 196052 433708 196064
rect 433760 196052 433766 196104
rect 367462 196024 367468 196036
rect 367388 195996 367468 196024
rect 367388 195968 367416 195996
rect 367462 195984 367468 195996
rect 367520 195984 367526 196036
rect 480254 195984 480260 196036
rect 480312 195984 480318 196036
rect 277486 195916 277492 195968
rect 277544 195956 277550 195968
rect 277670 195956 277676 195968
rect 277544 195928 277676 195956
rect 277544 195916 277550 195928
rect 277670 195916 277676 195928
rect 277728 195916 277734 195968
rect 367370 195916 367376 195968
rect 367428 195916 367434 195968
rect 376938 195916 376944 195968
rect 376996 195916 377002 195968
rect 387978 195916 387984 195968
rect 388036 195916 388042 195968
rect 376956 195832 376984 195916
rect 387996 195832 388024 195916
rect 480272 195888 480300 195984
rect 480346 195888 480352 195900
rect 480272 195860 480352 195888
rect 480346 195848 480352 195860
rect 480404 195848 480410 195900
rect 376938 195780 376944 195832
rect 376996 195780 377002 195832
rect 387978 195780 387984 195832
rect 388036 195780 388042 195832
rect 265250 193304 265256 193316
rect 265176 193276 265256 193304
rect 265176 193248 265204 193276
rect 265250 193264 265256 193276
rect 265308 193264 265314 193316
rect 356514 193304 356520 193316
rect 356440 193276 356520 193304
rect 356440 193248 356468 193276
rect 356514 193264 356520 193276
rect 356572 193264 356578 193316
rect 243081 193239 243139 193245
rect 243081 193205 243093 193239
rect 243127 193236 243139 193239
rect 243170 193236 243176 193248
rect 243127 193208 243176 193236
rect 243127 193205 243139 193208
rect 243081 193199 243139 193205
rect 243170 193196 243176 193208
rect 243228 193196 243234 193248
rect 252830 193196 252836 193248
rect 252888 193236 252894 193248
rect 253014 193236 253020 193248
rect 252888 193208 253020 193236
rect 252888 193196 252894 193208
rect 253014 193196 253020 193208
rect 253072 193196 253078 193248
rect 265158 193196 265164 193248
rect 265216 193196 265222 193248
rect 266998 193196 267004 193248
rect 267056 193236 267062 193248
rect 267090 193236 267096 193248
rect 267056 193208 267096 193236
rect 267056 193196 267062 193208
rect 267090 193196 267096 193208
rect 267148 193196 267154 193248
rect 288434 193196 288440 193248
rect 288492 193236 288498 193248
rect 288618 193236 288624 193248
rect 288492 193208 288624 193236
rect 288492 193196 288498 193208
rect 288618 193196 288624 193208
rect 288676 193196 288682 193248
rect 292758 193196 292764 193248
rect 292816 193236 292822 193248
rect 292942 193236 292948 193248
rect 292816 193208 292948 193236
rect 292816 193196 292822 193208
rect 292942 193196 292948 193208
rect 293000 193196 293006 193248
rect 298278 193196 298284 193248
rect 298336 193236 298342 193248
rect 298462 193236 298468 193248
rect 298336 193208 298468 193236
rect 298336 193196 298342 193208
rect 298462 193196 298468 193208
rect 298520 193196 298526 193248
rect 305178 193196 305184 193248
rect 305236 193236 305242 193248
rect 305362 193236 305368 193248
rect 305236 193208 305368 193236
rect 305236 193196 305242 193208
rect 305362 193196 305368 193208
rect 305420 193196 305426 193248
rect 308122 193196 308128 193248
rect 308180 193236 308186 193248
rect 308306 193236 308312 193248
rect 308180 193208 308312 193236
rect 308180 193196 308186 193208
rect 308306 193196 308312 193208
rect 308364 193196 308370 193248
rect 327258 193196 327264 193248
rect 327316 193236 327322 193248
rect 327350 193236 327356 193248
rect 327316 193208 327356 193236
rect 327316 193196 327322 193208
rect 327350 193196 327356 193208
rect 327408 193196 327414 193248
rect 330018 193196 330024 193248
rect 330076 193196 330082 193248
rect 334342 193196 334348 193248
rect 334400 193236 334406 193248
rect 334434 193236 334440 193248
rect 334400 193208 334440 193236
rect 334400 193196 334406 193208
rect 334434 193196 334440 193208
rect 334492 193196 334498 193248
rect 336734 193196 336740 193248
rect 336792 193236 336798 193248
rect 336826 193236 336832 193248
rect 336792 193208 336832 193236
rect 336792 193196 336798 193208
rect 336826 193196 336832 193208
rect 336884 193196 336890 193248
rect 346578 193196 346584 193248
rect 346636 193236 346642 193248
rect 346762 193236 346768 193248
rect 346636 193208 346768 193236
rect 346636 193196 346642 193208
rect 346762 193196 346768 193208
rect 346820 193196 346826 193248
rect 347958 193196 347964 193248
rect 348016 193236 348022 193248
rect 348142 193236 348148 193248
rect 348016 193208 348148 193236
rect 348016 193196 348022 193208
rect 348142 193196 348148 193208
rect 348200 193196 348206 193248
rect 353478 193196 353484 193248
rect 353536 193236 353542 193248
rect 353662 193236 353668 193248
rect 353536 193208 353668 193236
rect 353536 193196 353542 193208
rect 353662 193196 353668 193208
rect 353720 193196 353726 193248
rect 356422 193196 356428 193248
rect 356480 193196 356486 193248
rect 375558 193236 375564 193248
rect 375519 193208 375564 193236
rect 375558 193196 375564 193208
rect 375616 193196 375622 193248
rect 382274 193196 382280 193248
rect 382332 193236 382338 193248
rect 382458 193236 382464 193248
rect 382332 193208 382464 193236
rect 382332 193196 382338 193208
rect 382458 193196 382464 193208
rect 382516 193196 382522 193248
rect 392118 193196 392124 193248
rect 392176 193236 392182 193248
rect 392210 193236 392216 193248
rect 392176 193208 392216 193236
rect 392176 193196 392182 193208
rect 392210 193196 392216 193208
rect 392268 193196 392274 193248
rect 397730 193196 397736 193248
rect 397788 193236 397794 193248
rect 397914 193236 397920 193248
rect 397788 193208 397920 193236
rect 397788 193196 397794 193208
rect 397914 193196 397920 193208
rect 397972 193196 397978 193248
rect 408770 193196 408776 193248
rect 408828 193236 408834 193248
rect 408954 193236 408960 193248
rect 408828 193208 408960 193236
rect 408828 193196 408834 193208
rect 408954 193196 408960 193208
rect 409012 193196 409018 193248
rect 416958 193196 416964 193248
rect 417016 193236 417022 193248
rect 417142 193236 417148 193248
rect 417016 193208 417148 193236
rect 417016 193196 417022 193208
rect 417142 193196 417148 193208
rect 417200 193196 417206 193248
rect 433702 193236 433708 193248
rect 433663 193208 433708 193236
rect 433702 193196 433708 193208
rect 433760 193196 433766 193248
rect 472158 193196 472164 193248
rect 472216 193236 472222 193248
rect 472342 193236 472348 193248
rect 472216 193208 472348 193236
rect 472216 193196 472222 193208
rect 472342 193196 472348 193208
rect 472400 193196 472406 193248
rect 270586 193168 270592 193180
rect 270547 193140 270592 193168
rect 270586 193128 270592 193140
rect 270644 193128 270650 193180
rect 281902 193168 281908 193180
rect 281863 193140 281908 193168
rect 281902 193128 281908 193140
rect 281960 193128 281966 193180
rect 330036 193168 330064 193196
rect 330110 193168 330116 193180
rect 330036 193140 330116 193168
rect 330110 193128 330116 193140
rect 330168 193128 330174 193180
rect 352098 193168 352104 193180
rect 352059 193140 352104 193168
rect 352098 193128 352104 193140
rect 352156 193128 352162 193180
rect 369946 193168 369952 193180
rect 369907 193140 369952 193168
rect 369946 193128 369952 193140
rect 370004 193128 370010 193180
rect 231946 191768 231952 191820
rect 232004 191808 232010 191820
rect 232038 191808 232044 191820
rect 232004 191780 232044 191808
rect 232004 191768 232010 191780
rect 232038 191768 232044 191780
rect 232096 191768 232102 191820
rect 270586 191808 270592 191820
rect 270547 191780 270592 191808
rect 270586 191768 270592 191780
rect 270644 191768 270650 191820
rect 255498 190516 255504 190528
rect 255459 190488 255504 190516
rect 255498 190476 255504 190488
rect 255556 190476 255562 190528
rect 364518 190448 364524 190460
rect 364479 190420 364524 190448
rect 364518 190408 364524 190420
rect 364576 190408 364582 190460
rect 332778 189088 332784 189100
rect 332739 189060 332784 189088
rect 332778 189048 332784 189060
rect 332836 189048 332842 189100
rect 236270 187688 236276 187740
rect 236328 187728 236334 187740
rect 236454 187728 236460 187740
rect 236328 187700 236460 187728
rect 236328 187688 236334 187700
rect 236454 187688 236460 187700
rect 236512 187688 236518 187740
rect 359090 187688 359096 187740
rect 359148 187728 359154 187740
rect 359185 187731 359243 187737
rect 359185 187728 359197 187731
rect 359148 187700 359197 187728
rect 359148 187688 359154 187700
rect 359185 187697 359197 187700
rect 359231 187697 359243 187731
rect 359185 187691 359243 187697
rect 236270 187592 236276 187604
rect 236231 187564 236276 187592
rect 236270 187552 236276 187564
rect 236328 187552 236334 187604
rect 451642 186464 451648 186516
rect 451700 186464 451706 186516
rect 271969 186439 272027 186445
rect 271969 186405 271981 186439
rect 272015 186436 272027 186439
rect 272058 186436 272064 186448
rect 272015 186408 272064 186436
rect 272015 186405 272027 186408
rect 271969 186399 272027 186405
rect 272058 186396 272064 186408
rect 272116 186396 272122 186448
rect 277670 186396 277676 186448
rect 277728 186396 277734 186448
rect 298278 186436 298284 186448
rect 298239 186408 298284 186436
rect 298278 186396 298284 186408
rect 298336 186396 298342 186448
rect 321649 186439 321707 186445
rect 321649 186405 321661 186439
rect 321695 186436 321707 186439
rect 321738 186436 321744 186448
rect 321695 186408 321744 186436
rect 321695 186405 321707 186408
rect 321649 186399 321707 186405
rect 321738 186396 321744 186408
rect 321796 186396 321802 186448
rect 324409 186439 324467 186445
rect 324409 186405 324421 186439
rect 324455 186436 324467 186439
rect 324498 186436 324504 186448
rect 324455 186408 324504 186436
rect 324455 186405 324467 186408
rect 324409 186399 324467 186405
rect 324498 186396 324504 186408
rect 324556 186396 324562 186448
rect 327258 186436 327264 186448
rect 327184 186408 327264 186436
rect 233326 186328 233332 186380
rect 233384 186368 233390 186380
rect 233510 186368 233516 186380
rect 233384 186340 233516 186368
rect 233384 186328 233390 186340
rect 233510 186328 233516 186340
rect 233568 186328 233574 186380
rect 243170 186368 243176 186380
rect 243096 186340 243176 186368
rect 243096 186312 243124 186340
rect 243170 186328 243176 186340
rect 243228 186328 243234 186380
rect 243078 186260 243084 186312
rect 243136 186260 243142 186312
rect 277688 186244 277716 186396
rect 327184 186312 327212 186408
rect 327258 186396 327264 186408
rect 327316 186396 327322 186448
rect 357618 186436 357624 186448
rect 357579 186408 357624 186436
rect 357618 186396 357624 186408
rect 357676 186396 357682 186448
rect 451660 186380 451688 186464
rect 422294 186328 422300 186380
rect 422352 186368 422358 186380
rect 422478 186368 422484 186380
rect 422352 186340 422484 186368
rect 422352 186328 422358 186340
rect 422478 186328 422484 186340
rect 422536 186328 422542 186380
rect 427814 186328 427820 186380
rect 427872 186368 427878 186380
rect 427998 186368 428004 186380
rect 427872 186340 428004 186368
rect 427872 186328 427878 186340
rect 427998 186328 428004 186340
rect 428056 186328 428062 186380
rect 451642 186328 451648 186380
rect 451700 186328 451706 186380
rect 327166 186260 327172 186312
rect 327224 186260 327230 186312
rect 364518 186300 364524 186312
rect 364479 186272 364524 186300
rect 364518 186260 364524 186272
rect 364576 186260 364582 186312
rect 386598 186300 386604 186312
rect 386559 186272 386604 186300
rect 386598 186260 386604 186272
rect 386656 186260 386662 186312
rect 277670 186192 277676 186244
rect 277728 186192 277734 186244
rect 382458 183608 382464 183660
rect 382516 183608 382522 183660
rect 252830 183540 252836 183592
rect 252888 183580 252894 183592
rect 253014 183580 253020 183592
rect 252888 183552 253020 183580
rect 252888 183540 252894 183552
rect 253014 183540 253020 183552
rect 253072 183540 253078 183592
rect 271966 183580 271972 183592
rect 271927 183552 271972 183580
rect 271966 183540 271972 183552
rect 272024 183540 272030 183592
rect 287238 183540 287244 183592
rect 287296 183580 287302 183592
rect 287422 183580 287428 183592
rect 287296 183552 287428 183580
rect 287296 183540 287302 183552
rect 287422 183540 287428 183552
rect 287480 183540 287486 183592
rect 298278 183580 298284 183592
rect 298239 183552 298284 183580
rect 298278 183540 298284 183552
rect 298336 183540 298342 183592
rect 309321 183583 309379 183589
rect 309321 183549 309333 183583
rect 309367 183580 309379 183583
rect 309502 183580 309508 183592
rect 309367 183552 309508 183580
rect 309367 183549 309379 183552
rect 309321 183543 309379 183549
rect 309502 183540 309508 183552
rect 309560 183540 309566 183592
rect 321646 183580 321652 183592
rect 321607 183552 321652 183580
rect 321646 183540 321652 183552
rect 321704 183540 321710 183592
rect 324406 183580 324412 183592
rect 324367 183552 324412 183580
rect 324406 183540 324412 183552
rect 324464 183540 324470 183592
rect 329926 183540 329932 183592
rect 329984 183580 329990 183592
rect 330110 183580 330116 183592
rect 329984 183552 330116 183580
rect 329984 183540 329990 183552
rect 330110 183540 330116 183552
rect 330168 183540 330174 183592
rect 331398 183540 331404 183592
rect 331456 183580 331462 183592
rect 331490 183580 331496 183592
rect 331456 183552 331496 183580
rect 331456 183540 331462 183552
rect 331490 183540 331496 183552
rect 331548 183540 331554 183592
rect 334342 183540 334348 183592
rect 334400 183580 334406 183592
rect 334434 183580 334440 183592
rect 334400 183552 334440 183580
rect 334400 183540 334406 183552
rect 334434 183540 334440 183552
rect 334492 183540 334498 183592
rect 336734 183540 336740 183592
rect 336792 183580 336798 183592
rect 336826 183580 336832 183592
rect 336792 183552 336832 183580
rect 336792 183540 336798 183552
rect 336826 183540 336832 183552
rect 336884 183540 336890 183592
rect 347958 183540 347964 183592
rect 348016 183580 348022 183592
rect 348050 183580 348056 183592
rect 348016 183552 348056 183580
rect 348016 183540 348022 183552
rect 348050 183540 348056 183552
rect 348108 183540 348114 183592
rect 352006 183540 352012 183592
rect 352064 183580 352070 183592
rect 352190 183580 352196 183592
rect 352064 183552 352196 183580
rect 352064 183540 352070 183552
rect 352190 183540 352196 183552
rect 352248 183540 352254 183592
rect 353478 183540 353484 183592
rect 353536 183580 353542 183592
rect 353570 183580 353576 183592
rect 353536 183552 353576 183580
rect 353536 183540 353542 183552
rect 353570 183540 353576 183552
rect 353628 183540 353634 183592
rect 356422 183540 356428 183592
rect 356480 183580 356486 183592
rect 356514 183580 356520 183592
rect 356480 183552 356520 183580
rect 356480 183540 356486 183552
rect 356514 183540 356520 183552
rect 356572 183540 356578 183592
rect 382476 183524 382504 183608
rect 270589 183515 270647 183521
rect 270589 183481 270601 183515
rect 270635 183512 270647 183515
rect 270678 183512 270684 183524
rect 270635 183484 270684 183512
rect 270635 183481 270647 183484
rect 270589 183475 270647 183481
rect 270678 183472 270684 183484
rect 270736 183472 270742 183524
rect 295702 183512 295708 183524
rect 295663 183484 295708 183512
rect 295702 183472 295708 183484
rect 295760 183472 295766 183524
rect 382458 183472 382464 183524
rect 382516 183472 382522 183524
rect 416866 183472 416872 183524
rect 416924 183512 416930 183524
rect 416958 183512 416964 183524
rect 416924 183484 416964 183512
rect 416924 183472 416930 183484
rect 416958 183472 416964 183484
rect 417016 183472 417022 183524
rect 332778 182220 332784 182232
rect 332704 182192 332784 182220
rect 332704 182164 332732 182192
rect 332778 182180 332784 182192
rect 332836 182180 332842 182232
rect 231946 182112 231952 182164
rect 232004 182152 232010 182164
rect 232130 182152 232136 182164
rect 232004 182124 232136 182152
rect 232004 182112 232010 182124
rect 232130 182112 232136 182124
rect 232188 182112 232194 182164
rect 265158 182112 265164 182164
rect 265216 182152 265222 182164
rect 265250 182152 265256 182164
rect 265216 182124 265256 182152
rect 265216 182112 265222 182124
rect 265250 182112 265256 182124
rect 265308 182112 265314 182164
rect 267182 182152 267188 182164
rect 267143 182124 267188 182152
rect 267182 182112 267188 182124
rect 267240 182112 267246 182164
rect 287238 182112 287244 182164
rect 287296 182152 287302 182164
rect 287422 182152 287428 182164
rect 287296 182124 287428 182152
rect 287296 182112 287302 182124
rect 287422 182112 287428 182124
rect 287480 182112 287486 182164
rect 292850 182112 292856 182164
rect 292908 182152 292914 182164
rect 292942 182152 292948 182164
rect 292908 182124 292948 182152
rect 292908 182112 292914 182124
rect 292942 182112 292948 182124
rect 293000 182112 293006 182164
rect 298278 182112 298284 182164
rect 298336 182152 298342 182164
rect 298462 182152 298468 182164
rect 298336 182124 298468 182152
rect 298336 182112 298342 182124
rect 298462 182112 298468 182124
rect 298520 182112 298526 182164
rect 331490 182112 331496 182164
rect 331548 182152 331554 182164
rect 331582 182152 331588 182164
rect 331548 182124 331588 182152
rect 331548 182112 331554 182124
rect 331582 182112 331588 182124
rect 331640 182112 331646 182164
rect 332686 182112 332692 182164
rect 332744 182112 332750 182164
rect 334434 182112 334440 182164
rect 334492 182152 334498 182164
rect 334526 182152 334532 182164
rect 334492 182124 334532 182152
rect 334492 182112 334498 182124
rect 334526 182112 334532 182124
rect 334584 182112 334590 182164
rect 336826 182152 336832 182164
rect 336787 182124 336832 182152
rect 336826 182112 336832 182124
rect 336884 182112 336890 182164
rect 365714 182112 365720 182164
rect 365772 182152 365778 182164
rect 365898 182152 365904 182164
rect 365772 182124 365904 182152
rect 365772 182112 365778 182124
rect 365898 182112 365904 182124
rect 365956 182112 365962 182164
rect 372614 181160 372620 181212
rect 372672 181200 372678 181212
rect 382182 181200 382188 181212
rect 372672 181172 382188 181200
rect 372672 181160 372678 181172
rect 382182 181160 382188 181172
rect 382240 181160 382246 181212
rect 364334 181024 364340 181076
rect 364392 181024 364398 181076
rect 364352 180872 364380 181024
rect 553302 180956 553308 181008
rect 553360 180996 553366 181008
rect 554958 180996 554964 181008
rect 553360 180968 554964 180996
rect 553360 180956 553366 180968
rect 554958 180956 554964 180968
rect 555016 180956 555022 181008
rect 475930 180888 475936 180940
rect 475988 180928 475994 180940
rect 476114 180928 476120 180940
rect 475988 180900 476120 180928
rect 475988 180888 475994 180900
rect 476114 180888 476120 180900
rect 476172 180888 476178 180940
rect 364334 180820 364340 180872
rect 364392 180820 364398 180872
rect 425054 180820 425060 180872
rect 425112 180860 425118 180872
rect 434530 180860 434536 180872
rect 425112 180832 434536 180860
rect 425112 180820 425118 180832
rect 434530 180820 434536 180832
rect 434588 180820 434594 180872
rect 521654 180820 521660 180872
rect 521712 180860 521718 180872
rect 526438 180860 526444 180872
rect 521712 180832 526444 180860
rect 521712 180820 521718 180832
rect 526438 180820 526444 180832
rect 526496 180820 526502 180872
rect 255498 180792 255504 180804
rect 255459 180764 255504 180792
rect 255498 180752 255504 180764
rect 255556 180752 255562 180804
rect 347961 180795 348019 180801
rect 347961 180761 347973 180795
rect 348007 180792 348019 180795
rect 348050 180792 348056 180804
rect 348007 180764 348056 180792
rect 348007 180761 348019 180764
rect 347961 180755 348019 180761
rect 348050 180752 348056 180764
rect 348108 180752 348114 180804
rect 352006 180752 352012 180804
rect 352064 180792 352070 180804
rect 352101 180795 352159 180801
rect 352101 180792 352113 180795
rect 352064 180764 352113 180792
rect 352064 180752 352070 180764
rect 352101 180761 352113 180764
rect 352147 180761 352159 180795
rect 352101 180755 352159 180761
rect 353481 180795 353539 180801
rect 353481 180761 353493 180795
rect 353527 180792 353539 180795
rect 353570 180792 353576 180804
rect 353527 180764 353576 180792
rect 353527 180761 353539 180764
rect 353481 180755 353539 180761
rect 353570 180752 353576 180764
rect 353628 180752 353634 180804
rect 357618 179432 357624 179444
rect 357579 179404 357624 179432
rect 357618 179392 357624 179404
rect 357676 179392 357682 179444
rect 359090 179256 359096 179308
rect 359148 179296 359154 179308
rect 359182 179296 359188 179308
rect 359148 179268 359188 179296
rect 359148 179256 359154 179268
rect 359182 179256 359188 179268
rect 359240 179256 359246 179308
rect 252741 178823 252799 178829
rect 252741 178789 252753 178823
rect 252787 178820 252799 178823
rect 252830 178820 252836 178832
rect 252787 178792 252836 178820
rect 252787 178789 252799 178792
rect 252741 178783 252799 178789
rect 252830 178780 252836 178792
rect 252888 178780 252894 178832
rect 480346 178780 480352 178832
rect 480404 178780 480410 178832
rect 480364 178696 480392 178780
rect 480346 178644 480352 178696
rect 480404 178644 480410 178696
rect 236273 178075 236331 178081
rect 236273 178041 236285 178075
rect 236319 178072 236331 178075
rect 236454 178072 236460 178084
rect 236319 178044 236460 178072
rect 236319 178041 236331 178044
rect 236273 178035 236331 178041
rect 236454 178032 236460 178044
rect 236512 178032 236518 178084
rect 364610 176740 364616 176792
rect 364668 176740 364674 176792
rect 386690 176740 386696 176792
rect 386748 176740 386754 176792
rect 329926 176672 329932 176724
rect 329984 176672 329990 176724
rect 244458 176604 244464 176656
rect 244516 176604 244522 176656
rect 244476 176520 244504 176604
rect 329944 176576 329972 176672
rect 364628 176656 364656 176740
rect 386708 176656 386736 176740
rect 346578 176604 346584 176656
rect 346636 176604 346642 176656
rect 364610 176604 364616 176656
rect 364668 176604 364674 176656
rect 386690 176604 386696 176656
rect 386748 176604 386754 176656
rect 397730 176644 397736 176656
rect 397691 176616 397736 176644
rect 397730 176604 397736 176616
rect 397788 176604 397794 176656
rect 330018 176576 330024 176588
rect 329944 176548 330024 176576
rect 330018 176536 330024 176548
rect 330076 176536 330082 176588
rect 336826 176576 336832 176588
rect 336787 176548 336832 176576
rect 336826 176536 336832 176548
rect 336884 176536 336890 176588
rect 346596 176520 346624 176604
rect 244458 176468 244464 176520
rect 244516 176468 244522 176520
rect 249978 176468 249984 176520
rect 250036 176468 250042 176520
rect 346578 176468 346584 176520
rect 346636 176468 346642 176520
rect 249996 176384 250024 176468
rect 249978 176332 249984 176384
rect 250036 176332 250042 176384
rect 309502 174020 309508 174072
rect 309560 174020 309566 174072
rect 294230 173992 294236 174004
rect 294156 173964 294236 173992
rect 241790 173884 241796 173936
rect 241848 173924 241854 173936
rect 241974 173924 241980 173936
rect 241848 173896 241980 173924
rect 241848 173884 241854 173896
rect 241974 173884 241980 173896
rect 242032 173884 242038 173936
rect 243170 173884 243176 173936
rect 243228 173924 243234 173936
rect 243262 173924 243268 173936
rect 243228 173896 243268 173924
rect 243228 173884 243234 173896
rect 243262 173884 243268 173896
rect 243320 173884 243326 173936
rect 252738 173924 252744 173936
rect 252699 173896 252744 173924
rect 252738 173884 252744 173896
rect 252796 173884 252802 173936
rect 254118 173884 254124 173936
rect 254176 173924 254182 173936
rect 254302 173924 254308 173936
rect 254176 173896 254308 173924
rect 254176 173884 254182 173896
rect 254302 173884 254308 173896
rect 254360 173884 254366 173936
rect 259730 173884 259736 173936
rect 259788 173924 259794 173936
rect 259822 173924 259828 173936
rect 259788 173896 259828 173924
rect 259788 173884 259794 173896
rect 259822 173884 259828 173896
rect 259880 173884 259886 173936
rect 266446 173884 266452 173936
rect 266504 173924 266510 173936
rect 266538 173924 266544 173936
rect 266504 173896 266544 173924
rect 266504 173884 266510 173896
rect 266538 173884 266544 173896
rect 266596 173884 266602 173936
rect 270678 173884 270684 173936
rect 270736 173924 270742 173936
rect 270862 173924 270868 173936
rect 270736 173896 270868 173924
rect 270736 173884 270742 173896
rect 270862 173884 270868 173896
rect 270920 173884 270926 173936
rect 271966 173884 271972 173936
rect 272024 173924 272030 173936
rect 272058 173924 272064 173936
rect 272024 173896 272064 173924
rect 272024 173884 272030 173896
rect 272058 173884 272064 173896
rect 272116 173884 272122 173936
rect 288434 173884 288440 173936
rect 288492 173924 288498 173936
rect 288618 173924 288624 173936
rect 288492 173896 288624 173924
rect 288492 173884 288498 173896
rect 288618 173884 288624 173896
rect 288676 173884 288682 173936
rect 294156 173868 294184 173964
rect 294230 173952 294236 173964
rect 294288 173952 294294 174004
rect 308122 173884 308128 173936
rect 308180 173924 308186 173936
rect 308214 173924 308220 173936
rect 308180 173896 308220 173924
rect 308180 173884 308186 173896
rect 308214 173884 308220 173896
rect 308272 173884 308278 173936
rect 309520 173868 309548 174020
rect 310698 173884 310704 173936
rect 310756 173924 310762 173936
rect 310882 173924 310888 173936
rect 310756 173896 310888 173924
rect 310756 173884 310762 173896
rect 310882 173884 310888 173896
rect 310940 173884 310946 173936
rect 321646 173884 321652 173936
rect 321704 173924 321710 173936
rect 321738 173924 321744 173936
rect 321704 173896 321744 173924
rect 321704 173884 321710 173896
rect 321738 173884 321744 173896
rect 321796 173884 321802 173936
rect 324406 173884 324412 173936
rect 324464 173924 324470 173936
rect 324498 173924 324504 173936
rect 324464 173896 324504 173924
rect 324464 173884 324470 173896
rect 324498 173884 324504 173896
rect 324556 173884 324562 173936
rect 327166 173884 327172 173936
rect 327224 173924 327230 173936
rect 327258 173924 327264 173936
rect 327224 173896 327264 173924
rect 327224 173884 327230 173896
rect 327258 173884 327264 173896
rect 327316 173884 327322 173936
rect 370038 173884 370044 173936
rect 370096 173924 370102 173936
rect 370130 173924 370136 173936
rect 370096 173896 370136 173924
rect 370096 173884 370102 173896
rect 370130 173884 370136 173896
rect 370188 173884 370194 173936
rect 397730 173924 397736 173936
rect 397691 173896 397736 173924
rect 397730 173884 397736 173896
rect 397788 173884 397794 173936
rect 408770 173884 408776 173936
rect 408828 173924 408834 173936
rect 408954 173924 408960 173936
rect 408828 173896 408960 173924
rect 408828 173884 408834 173896
rect 408954 173884 408960 173896
rect 409012 173884 409018 173936
rect 422478 173884 422484 173936
rect 422536 173924 422542 173936
rect 422662 173924 422668 173936
rect 422536 173896 422668 173924
rect 422536 173884 422542 173896
rect 422662 173884 422668 173896
rect 422720 173884 422726 173936
rect 433610 173884 433616 173936
rect 433668 173924 433674 173936
rect 433702 173924 433708 173936
rect 433668 173896 433708 173924
rect 433668 173884 433674 173896
rect 433702 173884 433708 173896
rect 433760 173884 433766 173936
rect 472158 173884 472164 173936
rect 472216 173924 472222 173936
rect 472342 173924 472348 173936
rect 472216 173896 472348 173924
rect 472216 173884 472222 173896
rect 472342 173884 472348 173896
rect 472400 173884 472406 173936
rect 294138 173816 294144 173868
rect 294196 173816 294202 173868
rect 309502 173816 309508 173868
rect 309560 173816 309566 173868
rect 267182 173312 267188 173324
rect 267143 173284 267188 173312
rect 267182 173272 267188 173284
rect 267240 173272 267246 173324
rect 295610 172524 295616 172576
rect 295668 172564 295674 172576
rect 295702 172564 295708 172576
rect 295668 172536 295708 172564
rect 295668 172524 295674 172536
rect 295702 172524 295708 172536
rect 295760 172524 295766 172576
rect 254118 172496 254124 172508
rect 254079 172468 254124 172496
rect 254118 172456 254124 172468
rect 254176 172456 254182 172508
rect 259641 172499 259699 172505
rect 259641 172465 259653 172499
rect 259687 172496 259699 172499
rect 259730 172496 259736 172508
rect 259687 172468 259736 172496
rect 259687 172465 259699 172468
rect 259641 172459 259699 172465
rect 259730 172456 259736 172468
rect 259788 172456 259794 172508
rect 271969 172499 272027 172505
rect 271969 172465 271981 172499
rect 272015 172496 272027 172499
rect 272058 172496 272064 172508
rect 272015 172468 272064 172496
rect 272015 172465 272027 172468
rect 271969 172459 272027 172465
rect 272058 172456 272064 172468
rect 272116 172456 272122 172508
rect 292758 172496 292764 172508
rect 292719 172468 292764 172496
rect 292758 172456 292764 172468
rect 292816 172456 292822 172508
rect 332686 172456 332692 172508
rect 332744 172496 332750 172508
rect 332778 172496 332784 172508
rect 332744 172468 332784 172496
rect 332744 172456 332750 172468
rect 332778 172456 332784 172468
rect 332836 172456 332842 172508
rect 342349 172499 342407 172505
rect 342349 172465 342361 172499
rect 342395 172496 342407 172499
rect 342530 172496 342536 172508
rect 342395 172468 342536 172496
rect 342395 172465 342407 172468
rect 342349 172459 342407 172465
rect 342530 172456 342536 172468
rect 342588 172456 342594 172508
rect 451734 172456 451740 172508
rect 451792 172496 451798 172508
rect 452010 172496 452016 172508
rect 451792 172468 452016 172496
rect 451792 172456 451798 172468
rect 452010 172456 452016 172468
rect 452068 172456 452074 172508
rect 288342 170076 288348 170128
rect 288400 170116 288406 170128
rect 296622 170116 296628 170128
rect 288400 170088 296628 170116
rect 288400 170076 288406 170088
rect 296622 170076 296628 170088
rect 296680 170076 296686 170128
rect 328362 170008 328368 170060
rect 328420 170048 328426 170060
rect 336642 170048 336648 170060
rect 328420 170020 336648 170048
rect 328420 170008 328426 170020
rect 336642 170008 336648 170020
rect 336700 170008 336706 170060
rect 365714 169940 365720 169992
rect 365772 169980 365778 169992
rect 368290 169980 368296 169992
rect 365772 169952 368296 169980
rect 365772 169940 365778 169952
rect 368290 169940 368296 169952
rect 368348 169940 368354 169992
rect 454034 169940 454040 169992
rect 454092 169980 454098 169992
rect 458174 169980 458180 169992
rect 454092 169952 458180 169980
rect 454092 169940 454098 169952
rect 458174 169940 458180 169952
rect 458232 169940 458238 169992
rect 514570 169940 514576 169992
rect 514628 169980 514634 169992
rect 516870 169980 516876 169992
rect 514628 169952 516876 169980
rect 514628 169940 514634 169952
rect 516870 169940 516876 169952
rect 516928 169940 516934 169992
rect 475930 169872 475936 169924
rect 475988 169912 475994 169924
rect 476114 169912 476120 169924
rect 475988 169884 476120 169912
rect 475988 169872 475994 169884
rect 476114 169872 476120 169884
rect 476172 169872 476178 169924
rect 309042 169804 309048 169856
rect 309100 169844 309106 169856
rect 317322 169844 317328 169856
rect 309100 169816 317328 169844
rect 309100 169804 309106 169816
rect 317322 169804 317328 169816
rect 317380 169804 317386 169856
rect 425054 169804 425060 169856
rect 425112 169844 425118 169856
rect 434530 169844 434536 169856
rect 425112 169816 434536 169844
rect 425112 169804 425118 169816
rect 434530 169804 434536 169816
rect 434588 169804 434594 169856
rect 524230 169804 524236 169856
rect 524288 169844 524294 169856
rect 526438 169844 526444 169856
rect 524288 169816 526444 169844
rect 524288 169804 524294 169816
rect 526438 169804 526444 169816
rect 526496 169804 526502 169856
rect 299382 169668 299388 169720
rect 299440 169708 299446 169720
rect 302970 169708 302976 169720
rect 299440 169680 302976 169708
rect 299440 169668 299446 169680
rect 302970 169668 302976 169680
rect 303028 169668 303034 169720
rect 376938 169056 376944 169108
rect 376996 169096 377002 169108
rect 377122 169096 377128 169108
rect 376996 169068 377128 169096
rect 376996 169056 377002 169068
rect 377122 169056 377128 169068
rect 377180 169056 377186 169108
rect 480346 169056 480352 169108
rect 480404 169096 480410 169108
rect 480530 169096 480536 169108
rect 480404 169068 480536 169096
rect 480404 169056 480410 169068
rect 480530 169056 480536 169068
rect 480588 169056 480594 169108
rect 321462 168580 321468 168632
rect 321520 168620 321526 168632
rect 321738 168620 321744 168632
rect 321520 168592 321744 168620
rect 321520 168580 321526 168592
rect 321738 168580 321744 168592
rect 321796 168580 321802 168632
rect 382274 167628 382280 167680
rect 382332 167668 382338 167680
rect 382461 167671 382519 167677
rect 382461 167668 382473 167671
rect 382332 167640 382473 167668
rect 382332 167628 382338 167640
rect 382461 167637 382473 167640
rect 382507 167637 382519 167671
rect 382461 167631 382519 167637
rect 242989 167127 243047 167133
rect 242989 167093 243001 167127
rect 243035 167124 243047 167127
rect 243170 167124 243176 167136
rect 243035 167096 243176 167124
rect 243035 167093 243047 167096
rect 242989 167087 243047 167093
rect 243170 167084 243176 167096
rect 243228 167084 243234 167136
rect 356514 167124 356520 167136
rect 356440 167096 356520 167124
rect 233326 167016 233332 167068
rect 233384 167056 233390 167068
rect 233510 167056 233516 167068
rect 233384 167028 233516 167056
rect 233384 167016 233390 167028
rect 233510 167016 233516 167028
rect 233568 167016 233574 167068
rect 270678 167016 270684 167068
rect 270736 167016 270742 167068
rect 318886 167016 318892 167068
rect 318944 167056 318950 167068
rect 319070 167056 319076 167068
rect 318944 167028 319076 167056
rect 318944 167016 318950 167028
rect 319070 167016 319076 167028
rect 319128 167016 319134 167068
rect 254118 166988 254124 167000
rect 254079 166960 254124 166988
rect 254118 166948 254124 166960
rect 254176 166948 254182 167000
rect 255498 166988 255504 167000
rect 255459 166960 255504 166988
rect 255498 166948 255504 166960
rect 255556 166948 255562 167000
rect 270696 166920 270724 167016
rect 356440 166932 356468 167096
rect 356514 167084 356520 167096
rect 356572 167084 356578 167136
rect 400398 167016 400404 167068
rect 400456 167056 400462 167068
rect 400582 167056 400588 167068
rect 400456 167028 400588 167056
rect 400456 167016 400462 167028
rect 400582 167016 400588 167028
rect 400640 167016 400646 167068
rect 422294 167016 422300 167068
rect 422352 167056 422358 167068
rect 422478 167056 422484 167068
rect 422352 167028 422484 167056
rect 422352 167016 422358 167028
rect 422478 167016 422484 167028
rect 422536 167016 422542 167068
rect 466454 167016 466460 167068
rect 466512 167056 466518 167068
rect 466638 167056 466644 167068
rect 466512 167028 466644 167056
rect 466512 167016 466518 167028
rect 466638 167016 466644 167028
rect 466696 167016 466702 167068
rect 270770 166920 270776 166932
rect 270696 166892 270776 166920
rect 270770 166880 270776 166892
rect 270828 166880 270834 166932
rect 356422 166880 356428 166932
rect 356480 166880 356486 166932
rect 2774 165112 2780 165164
rect 2832 165152 2838 165164
rect 4798 165152 4804 165164
rect 2832 165124 4804 165152
rect 2832 165112 2838 165124
rect 4798 165112 4804 165124
rect 4856 165112 4862 165164
rect 231946 164228 231952 164280
rect 232004 164268 232010 164280
rect 232038 164268 232044 164280
rect 232004 164240 232044 164268
rect 232004 164228 232010 164240
rect 232038 164228 232044 164240
rect 232096 164228 232102 164280
rect 298186 164228 298192 164280
rect 298244 164268 298250 164280
rect 298278 164268 298284 164280
rect 298244 164240 298284 164268
rect 298244 164228 298250 164240
rect 298278 164228 298284 164240
rect 298336 164228 298342 164280
rect 393222 164228 393228 164280
rect 393280 164228 393286 164280
rect 265161 164203 265219 164209
rect 265161 164169 265173 164203
rect 265207 164200 265219 164203
rect 265250 164200 265256 164212
rect 265207 164172 265256 164200
rect 265207 164169 265219 164172
rect 265161 164163 265219 164169
rect 265250 164160 265256 164172
rect 265308 164160 265314 164212
rect 266906 164160 266912 164212
rect 266964 164200 266970 164212
rect 266998 164200 267004 164212
rect 266964 164172 267004 164200
rect 266964 164160 266970 164172
rect 266998 164160 267004 164172
rect 267056 164160 267062 164212
rect 292758 164200 292764 164212
rect 292719 164172 292764 164200
rect 292758 164160 292764 164172
rect 292816 164160 292822 164212
rect 308030 164160 308036 164212
rect 308088 164200 308094 164212
rect 308214 164200 308220 164212
rect 308088 164172 308220 164200
rect 308088 164160 308094 164172
rect 308214 164160 308220 164172
rect 308272 164160 308278 164212
rect 310698 164160 310704 164212
rect 310756 164200 310762 164212
rect 310882 164200 310888 164212
rect 310756 164172 310888 164200
rect 310756 164160 310762 164172
rect 310882 164160 310888 164172
rect 310940 164160 310946 164212
rect 327166 164160 327172 164212
rect 327224 164160 327230 164212
rect 329926 164160 329932 164212
rect 329984 164200 329990 164212
rect 330110 164200 330116 164212
rect 329984 164172 330116 164200
rect 329984 164160 329990 164172
rect 330110 164160 330116 164172
rect 330168 164160 330174 164212
rect 370041 164203 370099 164209
rect 370041 164169 370053 164203
rect 370087 164200 370099 164203
rect 370130 164200 370136 164212
rect 370087 164172 370136 164200
rect 370087 164169 370099 164172
rect 370041 164163 370099 164169
rect 370130 164160 370136 164172
rect 370188 164160 370194 164212
rect 376938 164200 376944 164212
rect 376899 164172 376944 164200
rect 376938 164160 376944 164172
rect 376996 164160 377002 164212
rect 386690 164160 386696 164212
rect 386748 164200 386754 164212
rect 386782 164200 386788 164212
rect 386748 164172 386788 164200
rect 386748 164160 386754 164172
rect 386782 164160 386788 164172
rect 386840 164160 386846 164212
rect 327184 164132 327212 164160
rect 393240 164144 393268 164228
rect 397730 164200 397736 164212
rect 397691 164172 397736 164200
rect 397730 164160 397736 164172
rect 397788 164160 397794 164212
rect 400490 164200 400496 164212
rect 400451 164172 400496 164200
rect 400490 164160 400496 164172
rect 400548 164160 400554 164212
rect 408402 164160 408408 164212
rect 408460 164200 408466 164212
rect 408586 164200 408592 164212
rect 408460 164172 408592 164200
rect 408460 164160 408466 164172
rect 408586 164160 408592 164172
rect 408644 164160 408650 164212
rect 416866 164160 416872 164212
rect 416924 164200 416930 164212
rect 416958 164200 416964 164212
rect 416924 164172 416964 164200
rect 416924 164160 416930 164172
rect 416958 164160 416964 164172
rect 417016 164160 417022 164212
rect 422386 164200 422392 164212
rect 422347 164172 422392 164200
rect 422386 164160 422392 164172
rect 422444 164160 422450 164212
rect 466546 164200 466552 164212
rect 466507 164172 466552 164200
rect 466546 164160 466552 164172
rect 466604 164160 466610 164212
rect 472066 164160 472072 164212
rect 472124 164200 472130 164212
rect 472342 164200 472348 164212
rect 472124 164172 472348 164200
rect 472124 164160 472130 164172
rect 472342 164160 472348 164172
rect 472400 164160 472406 164212
rect 480257 164203 480315 164209
rect 480257 164169 480269 164203
rect 480303 164200 480315 164203
rect 480346 164200 480352 164212
rect 480303 164172 480352 164200
rect 480303 164169 480315 164172
rect 480257 164163 480315 164169
rect 480346 164160 480352 164172
rect 480404 164160 480410 164212
rect 327258 164132 327264 164144
rect 327184 164104 327264 164132
rect 327258 164092 327264 164104
rect 327316 164092 327322 164144
rect 393222 164092 393228 164144
rect 393280 164092 393286 164144
rect 242986 162908 242992 162920
rect 242947 162880 242992 162908
rect 242986 162868 242992 162880
rect 243044 162868 243050 162920
rect 259638 162908 259644 162920
rect 259599 162880 259644 162908
rect 259638 162868 259644 162880
rect 259696 162868 259702 162920
rect 271966 162908 271972 162920
rect 271927 162880 271972 162908
rect 271966 162868 271972 162880
rect 272024 162868 272030 162920
rect 342346 162908 342352 162920
rect 342307 162880 342352 162908
rect 342346 162868 342352 162880
rect 342404 162868 342410 162920
rect 347958 162908 347964 162920
rect 347919 162880 347964 162908
rect 347958 162868 347964 162880
rect 348016 162868 348022 162920
rect 352098 162908 352104 162920
rect 352059 162880 352104 162908
rect 352098 162868 352104 162880
rect 352156 162868 352162 162920
rect 353478 162908 353484 162920
rect 353439 162880 353484 162908
rect 353478 162868 353484 162880
rect 353536 162868 353542 162920
rect 298278 162840 298284 162852
rect 298239 162812 298284 162840
rect 298278 162800 298284 162812
rect 298336 162800 298342 162852
rect 308214 162800 308220 162852
rect 308272 162840 308278 162852
rect 308398 162840 308404 162852
rect 308272 162812 308404 162840
rect 308272 162800 308278 162812
rect 308398 162800 308404 162812
rect 308456 162800 308462 162852
rect 327258 162800 327264 162852
rect 327316 162840 327322 162852
rect 327442 162840 327448 162852
rect 327316 162812 327448 162840
rect 327316 162800 327322 162812
rect 327442 162800 327448 162812
rect 327500 162800 327506 162852
rect 393222 162840 393228 162852
rect 393183 162812 393228 162840
rect 393222 162800 393228 162812
rect 393280 162800 393286 162852
rect 451553 162843 451611 162849
rect 451553 162809 451565 162843
rect 451599 162840 451611 162843
rect 451734 162840 451740 162852
rect 451599 162812 451740 162840
rect 451599 162809 451611 162812
rect 451553 162803 451611 162809
rect 451734 162800 451740 162812
rect 451792 162800 451798 162852
rect 334526 161412 334532 161424
rect 334487 161384 334532 161412
rect 334526 161372 334532 161384
rect 334584 161372 334590 161424
rect 356422 161344 356428 161356
rect 356383 161316 356428 161344
rect 356422 161304 356428 161316
rect 356480 161304 356486 161356
rect 321462 159332 321468 159384
rect 321520 159372 321526 159384
rect 321738 159372 321744 159384
rect 321520 159344 321744 159372
rect 321520 159332 321526 159344
rect 321738 159332 321744 159344
rect 321796 159332 321802 159384
rect 252554 157972 252560 158024
rect 252612 158012 252618 158024
rect 252738 158012 252744 158024
rect 252612 157984 252744 158012
rect 252612 157972 252618 157984
rect 252738 157972 252744 157984
rect 252796 157972 252802 158024
rect 271966 158012 271972 158024
rect 271927 157984 271972 158012
rect 271966 157972 271972 157984
rect 272024 157972 272030 158024
rect 405734 157700 405740 157752
rect 405792 157740 405798 157752
rect 415302 157740 415308 157752
rect 405792 157712 415308 157740
rect 405792 157700 405798 157712
rect 415302 157700 415308 157712
rect 415360 157700 415366 157752
rect 387978 157428 387984 157480
rect 388036 157428 388042 157480
rect 521654 157428 521660 157480
rect 521712 157468 521718 157480
rect 526438 157468 526444 157480
rect 521712 157440 526444 157468
rect 521712 157428 521718 157440
rect 526438 157428 526444 157440
rect 526496 157428 526502 157480
rect 232038 157360 232044 157412
rect 232096 157360 232102 157412
rect 324498 157400 324504 157412
rect 324424 157372 324504 157400
rect 232056 157332 232084 157360
rect 232130 157332 232136 157344
rect 232056 157304 232136 157332
rect 232130 157292 232136 157304
rect 232188 157292 232194 157344
rect 298278 157332 298284 157344
rect 298239 157304 298284 157332
rect 298278 157292 298284 157304
rect 298336 157292 298342 157344
rect 324424 157276 324452 157372
rect 324498 157360 324504 157372
rect 324556 157360 324562 157412
rect 387996 157344 388024 157428
rect 346578 157292 346584 157344
rect 346636 157292 346642 157344
rect 387978 157292 387984 157344
rect 388036 157292 388042 157344
rect 400490 157332 400496 157344
rect 400451 157304 400496 157332
rect 400490 157292 400496 157304
rect 400548 157292 400554 157344
rect 422386 157332 422392 157344
rect 422347 157304 422392 157332
rect 422386 157292 422392 157304
rect 422444 157292 422450 157344
rect 466546 157332 466552 157344
rect 466507 157304 466552 157332
rect 466546 157292 466552 157304
rect 466604 157292 466610 157344
rect 324406 157224 324412 157276
rect 324464 157224 324470 157276
rect 346596 157208 346624 157292
rect 346578 157156 346584 157208
rect 346636 157156 346642 157208
rect 292761 155907 292819 155913
rect 292761 155873 292773 155907
rect 292807 155904 292819 155907
rect 292850 155904 292856 155916
rect 292807 155876 292856 155904
rect 292807 155873 292819 155876
rect 292761 155867 292819 155873
rect 292850 155864 292856 155876
rect 292908 155864 292914 155916
rect 265158 154680 265164 154692
rect 265119 154652 265164 154680
rect 265158 154640 265164 154652
rect 265216 154640 265222 154692
rect 266538 154572 266544 154624
rect 266596 154612 266602 154624
rect 266630 154612 266636 154624
rect 266596 154584 266636 154612
rect 266596 154572 266602 154584
rect 266630 154572 266636 154584
rect 266688 154572 266694 154624
rect 370038 154612 370044 154624
rect 369999 154584 370044 154612
rect 370038 154572 370044 154584
rect 370096 154572 370102 154624
rect 376938 154612 376944 154624
rect 376899 154584 376944 154612
rect 376938 154572 376944 154584
rect 376996 154572 377002 154624
rect 382458 154612 382464 154624
rect 382419 154584 382464 154612
rect 382458 154572 382464 154584
rect 382516 154572 382522 154624
rect 397730 154612 397736 154624
rect 397691 154584 397736 154612
rect 397730 154572 397736 154584
rect 397788 154572 397794 154624
rect 242986 154544 242992 154556
rect 242947 154516 242992 154544
rect 242986 154504 242992 154516
rect 243044 154504 243050 154556
rect 331398 154544 331404 154556
rect 331359 154516 331404 154544
rect 331398 154504 331404 154516
rect 331456 154504 331462 154556
rect 375558 154544 375564 154556
rect 375519 154516 375564 154544
rect 375558 154504 375564 154516
rect 375616 154504 375622 154556
rect 381078 154544 381084 154556
rect 381039 154516 381084 154544
rect 381078 154504 381084 154516
rect 381136 154504 381142 154556
rect 386598 154504 386604 154556
rect 386656 154544 386662 154556
rect 386782 154544 386788 154556
rect 386656 154516 386788 154544
rect 386656 154504 386662 154516
rect 386782 154504 386788 154516
rect 386840 154504 386846 154556
rect 392118 154544 392124 154556
rect 392079 154516 392124 154544
rect 392118 154504 392124 154516
rect 392176 154504 392182 154556
rect 254118 153212 254124 153264
rect 254176 153252 254182 153264
rect 254394 153252 254400 153264
rect 254176 153224 254400 153252
rect 254176 153212 254182 153224
rect 254394 153212 254400 153224
rect 254452 153212 254458 153264
rect 480254 153252 480260 153264
rect 480215 153224 480260 153252
rect 480254 153212 480260 153224
rect 480312 153212 480318 153264
rect 240226 153144 240232 153196
rect 240284 153184 240290 153196
rect 240502 153184 240508 153196
rect 240284 153156 240508 153184
rect 240284 153144 240290 153156
rect 240502 153144 240508 153156
rect 240560 153144 240566 153196
rect 281718 153144 281724 153196
rect 281776 153184 281782 153196
rect 281810 153184 281816 153196
rect 281776 153156 281816 153184
rect 281776 153144 281782 153156
rect 281810 153144 281816 153156
rect 281868 153144 281874 153196
rect 334529 153187 334587 153193
rect 334529 153153 334541 153187
rect 334575 153184 334587 153187
rect 334618 153184 334624 153196
rect 334575 153156 334624 153184
rect 334575 153153 334587 153156
rect 334529 153147 334587 153153
rect 334618 153144 334624 153156
rect 334676 153144 334682 153196
rect 254394 153116 254400 153128
rect 254355 153088 254400 153116
rect 254394 153076 254400 153088
rect 254452 153076 254458 153128
rect 356422 151824 356428 151836
rect 356383 151796 356428 151824
rect 356422 151784 356428 151796
rect 356480 151784 356486 151836
rect 236362 151756 236368 151768
rect 236323 151728 236368 151756
rect 236362 151716 236368 151728
rect 236420 151716 236426 151768
rect 334437 151759 334495 151765
rect 334437 151725 334449 151759
rect 334483 151756 334495 151759
rect 334618 151756 334624 151768
rect 334483 151728 334624 151756
rect 334483 151725 334495 151728
rect 334437 151719 334495 151725
rect 334618 151716 334624 151728
rect 334676 151716 334682 151768
rect 271966 148628 271972 148640
rect 271927 148600 271972 148628
rect 271966 148588 271972 148600
rect 272024 148588 272030 148640
rect 265158 147704 265164 147756
rect 265216 147704 265222 147756
rect 433610 147704 433616 147756
rect 433668 147704 433674 147756
rect 233326 147636 233332 147688
rect 233384 147676 233390 147688
rect 233510 147676 233516 147688
rect 233384 147648 233516 147676
rect 233384 147636 233390 147648
rect 233510 147636 233516 147648
rect 233568 147636 233574 147688
rect 265176 147620 265204 147704
rect 309318 147636 309324 147688
rect 309376 147636 309382 147688
rect 318886 147636 318892 147688
rect 318944 147676 318950 147688
rect 319070 147676 319076 147688
rect 318944 147648 319076 147676
rect 318944 147636 318950 147648
rect 319070 147636 319076 147648
rect 319128 147636 319134 147688
rect 364518 147636 364524 147688
rect 364576 147636 364582 147688
rect 370038 147636 370044 147688
rect 370096 147636 370102 147688
rect 400398 147636 400404 147688
rect 400456 147676 400462 147688
rect 400582 147676 400588 147688
rect 400456 147648 400588 147676
rect 400456 147636 400462 147648
rect 400582 147636 400588 147648
rect 400640 147636 400646 147688
rect 422294 147636 422300 147688
rect 422352 147676 422358 147688
rect 422478 147676 422484 147688
rect 422352 147648 422484 147676
rect 422352 147636 422358 147648
rect 422478 147636 422484 147648
rect 422536 147636 422542 147688
rect 242989 147611 243047 147617
rect 242989 147577 243001 147611
rect 243035 147608 243047 147611
rect 243078 147608 243084 147620
rect 243035 147580 243084 147608
rect 243035 147577 243047 147580
rect 242989 147571 243047 147577
rect 243078 147568 243084 147580
rect 243136 147568 243142 147620
rect 265158 147568 265164 147620
rect 265216 147568 265222 147620
rect 292758 147608 292764 147620
rect 292719 147580 292764 147608
rect 292758 147568 292764 147580
rect 292816 147568 292822 147620
rect 309336 147608 309364 147636
rect 309410 147608 309416 147620
rect 309336 147580 309416 147608
rect 309410 147568 309416 147580
rect 309468 147568 309474 147620
rect 364536 147608 364564 147636
rect 364610 147608 364616 147620
rect 364536 147580 364616 147608
rect 364610 147568 364616 147580
rect 364668 147568 364674 147620
rect 370056 147608 370084 147636
rect 433628 147620 433656 147704
rect 466454 147636 466460 147688
rect 466512 147676 466518 147688
rect 466638 147676 466644 147688
rect 466512 147648 466644 147676
rect 466512 147636 466518 147648
rect 466638 147636 466644 147648
rect 466696 147636 466702 147688
rect 370130 147608 370136 147620
rect 370056 147580 370136 147608
rect 370130 147568 370136 147580
rect 370188 147568 370194 147620
rect 375558 147608 375564 147620
rect 375519 147580 375564 147608
rect 375558 147568 375564 147580
rect 375616 147568 375622 147620
rect 381078 147608 381084 147620
rect 381039 147580 381084 147608
rect 381078 147568 381084 147580
rect 381136 147568 381142 147620
rect 392118 147608 392124 147620
rect 392079 147580 392124 147608
rect 392118 147568 392124 147580
rect 392176 147568 392182 147620
rect 433610 147568 433616 147620
rect 433668 147568 433674 147620
rect 451550 147608 451556 147620
rect 451511 147580 451556 147608
rect 451550 147568 451556 147580
rect 451608 147568 451614 147620
rect 331401 147475 331459 147481
rect 331401 147441 331413 147475
rect 331447 147472 331459 147475
rect 331490 147472 331496 147484
rect 331447 147444 331496 147472
rect 331447 147441 331459 147444
rect 331401 147435 331459 147441
rect 331490 147432 331496 147444
rect 331548 147432 331554 147484
rect 393222 145024 393228 145036
rect 393183 144996 393228 145024
rect 393222 144984 393228 144996
rect 393280 144984 393286 145036
rect 252738 144916 252744 144968
rect 252796 144956 252802 144968
rect 252830 144956 252836 144968
rect 252796 144928 252836 144956
rect 252796 144916 252802 144928
rect 252830 144916 252836 144928
rect 252888 144916 252894 144968
rect 283098 144956 283104 144968
rect 283024 144928 283104 144956
rect 283024 144900 283052 144928
rect 283098 144916 283104 144928
rect 283156 144916 283162 144968
rect 308122 144916 308128 144968
rect 308180 144956 308186 144968
rect 308214 144956 308220 144968
rect 308180 144928 308220 144956
rect 308180 144916 308186 144928
rect 308214 144916 308220 144928
rect 308272 144916 308278 144968
rect 397730 144956 397736 144968
rect 397691 144928 397736 144956
rect 397730 144916 397736 144928
rect 397788 144916 397794 144968
rect 243170 144848 243176 144900
rect 243228 144888 243234 144900
rect 243262 144888 243268 144900
rect 243228 144860 243268 144888
rect 243228 144848 243234 144860
rect 243262 144848 243268 144860
rect 243320 144848 243326 144900
rect 271966 144848 271972 144900
rect 272024 144888 272030 144900
rect 272058 144888 272064 144900
rect 272024 144860 272064 144888
rect 272024 144848 272030 144860
rect 272058 144848 272064 144860
rect 272116 144848 272122 144900
rect 283006 144848 283012 144900
rect 283064 144848 283070 144900
rect 292758 144888 292764 144900
rect 292719 144860 292764 144888
rect 292758 144848 292764 144860
rect 292816 144848 292822 144900
rect 294046 144848 294052 144900
rect 294104 144888 294110 144900
rect 294230 144888 294236 144900
rect 294104 144860 294236 144888
rect 294104 144848 294110 144860
rect 294230 144848 294236 144860
rect 294288 144848 294294 144900
rect 295610 144848 295616 144900
rect 295668 144888 295674 144900
rect 295702 144888 295708 144900
rect 295668 144860 295708 144888
rect 295668 144848 295674 144860
rect 295702 144848 295708 144860
rect 295760 144848 295766 144900
rect 298278 144848 298284 144900
rect 298336 144888 298342 144900
rect 298462 144888 298468 144900
rect 298336 144860 298468 144888
rect 298336 144848 298342 144860
rect 298462 144848 298468 144860
rect 298520 144848 298526 144900
rect 347958 144848 347964 144900
rect 348016 144888 348022 144900
rect 348050 144888 348056 144900
rect 348016 144860 348056 144888
rect 348016 144848 348022 144860
rect 348050 144848 348056 144860
rect 348108 144848 348114 144900
rect 352006 144848 352012 144900
rect 352064 144888 352070 144900
rect 352190 144888 352196 144900
rect 352064 144860 352196 144888
rect 352064 144848 352070 144860
rect 352190 144848 352196 144860
rect 352248 144848 352254 144900
rect 353478 144848 353484 144900
rect 353536 144888 353542 144900
rect 353570 144888 353576 144900
rect 353536 144860 353576 144888
rect 353536 144848 353542 144860
rect 353570 144848 353576 144860
rect 353628 144848 353634 144900
rect 357526 144848 357532 144900
rect 357584 144888 357590 144900
rect 357710 144888 357716 144900
rect 357584 144860 357716 144888
rect 357584 144848 357590 144860
rect 357710 144848 357716 144860
rect 357768 144848 357774 144900
rect 358998 144848 359004 144900
rect 359056 144888 359062 144900
rect 359182 144888 359188 144900
rect 359056 144860 359188 144888
rect 359056 144848 359062 144860
rect 359182 144848 359188 144860
rect 359240 144848 359246 144900
rect 364518 144848 364524 144900
rect 364576 144888 364582 144900
rect 364610 144888 364616 144900
rect 364576 144860 364616 144888
rect 364576 144848 364582 144860
rect 364610 144848 364616 144860
rect 364668 144848 364674 144900
rect 370130 144848 370136 144900
rect 370188 144888 370194 144900
rect 370222 144888 370228 144900
rect 370188 144860 370228 144888
rect 370188 144848 370194 144860
rect 370222 144848 370228 144860
rect 370280 144848 370286 144900
rect 375558 144848 375564 144900
rect 375616 144888 375622 144900
rect 375650 144888 375656 144900
rect 375616 144860 375656 144888
rect 375616 144848 375622 144860
rect 375650 144848 375656 144860
rect 375708 144848 375714 144900
rect 400490 144888 400496 144900
rect 400451 144860 400496 144888
rect 400490 144848 400496 144860
rect 400548 144848 400554 144900
rect 422386 144888 422392 144900
rect 422347 144860 422392 144888
rect 422386 144848 422392 144860
rect 422444 144848 422450 144900
rect 427722 144848 427728 144900
rect 427780 144888 427786 144900
rect 427998 144888 428004 144900
rect 427780 144860 428004 144888
rect 427780 144848 427786 144860
rect 427998 144848 428004 144860
rect 428056 144848 428062 144900
rect 466546 144888 466552 144900
rect 466507 144860 466552 144888
rect 466546 144848 466552 144860
rect 466604 144848 466610 144900
rect 381081 144823 381139 144829
rect 381081 144789 381093 144823
rect 381127 144820 381139 144823
rect 381170 144820 381176 144832
rect 381127 144792 381176 144820
rect 381127 144789 381139 144792
rect 381081 144783 381139 144789
rect 381170 144780 381176 144792
rect 381228 144780 381234 144832
rect 254118 143556 254124 143608
rect 254176 143596 254182 143608
rect 254397 143599 254455 143605
rect 254397 143596 254409 143599
rect 254176 143568 254409 143596
rect 254176 143556 254182 143568
rect 254397 143565 254409 143568
rect 254443 143565 254455 143599
rect 254397 143559 254455 143565
rect 397730 143556 397736 143608
rect 397788 143596 397794 143608
rect 397788 143568 397833 143596
rect 397788 143556 397794 143568
rect 252738 143488 252744 143540
rect 252796 143528 252802 143540
rect 252922 143528 252928 143540
rect 252796 143500 252928 143528
rect 252796 143488 252802 143500
rect 252922 143488 252928 143500
rect 252980 143488 252986 143540
rect 254210 143528 254216 143540
rect 254171 143500 254216 143528
rect 254210 143488 254216 143500
rect 254268 143488 254274 143540
rect 259641 143531 259699 143537
rect 259641 143497 259653 143531
rect 259687 143528 259699 143531
rect 259730 143528 259736 143540
rect 259687 143500 259736 143528
rect 259687 143497 259699 143500
rect 259641 143491 259699 143497
rect 259730 143488 259736 143500
rect 259788 143488 259794 143540
rect 266446 143488 266452 143540
rect 266504 143528 266510 143540
rect 266722 143528 266728 143540
rect 266504 143500 266728 143528
rect 266504 143488 266510 143500
rect 266722 143488 266728 143500
rect 266780 143488 266786 143540
rect 287238 143528 287244 143540
rect 287199 143500 287244 143528
rect 287238 143488 287244 143500
rect 287296 143488 287302 143540
rect 305086 143528 305092 143540
rect 305047 143500 305092 143528
rect 305086 143488 305092 143500
rect 305144 143488 305150 143540
rect 309410 143488 309416 143540
rect 309468 143528 309474 143540
rect 309686 143528 309692 143540
rect 309468 143500 309692 143528
rect 309468 143488 309474 143500
rect 309686 143488 309692 143500
rect 309744 143488 309750 143540
rect 321646 143528 321652 143540
rect 321607 143500 321652 143528
rect 321646 143488 321652 143500
rect 321704 143488 321710 143540
rect 393222 143528 393228 143540
rect 393183 143500 393228 143528
rect 393222 143488 393228 143500
rect 393280 143488 393286 143540
rect 480254 143488 480260 143540
rect 480312 143528 480318 143540
rect 480438 143528 480444 143540
rect 480312 143500 480444 143528
rect 480312 143488 480318 143500
rect 480438 143488 480444 143500
rect 480496 143488 480502 143540
rect 236362 143460 236368 143472
rect 236323 143432 236368 143460
rect 236362 143420 236368 143432
rect 236420 143420 236426 143472
rect 334434 142168 334440 142180
rect 334395 142140 334440 142168
rect 334434 142128 334440 142140
rect 334492 142128 334498 142180
rect 283006 142100 283012 142112
rect 282967 142072 283012 142100
rect 283006 142060 283012 142072
rect 283064 142060 283070 142112
rect 408862 140020 408868 140072
rect 408920 140060 408926 140072
rect 409046 140060 409052 140072
rect 408920 140032 409052 140060
rect 408920 140020 408926 140032
rect 409046 140020 409052 140032
rect 409104 140020 409110 140072
rect 277670 138088 277676 138100
rect 277596 138060 277676 138088
rect 277596 137964 277624 138060
rect 277670 138048 277676 138060
rect 277728 138048 277734 138100
rect 376938 137980 376944 138032
rect 376996 137980 377002 138032
rect 382458 137980 382464 138032
rect 382516 137980 382522 138032
rect 416866 137980 416872 138032
rect 416924 137980 416930 138032
rect 451550 137980 451556 138032
rect 451608 137980 451614 138032
rect 472066 137980 472072 138032
rect 472124 137980 472130 138032
rect 277578 137912 277584 137964
rect 277636 137912 277642 137964
rect 376956 137896 376984 137980
rect 382476 137896 382504 137980
rect 400490 137952 400496 137964
rect 400451 137924 400496 137952
rect 400490 137912 400496 137924
rect 400548 137912 400554 137964
rect 416774 137912 416780 137964
rect 416832 137952 416838 137964
rect 416884 137952 416912 137980
rect 422386 137952 422392 137964
rect 416832 137924 416912 137952
rect 422347 137924 422392 137952
rect 416832 137912 416838 137924
rect 422386 137912 422392 137924
rect 422444 137912 422450 137964
rect 451568 137952 451596 137980
rect 451734 137952 451740 137964
rect 451568 137924 451740 137952
rect 451734 137912 451740 137924
rect 451792 137912 451798 137964
rect 466546 137952 466552 137964
rect 466507 137924 466552 137952
rect 466546 137912 466552 137924
rect 466604 137912 466610 137964
rect 471974 137912 471980 137964
rect 472032 137952 472038 137964
rect 472084 137952 472112 137980
rect 472032 137924 472112 137952
rect 472032 137912 472038 137924
rect 376938 137844 376944 137896
rect 376996 137844 377002 137896
rect 382458 137844 382464 137896
rect 382516 137844 382522 137896
rect 292758 135300 292764 135312
rect 292719 135272 292764 135300
rect 292758 135260 292764 135272
rect 292816 135260 292822 135312
rect 365990 135300 365996 135312
rect 365916 135272 365996 135300
rect 365916 135244 365944 135272
rect 365990 135260 365996 135272
rect 366048 135260 366054 135312
rect 381078 135300 381084 135312
rect 381039 135272 381084 135300
rect 381078 135260 381084 135272
rect 381136 135260 381142 135312
rect 243078 135192 243084 135244
rect 243136 135232 243142 135244
rect 243262 135232 243268 135244
rect 243136 135204 243268 135232
rect 243136 135192 243142 135204
rect 243262 135192 243268 135204
rect 243320 135192 243326 135244
rect 271874 135192 271880 135244
rect 271932 135232 271938 135244
rect 271966 135232 271972 135244
rect 271932 135204 271972 135232
rect 271932 135192 271938 135204
rect 271966 135192 271972 135204
rect 272024 135192 272030 135244
rect 321646 135232 321652 135244
rect 321607 135204 321652 135232
rect 321646 135192 321652 135204
rect 321704 135192 321710 135244
rect 365898 135192 365904 135244
rect 365956 135192 365962 135244
rect 367370 135192 367376 135244
rect 367428 135232 367434 135244
rect 367554 135232 367560 135244
rect 367428 135204 367560 135232
rect 367428 135192 367434 135204
rect 367554 135192 367560 135204
rect 367612 135192 367618 135244
rect 298002 134104 298008 134156
rect 298060 134144 298066 134156
rect 301590 134144 301596 134156
rect 298060 134116 301596 134144
rect 298060 134104 298066 134116
rect 301590 134104 301596 134116
rect 301648 134104 301654 134156
rect 383654 134036 383660 134088
rect 383712 134076 383718 134088
rect 385218 134076 385224 134088
rect 383712 134048 385224 134076
rect 383712 134036 383718 134048
rect 385218 134036 385224 134048
rect 385276 134036 385282 134088
rect 287238 133940 287244 133952
rect 287199 133912 287244 133940
rect 287238 133900 287244 133912
rect 287296 133900 287302 133952
rect 305086 133940 305092 133952
rect 305047 133912 305092 133940
rect 305086 133900 305092 133912
rect 305144 133900 305150 133952
rect 393222 133940 393228 133952
rect 393183 133912 393228 133940
rect 393222 133900 393228 133912
rect 393280 133900 393286 133952
rect 521654 133900 521660 133952
rect 521712 133940 521718 133952
rect 526438 133940 526444 133952
rect 521712 133912 526444 133940
rect 521712 133900 521718 133912
rect 526438 133900 526444 133912
rect 526496 133900 526502 133952
rect 243262 133872 243268 133884
rect 243223 133844 243268 133872
rect 243262 133832 243268 133844
rect 243320 133832 243326 133884
rect 292758 133872 292764 133884
rect 292719 133844 292764 133872
rect 292758 133832 292764 133844
rect 292816 133832 292822 133884
rect 334434 133872 334440 133884
rect 334395 133844 334440 133872
rect 334434 133832 334440 133844
rect 334492 133832 334498 133884
rect 353478 133872 353484 133884
rect 353439 133844 353484 133872
rect 353478 133832 353484 133844
rect 353536 133832 353542 133884
rect 356422 133872 356428 133884
rect 356383 133844 356428 133872
rect 356422 133832 356428 133844
rect 356480 133832 356486 133884
rect 386598 133872 386604 133884
rect 386559 133844 386604 133872
rect 386598 133832 386604 133844
rect 386656 133832 386662 133884
rect 259641 133807 259699 133813
rect 259641 133773 259653 133807
rect 259687 133804 259699 133807
rect 259730 133804 259736 133816
rect 259687 133776 259736 133804
rect 259687 133773 259699 133776
rect 259641 133767 259699 133773
rect 259730 133764 259736 133776
rect 259788 133764 259794 133816
rect 283009 132515 283067 132521
rect 283009 132481 283021 132515
rect 283055 132512 283067 132515
rect 283098 132512 283104 132524
rect 283055 132484 283104 132512
rect 283055 132481 283067 132484
rect 283009 132475 283067 132481
rect 283098 132472 283104 132484
rect 283156 132472 283162 132524
rect 267185 132447 267243 132453
rect 267185 132413 267197 132447
rect 267231 132444 267243 132447
rect 267274 132444 267280 132456
rect 267231 132416 267280 132444
rect 267231 132413 267243 132416
rect 267185 132407 267243 132413
rect 267274 132404 267280 132416
rect 267332 132404 267338 132456
rect 330018 128432 330024 128444
rect 329944 128404 330024 128432
rect 233326 128324 233332 128376
rect 233384 128364 233390 128376
rect 233510 128364 233516 128376
rect 233384 128336 233516 128364
rect 233384 128324 233390 128336
rect 233510 128324 233516 128336
rect 233568 128324 233574 128376
rect 318886 128324 318892 128376
rect 318944 128364 318950 128376
rect 319070 128364 319076 128376
rect 318944 128336 319076 128364
rect 318944 128324 318950 128336
rect 319070 128324 319076 128336
rect 319128 128324 319134 128376
rect 329944 128308 329972 128404
rect 330018 128392 330024 128404
rect 330076 128392 330082 128444
rect 422294 128324 422300 128376
rect 422352 128364 422358 128376
rect 422478 128364 422484 128376
rect 422352 128336 422484 128364
rect 422352 128324 422358 128336
rect 422478 128324 422484 128336
rect 422536 128324 422542 128376
rect 451550 128324 451556 128376
rect 451608 128364 451614 128376
rect 451734 128364 451740 128376
rect 451608 128336 451740 128364
rect 451608 128324 451614 128336
rect 451734 128324 451740 128336
rect 451792 128324 451798 128376
rect 329926 128256 329932 128308
rect 329984 128256 329990 128308
rect 236270 125740 236276 125792
rect 236328 125740 236334 125792
rect 236288 125656 236316 125740
rect 304905 125715 304963 125721
rect 304905 125681 304917 125715
rect 304951 125712 304963 125715
rect 305086 125712 305092 125724
rect 304951 125684 305092 125712
rect 304951 125681 304963 125684
rect 304905 125675 304963 125681
rect 305086 125672 305092 125684
rect 305144 125672 305150 125724
rect 236270 125604 236276 125656
rect 236328 125604 236334 125656
rect 240134 125604 240140 125656
rect 240192 125644 240198 125656
rect 240318 125644 240324 125656
rect 240192 125616 240324 125644
rect 240192 125604 240198 125616
rect 240318 125604 240324 125616
rect 240376 125604 240382 125656
rect 347958 125604 347964 125656
rect 348016 125604 348022 125656
rect 364518 125604 364524 125656
rect 364576 125604 364582 125656
rect 365898 125604 365904 125656
rect 365956 125644 365962 125656
rect 365990 125644 365996 125656
rect 365956 125616 365996 125644
rect 365956 125604 365962 125616
rect 365990 125604 365996 125616
rect 366048 125604 366054 125656
rect 400490 125604 400496 125656
rect 400548 125644 400554 125656
rect 400582 125644 400588 125656
rect 400548 125616 400588 125644
rect 400548 125604 400554 125616
rect 400582 125604 400588 125616
rect 400640 125604 400646 125656
rect 270586 125536 270592 125588
rect 270644 125576 270650 125588
rect 270770 125576 270776 125588
rect 270644 125548 270776 125576
rect 270644 125536 270650 125548
rect 270770 125536 270776 125548
rect 270828 125536 270834 125588
rect 271966 125536 271972 125588
rect 272024 125576 272030 125588
rect 272058 125576 272064 125588
rect 272024 125548 272064 125576
rect 272024 125536 272030 125548
rect 272058 125536 272064 125548
rect 272116 125536 272122 125588
rect 292758 125576 292764 125588
rect 292719 125548 292764 125576
rect 292758 125536 292764 125548
rect 292816 125536 292822 125588
rect 310698 125576 310704 125588
rect 310659 125548 310704 125576
rect 310698 125536 310704 125548
rect 310756 125536 310762 125588
rect 342438 125536 342444 125588
rect 342496 125576 342502 125588
rect 342622 125576 342628 125588
rect 342496 125548 342628 125576
rect 342496 125536 342502 125548
rect 342622 125536 342628 125548
rect 342680 125536 342686 125588
rect 347976 125508 348004 125604
rect 348050 125508 348056 125520
rect 347976 125480 348056 125508
rect 348050 125468 348056 125480
rect 348108 125468 348114 125520
rect 364536 125508 364564 125604
rect 369946 125536 369952 125588
rect 370004 125576 370010 125588
rect 370130 125576 370136 125588
rect 370004 125548 370136 125576
rect 370004 125536 370010 125548
rect 370130 125536 370136 125548
rect 370188 125536 370194 125588
rect 371418 125536 371424 125588
rect 371476 125576 371482 125588
rect 371510 125576 371516 125588
rect 371476 125548 371516 125576
rect 371476 125536 371482 125548
rect 371510 125536 371516 125548
rect 371568 125536 371574 125588
rect 381170 125576 381176 125588
rect 381131 125548 381176 125576
rect 381170 125536 381176 125548
rect 381228 125536 381234 125588
rect 433610 125576 433616 125588
rect 433571 125548 433616 125576
rect 433610 125536 433616 125548
rect 433668 125536 433674 125588
rect 364610 125508 364616 125520
rect 364536 125480 364616 125508
rect 364610 125468 364616 125480
rect 364668 125468 364674 125520
rect 259730 124312 259736 124364
rect 259788 124312 259794 124364
rect 259748 124228 259776 124312
rect 243265 124219 243323 124225
rect 243265 124185 243277 124219
rect 243311 124216 243323 124219
rect 243354 124216 243360 124228
rect 243311 124188 243360 124216
rect 243311 124185 243323 124188
rect 243265 124179 243323 124185
rect 243354 124176 243360 124188
rect 243412 124176 243418 124228
rect 254210 124216 254216 124228
rect 254171 124188 254216 124216
rect 254210 124176 254216 124188
rect 254268 124176 254274 124228
rect 259730 124176 259736 124228
rect 259788 124176 259794 124228
rect 304902 124216 304908 124228
rect 304863 124188 304908 124216
rect 304902 124176 304908 124188
rect 304960 124176 304966 124228
rect 334434 124216 334440 124228
rect 334395 124188 334440 124216
rect 334434 124176 334440 124188
rect 334492 124176 334498 124228
rect 353481 124219 353539 124225
rect 353481 124185 353493 124219
rect 353527 124216 353539 124219
rect 353570 124216 353576 124228
rect 353527 124188 353576 124216
rect 353527 124185 353539 124188
rect 353481 124179 353539 124185
rect 353570 124176 353576 124188
rect 353628 124176 353634 124228
rect 356422 124216 356428 124228
rect 356383 124188 356428 124216
rect 356422 124176 356428 124188
rect 356480 124176 356486 124228
rect 397730 124176 397736 124228
rect 397788 124216 397794 124228
rect 397914 124216 397920 124228
rect 397788 124188 397920 124216
rect 397788 124176 397794 124188
rect 397914 124176 397920 124188
rect 397972 124176 397978 124228
rect 240134 124108 240140 124160
rect 240192 124148 240198 124160
rect 249978 124148 249984 124160
rect 240192 124120 240237 124148
rect 249939 124120 249984 124148
rect 240192 124108 240198 124120
rect 249978 124108 249984 124120
rect 250036 124108 250042 124160
rect 271966 124148 271972 124160
rect 271927 124120 271972 124148
rect 271966 124108 271972 124120
rect 272024 124108 272030 124160
rect 287149 124151 287207 124157
rect 287149 124117 287161 124151
rect 287195 124148 287207 124151
rect 287238 124148 287244 124160
rect 287195 124120 287244 124148
rect 287195 124117 287207 124120
rect 287149 124111 287207 124117
rect 287238 124108 287244 124120
rect 287296 124108 287302 124160
rect 292850 124148 292856 124160
rect 292811 124120 292856 124148
rect 292850 124108 292856 124120
rect 292908 124108 292914 124160
rect 295518 124108 295524 124160
rect 295576 124148 295582 124160
rect 295610 124148 295616 124160
rect 295576 124120 295616 124148
rect 295576 124108 295582 124120
rect 295610 124108 295616 124120
rect 295668 124108 295674 124160
rect 309502 124108 309508 124160
rect 309560 124148 309566 124160
rect 309560 124120 309640 124148
rect 309560 124108 309566 124120
rect 309318 123972 309324 124024
rect 309376 124012 309382 124024
rect 309612 124012 309640 124120
rect 327166 124108 327172 124160
rect 327224 124148 327230 124160
rect 327258 124148 327264 124160
rect 327224 124120 327264 124148
rect 327224 124108 327230 124120
rect 327258 124108 327264 124120
rect 327316 124108 327322 124160
rect 342622 124148 342628 124160
rect 342583 124120 342628 124148
rect 342622 124108 342628 124120
rect 342680 124108 342686 124160
rect 365898 124148 365904 124160
rect 365859 124120 365904 124148
rect 365898 124108 365904 124120
rect 365956 124108 365962 124160
rect 407758 124148 407764 124160
rect 407719 124120 407764 124148
rect 407758 124108 407764 124120
rect 407816 124108 407822 124160
rect 466638 124148 466644 124160
rect 466599 124120 466644 124148
rect 466638 124108 466644 124120
rect 466696 124108 466702 124160
rect 309376 123984 309640 124012
rect 309376 123972 309382 123984
rect 345934 123224 345940 123276
rect 345992 123264 345998 123276
rect 354582 123264 354588 123276
rect 345992 123236 354588 123264
rect 345992 123224 345998 123236
rect 354582 123224 354588 123236
rect 354640 123224 354646 123276
rect 454034 123020 454040 123072
rect 454092 123060 454098 123072
rect 458174 123060 458180 123072
rect 454092 123032 458180 123060
rect 454092 123020 454098 123032
rect 458174 123020 458180 123032
rect 458232 123020 458238 123072
rect 514570 123020 514576 123072
rect 514628 123060 514634 123072
rect 516870 123060 516876 123072
rect 514628 123032 516876 123060
rect 514628 123020 514634 123032
rect 516870 123020 516876 123032
rect 516928 123020 516934 123072
rect 475930 122952 475936 123004
rect 475988 122992 475994 123004
rect 478138 122992 478144 123004
rect 475988 122964 478144 122992
rect 475988 122952 475994 122964
rect 478138 122952 478144 122964
rect 478196 122952 478202 123004
rect 386601 122927 386659 122933
rect 386601 122893 386613 122927
rect 386647 122924 386659 122927
rect 386690 122924 386696 122936
rect 386647 122896 386696 122924
rect 386647 122893 386659 122896
rect 386601 122887 386659 122893
rect 386690 122884 386696 122896
rect 386748 122884 386754 122936
rect 425054 122884 425060 122936
rect 425112 122924 425118 122936
rect 434530 122924 434536 122936
rect 425112 122896 434536 122924
rect 425112 122884 425118 122896
rect 434530 122884 434536 122896
rect 434588 122884 434594 122936
rect 524230 122884 524236 122936
rect 524288 122924 524294 122936
rect 526438 122924 526444 122936
rect 524288 122896 526444 122924
rect 524288 122884 524294 122896
rect 526438 122884 526444 122896
rect 526496 122884 526502 122936
rect 266630 122816 266636 122868
rect 266688 122856 266694 122868
rect 266722 122856 266728 122868
rect 266688 122828 266728 122856
rect 266688 122816 266694 122828
rect 266722 122816 266728 122828
rect 266780 122816 266786 122868
rect 267182 122856 267188 122868
rect 267143 122828 267188 122856
rect 267182 122816 267188 122828
rect 267240 122816 267246 122868
rect 259730 122748 259736 122800
rect 259788 122788 259794 122800
rect 259822 122788 259828 122800
rect 259788 122760 259828 122788
rect 259788 122748 259794 122760
rect 259822 122748 259828 122760
rect 259880 122748 259886 122800
rect 327258 122788 327264 122800
rect 327219 122760 327264 122788
rect 327258 122748 327264 122760
rect 327316 122748 327322 122800
rect 2958 122204 2964 122256
rect 3016 122244 3022 122256
rect 6178 122244 6184 122256
rect 3016 122216 6184 122244
rect 3016 122204 3022 122216
rect 6178 122204 6184 122216
rect 6236 122204 6242 122256
rect 386598 121388 386604 121440
rect 386656 121428 386662 121440
rect 386877 121431 386935 121437
rect 386877 121428 386889 121431
rect 386656 121400 386889 121428
rect 386656 121388 386662 121400
rect 386877 121397 386889 121400
rect 386923 121397 386935 121431
rect 386877 121391 386935 121397
rect 265066 120708 265072 120760
rect 265124 120748 265130 120760
rect 265250 120748 265256 120760
rect 265124 120720 265256 120748
rect 265124 120708 265130 120720
rect 265250 120708 265256 120720
rect 265308 120708 265314 120760
rect 329926 120232 329932 120284
rect 329984 120272 329990 120284
rect 330021 120275 330079 120281
rect 330021 120272 330033 120275
rect 329984 120244 330033 120272
rect 329984 120232 329990 120244
rect 330021 120241 330033 120244
rect 330067 120241 330079 120275
rect 330021 120235 330079 120241
rect 252554 119348 252560 119400
rect 252612 119388 252618 119400
rect 252741 119391 252799 119397
rect 252741 119388 252753 119391
rect 252612 119360 252753 119388
rect 252612 119348 252618 119360
rect 252741 119357 252753 119360
rect 252787 119357 252799 119391
rect 252741 119351 252799 119357
rect 321738 118844 321744 118856
rect 321699 118816 321744 118844
rect 321738 118804 321744 118816
rect 321796 118804 321802 118856
rect 324498 118844 324504 118856
rect 324459 118816 324504 118844
rect 324498 118804 324504 118816
rect 324556 118804 324562 118856
rect 298189 118779 298247 118785
rect 298189 118745 298201 118779
rect 298235 118776 298247 118779
rect 298278 118776 298284 118788
rect 298235 118748 298284 118776
rect 298235 118745 298247 118748
rect 298189 118739 298247 118745
rect 298278 118736 298284 118748
rect 298336 118736 298342 118788
rect 357618 118736 357624 118788
rect 357676 118736 357682 118788
rect 451734 118736 451740 118788
rect 451792 118736 451798 118788
rect 231854 118668 231860 118720
rect 231912 118708 231918 118720
rect 232038 118708 232044 118720
rect 231912 118680 232044 118708
rect 231912 118668 231918 118680
rect 232038 118668 232044 118680
rect 232096 118668 232102 118720
rect 244366 118668 244372 118720
rect 244424 118708 244430 118720
rect 244424 118680 244504 118708
rect 244424 118668 244430 118680
rect 244476 118652 244504 118680
rect 308122 118668 308128 118720
rect 308180 118668 308186 118720
rect 332778 118668 332784 118720
rect 332836 118668 332842 118720
rect 336826 118668 336832 118720
rect 336884 118668 336890 118720
rect 346578 118668 346584 118720
rect 346636 118668 346642 118720
rect 244458 118600 244464 118652
rect 244516 118600 244522 118652
rect 308140 118584 308168 118668
rect 310698 118640 310704 118652
rect 310659 118612 310704 118640
rect 310698 118600 310704 118612
rect 310756 118600 310762 118652
rect 332796 118584 332824 118668
rect 336844 118584 336872 118668
rect 346596 118584 346624 118668
rect 357636 118652 357664 118736
rect 416866 118668 416872 118720
rect 416924 118668 416930 118720
rect 422386 118668 422392 118720
rect 422444 118668 422450 118720
rect 357618 118600 357624 118652
rect 357676 118600 357682 118652
rect 365898 118640 365904 118652
rect 365859 118612 365904 118640
rect 365898 118600 365904 118612
rect 365956 118600 365962 118652
rect 416774 118600 416780 118652
rect 416832 118640 416838 118652
rect 416884 118640 416912 118668
rect 416832 118612 416912 118640
rect 422404 118640 422432 118668
rect 451752 118652 451780 118736
rect 472066 118668 472072 118720
rect 472124 118668 472130 118720
rect 422478 118640 422484 118652
rect 422404 118612 422484 118640
rect 416832 118600 416838 118612
rect 422478 118600 422484 118612
rect 422536 118600 422542 118652
rect 451734 118600 451740 118652
rect 451792 118600 451798 118652
rect 471974 118600 471980 118652
rect 472032 118640 472038 118652
rect 472084 118640 472112 118668
rect 472032 118612 472112 118640
rect 472032 118600 472038 118612
rect 308122 118532 308128 118584
rect 308180 118532 308186 118584
rect 332778 118532 332784 118584
rect 332836 118532 332842 118584
rect 336826 118532 336832 118584
rect 336884 118532 336890 118584
rect 346578 118532 346584 118584
rect 346636 118532 346642 118584
rect 236270 117988 236276 118040
rect 236328 118028 236334 118040
rect 236454 118028 236460 118040
rect 236328 118000 236460 118028
rect 236328 117988 236334 118000
rect 236454 117988 236460 118000
rect 236512 117988 236518 118040
rect 266906 117784 266912 117836
rect 266964 117824 266970 117836
rect 267182 117824 267188 117836
rect 266964 117796 267188 117824
rect 266964 117784 266970 117796
rect 267182 117784 267188 117796
rect 267240 117784 267246 117836
rect 381170 115988 381176 116000
rect 381131 115960 381176 115988
rect 381170 115948 381176 115960
rect 381228 115948 381234 116000
rect 400398 115948 400404 116000
rect 400456 115988 400462 116000
rect 400490 115988 400496 116000
rect 400456 115960 400496 115988
rect 400456 115948 400462 115960
rect 400490 115948 400496 115960
rect 400548 115948 400554 116000
rect 433610 115988 433616 116000
rect 433571 115960 433616 115988
rect 433610 115948 433616 115960
rect 433668 115948 433674 116000
rect 254118 115880 254124 115932
rect 254176 115920 254182 115932
rect 254210 115920 254216 115932
rect 254176 115892 254216 115920
rect 254176 115880 254182 115892
rect 254210 115880 254216 115892
rect 254268 115880 254274 115932
rect 277486 115880 277492 115932
rect 277544 115920 277550 115932
rect 277670 115920 277676 115932
rect 277544 115892 277676 115920
rect 277544 115880 277550 115892
rect 277670 115880 277676 115892
rect 277728 115880 277734 115932
rect 305086 115920 305092 115932
rect 305047 115892 305092 115920
rect 305086 115880 305092 115892
rect 305144 115880 305150 115932
rect 271966 115376 271972 115388
rect 271927 115348 271972 115376
rect 271966 115336 271972 115348
rect 272024 115336 272030 115388
rect 393222 114656 393228 114708
rect 393280 114656 393286 114708
rect 294046 114588 294052 114640
rect 294104 114588 294110 114640
rect 353570 114628 353576 114640
rect 353496 114600 353576 114628
rect 240137 114563 240195 114569
rect 240137 114529 240149 114563
rect 240183 114560 240195 114563
rect 240226 114560 240232 114572
rect 240183 114532 240232 114560
rect 240183 114529 240195 114532
rect 240137 114523 240195 114529
rect 240226 114520 240232 114532
rect 240284 114520 240290 114572
rect 243170 114520 243176 114572
rect 243228 114560 243234 114572
rect 243354 114560 243360 114572
rect 243228 114532 243360 114560
rect 243228 114520 243234 114532
rect 243354 114520 243360 114532
rect 243412 114520 243418 114572
rect 249978 114560 249984 114572
rect 249939 114532 249984 114560
rect 249978 114520 249984 114532
rect 250036 114520 250042 114572
rect 283098 114520 283104 114572
rect 283156 114560 283162 114572
rect 283190 114560 283196 114572
rect 283156 114532 283196 114560
rect 283156 114520 283162 114532
rect 283190 114520 283196 114532
rect 283248 114520 283254 114572
rect 287146 114560 287152 114572
rect 287107 114532 287152 114560
rect 287146 114520 287152 114532
rect 287204 114520 287210 114572
rect 294064 114560 294092 114588
rect 353496 114572 353524 114600
rect 353570 114588 353576 114600
rect 353628 114588 353634 114640
rect 356422 114588 356428 114640
rect 356480 114588 356486 114640
rect 369946 114588 369952 114640
rect 370004 114628 370010 114640
rect 370004 114600 370084 114628
rect 370004 114588 370010 114600
rect 294138 114560 294144 114572
rect 294064 114532 294144 114560
rect 294138 114520 294144 114532
rect 294196 114520 294202 114572
rect 321738 114560 321744 114572
rect 321699 114532 321744 114560
rect 321738 114520 321744 114532
rect 321796 114520 321802 114572
rect 324498 114560 324504 114572
rect 324459 114532 324504 114560
rect 324498 114520 324504 114532
rect 324556 114520 324562 114572
rect 342622 114560 342628 114572
rect 342583 114532 342628 114560
rect 342622 114520 342628 114532
rect 342680 114520 342686 114572
rect 348050 114560 348056 114572
rect 348011 114532 348056 114560
rect 348050 114520 348056 114532
rect 348108 114520 348114 114572
rect 353478 114520 353484 114572
rect 353536 114520 353542 114572
rect 356440 114560 356468 114588
rect 370056 114572 370084 114600
rect 393240 114572 393268 114656
rect 408586 114588 408592 114640
rect 408644 114628 408650 114640
rect 408770 114628 408776 114640
rect 408644 114600 408776 114628
rect 408644 114588 408650 114600
rect 408770 114588 408776 114600
rect 408828 114588 408834 114640
rect 356514 114560 356520 114572
rect 356440 114532 356520 114560
rect 356514 114520 356520 114532
rect 356572 114520 356578 114572
rect 370038 114520 370044 114572
rect 370096 114520 370102 114572
rect 393222 114520 393228 114572
rect 393280 114520 393286 114572
rect 407758 114560 407764 114572
rect 407719 114532 407764 114560
rect 407758 114520 407764 114532
rect 407816 114520 407822 114572
rect 466641 114563 466699 114569
rect 466641 114529 466653 114563
rect 466687 114560 466699 114563
rect 466822 114560 466828 114572
rect 466687 114532 466828 114560
rect 466687 114529 466699 114532
rect 466641 114523 466699 114529
rect 466822 114520 466828 114532
rect 466880 114520 466886 114572
rect 254118 114452 254124 114504
rect 254176 114492 254182 114504
rect 254210 114492 254216 114504
rect 254176 114464 254216 114492
rect 254176 114452 254182 114464
rect 254210 114452 254216 114464
rect 254268 114452 254274 114504
rect 397641 114495 397699 114501
rect 397641 114461 397653 114495
rect 397687 114492 397699 114495
rect 397730 114492 397736 114504
rect 397687 114464 397736 114492
rect 397687 114461 397699 114464
rect 397641 114455 397699 114461
rect 397730 114452 397736 114464
rect 397788 114452 397794 114504
rect 408681 114495 408739 114501
rect 408681 114461 408693 114495
rect 408727 114492 408739 114495
rect 408770 114492 408776 114504
rect 408727 114464 408776 114492
rect 408727 114461 408739 114464
rect 408681 114455 408739 114461
rect 408770 114452 408776 114464
rect 408828 114452 408834 114504
rect 292853 113203 292911 113209
rect 292853 113169 292865 113203
rect 292899 113200 292911 113203
rect 292942 113200 292948 113212
rect 292899 113172 292948 113200
rect 292899 113169 292911 113172
rect 292853 113163 292911 113169
rect 292942 113160 292948 113172
rect 293000 113160 293006 113212
rect 327258 113200 327264 113212
rect 327219 113172 327264 113200
rect 327258 113160 327264 113172
rect 327316 113160 327322 113212
rect 348050 113200 348056 113212
rect 348011 113172 348056 113200
rect 348050 113160 348056 113172
rect 348108 113160 348114 113212
rect 236273 113135 236331 113141
rect 236273 113101 236285 113135
rect 236319 113132 236331 113135
rect 236362 113132 236368 113144
rect 236319 113104 236368 113132
rect 236319 113101 236331 113104
rect 236273 113095 236331 113101
rect 236362 113092 236368 113104
rect 236420 113092 236426 113144
rect 295518 113132 295524 113144
rect 295479 113104 295524 113132
rect 295518 113092 295524 113104
rect 295576 113092 295582 113144
rect 298189 111843 298247 111849
rect 298189 111809 298201 111843
rect 298235 111809 298247 111843
rect 298189 111803 298247 111809
rect 298204 111704 298232 111803
rect 298373 111707 298431 111713
rect 298373 111704 298385 111707
rect 298204 111676 298385 111704
rect 298373 111673 298385 111676
rect 298419 111673 298431 111707
rect 298373 111667 298431 111673
rect 336734 110712 336740 110764
rect 336792 110752 336798 110764
rect 346210 110752 346216 110764
rect 336792 110724 346216 110752
rect 336792 110712 336798 110724
rect 346210 110712 346216 110724
rect 346268 110712 346274 110764
rect 425054 110508 425060 110560
rect 425112 110548 425118 110560
rect 434530 110548 434536 110560
rect 425112 110520 434536 110548
rect 425112 110508 425118 110520
rect 434530 110508 434536 110520
rect 434588 110508 434594 110560
rect 521654 110508 521660 110560
rect 521712 110548 521718 110560
rect 526438 110548 526444 110560
rect 521712 110520 526444 110548
rect 521712 110508 521718 110520
rect 526438 110508 526444 110520
rect 526496 110508 526502 110560
rect 243078 109732 243084 109744
rect 243039 109704 243084 109732
rect 243078 109692 243084 109704
rect 243136 109692 243142 109744
rect 282914 109692 282920 109744
rect 282972 109732 282978 109744
rect 283098 109732 283104 109744
rect 282972 109704 283104 109732
rect 282972 109692 282978 109704
rect 283098 109692 283104 109704
rect 283156 109692 283162 109744
rect 294138 109692 294144 109744
rect 294196 109692 294202 109744
rect 294156 109608 294184 109692
rect 294138 109556 294144 109608
rect 294196 109556 294202 109608
rect 364518 109080 364524 109132
rect 364576 109120 364582 109132
rect 364702 109120 364708 109132
rect 364576 109092 364708 109120
rect 364576 109080 364582 109092
rect 364702 109080 364708 109092
rect 364760 109080 364766 109132
rect 233326 109012 233332 109064
rect 233384 109052 233390 109064
rect 233510 109052 233516 109064
rect 233384 109024 233516 109052
rect 233384 109012 233390 109024
rect 233510 109012 233516 109024
rect 233568 109012 233574 109064
rect 422294 109012 422300 109064
rect 422352 109052 422358 109064
rect 422478 109052 422484 109064
rect 422352 109024 422484 109052
rect 422352 109012 422358 109024
rect 422478 109012 422484 109024
rect 422536 109012 422542 109064
rect 252738 106332 252744 106344
rect 252699 106304 252744 106332
rect 252738 106292 252744 106304
rect 252796 106292 252802 106344
rect 305089 106335 305147 106341
rect 305089 106301 305101 106335
rect 305135 106332 305147 106335
rect 305178 106332 305184 106344
rect 305135 106304 305184 106332
rect 305135 106301 305147 106304
rect 305089 106295 305147 106301
rect 305178 106292 305184 106304
rect 305236 106292 305242 106344
rect 319070 106292 319076 106344
rect 319128 106292 319134 106344
rect 330018 106332 330024 106344
rect 329979 106304 330024 106332
rect 330018 106292 330024 106304
rect 330076 106292 330082 106344
rect 342530 106292 342536 106344
rect 342588 106332 342594 106344
rect 342622 106332 342628 106344
rect 342588 106304 342628 106332
rect 342588 106292 342594 106304
rect 342622 106292 342628 106304
rect 342680 106292 342686 106344
rect 370038 106292 370044 106344
rect 370096 106292 370102 106344
rect 240137 106267 240195 106273
rect 240137 106233 240149 106267
rect 240183 106264 240195 106267
rect 240226 106264 240232 106276
rect 240183 106236 240232 106264
rect 240183 106233 240195 106236
rect 240137 106227 240195 106233
rect 240226 106224 240232 106236
rect 240284 106224 240290 106276
rect 241790 106224 241796 106276
rect 241848 106264 241854 106276
rect 241974 106264 241980 106276
rect 241848 106236 241980 106264
rect 241848 106224 241854 106236
rect 241974 106224 241980 106236
rect 242032 106224 242038 106276
rect 281626 106264 281632 106276
rect 281587 106236 281632 106264
rect 281626 106224 281632 106236
rect 281684 106224 281690 106276
rect 309226 106224 309232 106276
rect 309284 106264 309290 106276
rect 309318 106264 309324 106276
rect 309284 106236 309324 106264
rect 309284 106224 309290 106236
rect 309318 106224 309324 106236
rect 309376 106224 309382 106276
rect 319088 106208 319116 106292
rect 324498 106264 324504 106276
rect 324459 106236 324504 106264
rect 324498 106224 324504 106236
rect 324556 106224 324562 106276
rect 357618 106264 357624 106276
rect 357579 106236 357624 106264
rect 357618 106224 357624 106236
rect 357676 106224 357682 106276
rect 243081 106199 243139 106205
rect 243081 106165 243093 106199
rect 243127 106196 243139 106199
rect 243262 106196 243268 106208
rect 243127 106168 243268 106196
rect 243127 106165 243139 106168
rect 243081 106159 243139 106165
rect 243262 106156 243268 106168
rect 243320 106156 243326 106208
rect 319070 106156 319076 106208
rect 319128 106156 319134 106208
rect 370056 106196 370084 106292
rect 392026 106224 392032 106276
rect 392084 106264 392090 106276
rect 392302 106264 392308 106276
rect 392084 106236 392308 106264
rect 392084 106224 392090 106236
rect 392302 106224 392308 106236
rect 392360 106224 392366 106276
rect 422386 106264 422392 106276
rect 422347 106236 422392 106264
rect 422386 106224 422392 106236
rect 422444 106224 422450 106276
rect 427906 106264 427912 106276
rect 427867 106236 427912 106264
rect 427906 106224 427912 106236
rect 427964 106224 427970 106276
rect 433610 106264 433616 106276
rect 433571 106236 433616 106264
rect 433610 106224 433616 106236
rect 433668 106224 433674 106276
rect 370130 106196 370136 106208
rect 370056 106168 370136 106196
rect 370130 106156 370136 106168
rect 370188 106156 370194 106208
rect 327258 104972 327264 104984
rect 327184 104944 327264 104972
rect 327184 104916 327212 104944
rect 327258 104932 327264 104944
rect 327316 104932 327322 104984
rect 397638 104972 397644 104984
rect 397599 104944 397644 104972
rect 397638 104932 397644 104944
rect 397696 104932 397702 104984
rect 271874 104864 271880 104916
rect 271932 104904 271938 104916
rect 271966 104904 271972 104916
rect 271932 104876 271972 104904
rect 271932 104864 271938 104876
rect 271966 104864 271972 104876
rect 272024 104864 272030 104916
rect 292758 104864 292764 104916
rect 292816 104904 292822 104916
rect 292942 104904 292948 104916
rect 292816 104876 292948 104904
rect 292816 104864 292822 104876
rect 292942 104864 292948 104876
rect 293000 104864 293006 104916
rect 327166 104864 327172 104916
rect 327224 104864 327230 104916
rect 347866 104864 347872 104916
rect 347924 104904 347930 104916
rect 348050 104904 348056 104916
rect 347924 104876 348056 104904
rect 347924 104864 347930 104876
rect 348050 104864 348056 104876
rect 348108 104864 348114 104916
rect 408678 104904 408684 104916
rect 408639 104876 408684 104904
rect 408678 104864 408684 104876
rect 408736 104864 408742 104916
rect 282914 104836 282920 104848
rect 282875 104808 282920 104836
rect 282914 104796 282920 104808
rect 282972 104796 282978 104848
rect 309226 104836 309232 104848
rect 309187 104808 309232 104836
rect 309226 104796 309232 104808
rect 309284 104796 309290 104848
rect 319070 104836 319076 104848
rect 319031 104808 319076 104836
rect 319070 104796 319076 104808
rect 319128 104796 319134 104848
rect 393133 104839 393191 104845
rect 393133 104805 393145 104839
rect 393179 104836 393191 104839
rect 393222 104836 393228 104848
rect 393179 104808 393228 104836
rect 393179 104805 393191 104808
rect 393133 104799 393191 104805
rect 393222 104796 393228 104808
rect 393280 104796 393286 104848
rect 397638 104796 397644 104848
rect 397696 104796 397702 104848
rect 400490 104836 400496 104848
rect 400451 104808 400496 104836
rect 400490 104796 400496 104808
rect 400548 104796 400554 104848
rect 407758 104836 407764 104848
rect 407719 104808 407764 104836
rect 407758 104796 407764 104808
rect 407816 104796 407822 104848
rect 480438 104836 480444 104848
rect 480399 104808 480444 104836
rect 480438 104796 480444 104808
rect 480496 104796 480502 104848
rect 397656 104768 397684 104796
rect 397822 104768 397828 104780
rect 397656 104740 397828 104768
rect 397822 104728 397828 104740
rect 397880 104728 397886 104780
rect 364518 103708 364524 103760
rect 364576 103748 364582 103760
rect 364702 103748 364708 103760
rect 364576 103720 364708 103748
rect 364576 103708 364582 103720
rect 364702 103708 364708 103720
rect 364760 103708 364766 103760
rect 236270 103544 236276 103556
rect 236231 103516 236276 103544
rect 236270 103504 236276 103516
rect 236328 103504 236334 103556
rect 295518 103544 295524 103556
rect 295479 103516 295524 103544
rect 295518 103504 295524 103516
rect 295576 103504 295582 103556
rect 386874 103504 386880 103556
rect 386932 103544 386938 103556
rect 386932 103516 386977 103544
rect 386932 103504 386938 103516
rect 254210 103476 254216 103488
rect 254171 103448 254216 103476
rect 254210 103436 254216 103448
rect 254268 103436 254274 103488
rect 353481 103479 353539 103485
rect 353481 103445 353493 103479
rect 353527 103476 353539 103479
rect 353570 103476 353576 103488
rect 353527 103448 353576 103476
rect 353527 103445 353539 103448
rect 353481 103439 353539 103445
rect 353570 103436 353576 103448
rect 353628 103436 353634 103488
rect 356606 103436 356612 103488
rect 356664 103436 356670 103488
rect 370130 103436 370136 103488
rect 370188 103476 370194 103488
rect 370314 103476 370320 103488
rect 370188 103448 370320 103476
rect 370188 103436 370194 103448
rect 370314 103436 370320 103448
rect 370372 103436 370378 103488
rect 356422 103368 356428 103420
rect 356480 103408 356486 103420
rect 356624 103408 356652 103436
rect 356480 103380 356652 103408
rect 356480 103368 356486 103380
rect 236270 103096 236276 103148
rect 236328 103136 236334 103148
rect 236454 103136 236460 103148
rect 236328 103108 236460 103136
rect 236328 103096 236334 103108
rect 236454 103096 236460 103108
rect 236512 103096 236518 103148
rect 298370 102184 298376 102196
rect 298331 102156 298376 102184
rect 298370 102144 298376 102156
rect 298428 102144 298434 102196
rect 266449 102119 266507 102125
rect 266449 102085 266461 102119
rect 266495 102116 266507 102119
rect 266538 102116 266544 102128
rect 266495 102088 266544 102116
rect 266495 102085 266507 102088
rect 266449 102079 266507 102085
rect 266538 102076 266544 102088
rect 266596 102076 266602 102128
rect 231854 101396 231860 101448
rect 231912 101436 231918 101448
rect 232038 101436 232044 101448
rect 231912 101408 232044 101436
rect 231912 101396 231918 101408
rect 232038 101396 232044 101408
rect 232096 101396 232102 101448
rect 281626 101368 281632 101380
rect 281587 101340 281632 101368
rect 281626 101328 281632 101340
rect 281684 101328 281690 101380
rect 408770 100076 408776 100088
rect 408731 100048 408776 100076
rect 408770 100036 408776 100048
rect 408828 100036 408834 100088
rect 244458 99424 244464 99476
rect 244516 99424 244522 99476
rect 277578 99424 277584 99476
rect 277636 99424 277642 99476
rect 298370 99464 298376 99476
rect 298331 99436 298376 99464
rect 298370 99424 298376 99436
rect 298428 99424 298434 99476
rect 244476 99340 244504 99424
rect 277596 99340 277624 99424
rect 288618 99396 288624 99408
rect 288579 99368 288624 99396
rect 288618 99356 288624 99368
rect 288676 99356 288682 99408
rect 308122 99396 308128 99408
rect 308083 99368 308128 99396
rect 308122 99356 308128 99368
rect 308180 99356 308186 99408
rect 310698 99396 310704 99408
rect 310659 99368 310704 99396
rect 310698 99356 310704 99368
rect 310756 99356 310762 99408
rect 416866 99356 416872 99408
rect 416924 99356 416930 99408
rect 472066 99356 472072 99408
rect 472124 99356 472130 99408
rect 244458 99288 244464 99340
rect 244516 99288 244522 99340
rect 271874 99288 271880 99340
rect 271932 99328 271938 99340
rect 272058 99328 272064 99340
rect 271932 99300 272064 99328
rect 271932 99288 271938 99300
rect 272058 99288 272064 99300
rect 272116 99288 272122 99340
rect 277578 99288 277584 99340
rect 277636 99288 277642 99340
rect 416774 99288 416780 99340
rect 416832 99328 416838 99340
rect 416884 99328 416912 99356
rect 422386 99328 422392 99340
rect 416832 99300 416912 99328
rect 422347 99300 422392 99328
rect 416832 99288 416838 99300
rect 422386 99288 422392 99300
rect 422444 99288 422450 99340
rect 427906 99328 427912 99340
rect 427867 99300 427912 99328
rect 427906 99288 427912 99300
rect 427964 99288 427970 99340
rect 433610 99328 433616 99340
rect 433571 99300 433616 99328
rect 433610 99288 433616 99300
rect 433668 99288 433674 99340
rect 471974 99288 471980 99340
rect 472032 99328 472038 99340
rect 472084 99328 472112 99356
rect 472032 99300 472112 99328
rect 472032 99288 472038 99300
rect 393130 98716 393136 98728
rect 393091 98688 393136 98716
rect 393130 98676 393136 98688
rect 393188 98676 393194 98728
rect 240134 96676 240140 96688
rect 240095 96648 240140 96676
rect 240134 96636 240140 96648
rect 240192 96636 240198 96688
rect 288618 96676 288624 96688
rect 288579 96648 288624 96676
rect 288618 96636 288624 96648
rect 288676 96636 288682 96688
rect 308122 96676 308128 96688
rect 308083 96648 308128 96676
rect 308122 96636 308128 96648
rect 308180 96636 308186 96688
rect 310698 96676 310704 96688
rect 310659 96648 310704 96676
rect 310698 96636 310704 96648
rect 310756 96636 310762 96688
rect 324498 96676 324504 96688
rect 324459 96648 324504 96676
rect 324498 96636 324504 96648
rect 324556 96636 324562 96688
rect 357621 96543 357679 96549
rect 357621 96509 357633 96543
rect 357667 96540 357679 96543
rect 357710 96540 357716 96552
rect 357667 96512 357716 96540
rect 357667 96509 357679 96512
rect 357621 96503 357679 96509
rect 357710 96500 357716 96512
rect 357768 96500 357774 96552
rect 259638 95208 259644 95260
rect 259696 95248 259702 95260
rect 259822 95248 259828 95260
rect 259696 95220 259828 95248
rect 259696 95208 259702 95220
rect 259822 95208 259828 95220
rect 259880 95208 259886 95260
rect 266906 95208 266912 95260
rect 266964 95248 266970 95260
rect 267090 95248 267096 95260
rect 266964 95220 267096 95248
rect 266964 95208 266970 95220
rect 267090 95208 267096 95220
rect 267148 95208 267154 95260
rect 282914 95248 282920 95260
rect 282875 95220 282920 95248
rect 282914 95208 282920 95220
rect 282972 95208 282978 95260
rect 295518 95208 295524 95260
rect 295576 95208 295582 95260
rect 319070 95248 319076 95260
rect 319031 95220 319076 95248
rect 319070 95208 319076 95220
rect 319128 95208 319134 95260
rect 327166 95208 327172 95260
rect 327224 95248 327230 95260
rect 327258 95248 327264 95260
rect 327224 95220 327264 95248
rect 327224 95208 327230 95220
rect 327258 95208 327264 95220
rect 327316 95208 327322 95260
rect 400493 95251 400551 95257
rect 400493 95217 400505 95251
rect 400539 95248 400551 95251
rect 400582 95248 400588 95260
rect 400539 95220 400588 95248
rect 400539 95217 400551 95220
rect 400493 95211 400551 95217
rect 400582 95208 400588 95220
rect 400640 95208 400646 95260
rect 466546 95208 466552 95260
rect 466604 95248 466610 95260
rect 466822 95248 466828 95260
rect 466604 95220 466828 95248
rect 466604 95208 466610 95220
rect 466822 95208 466828 95220
rect 466880 95208 466886 95260
rect 480441 95251 480499 95257
rect 480441 95217 480453 95251
rect 480487 95248 480499 95251
rect 480530 95248 480536 95260
rect 480487 95220 480536 95248
rect 480487 95217 480499 95220
rect 480441 95211 480499 95217
rect 480530 95208 480536 95220
rect 480588 95208 480594 95260
rect 236273 95183 236331 95189
rect 236273 95149 236285 95183
rect 236319 95180 236331 95183
rect 236362 95180 236368 95192
rect 236319 95152 236368 95180
rect 236319 95149 236331 95152
rect 236273 95143 236331 95149
rect 236362 95140 236368 95152
rect 236420 95140 236426 95192
rect 240134 95140 240140 95192
rect 240192 95180 240198 95192
rect 287149 95183 287207 95189
rect 240192 95152 240237 95180
rect 240192 95140 240198 95152
rect 287149 95149 287161 95183
rect 287195 95180 287207 95183
rect 287238 95180 287244 95192
rect 287195 95152 287244 95180
rect 287195 95149 287207 95152
rect 287149 95143 287207 95149
rect 287238 95140 287244 95152
rect 287296 95140 287302 95192
rect 295536 95112 295564 95208
rect 295610 95112 295616 95124
rect 295536 95084 295616 95112
rect 295610 95072 295616 95084
rect 295668 95072 295674 95124
rect 351822 95072 351828 95124
rect 351880 95112 351886 95124
rect 352190 95112 352196 95124
rect 351880 95084 352196 95112
rect 351880 95072 351886 95084
rect 352190 95072 352196 95084
rect 352248 95072 352254 95124
rect 386782 93916 386788 93968
rect 386840 93956 386846 93968
rect 386840 93928 386920 93956
rect 386840 93916 386846 93928
rect 386892 93900 386920 93928
rect 254210 93888 254216 93900
rect 254171 93860 254216 93888
rect 254210 93848 254216 93860
rect 254268 93848 254274 93900
rect 353478 93888 353484 93900
rect 353439 93860 353484 93888
rect 353478 93848 353484 93860
rect 353536 93848 353542 93900
rect 386874 93848 386880 93900
rect 386932 93848 386938 93900
rect 294138 93780 294144 93832
rect 294196 93780 294202 93832
rect 298370 93820 298376 93832
rect 298331 93792 298376 93820
rect 298370 93780 298376 93792
rect 298428 93780 298434 93832
rect 364521 93823 364579 93829
rect 364521 93789 364533 93823
rect 364567 93820 364579 93823
rect 364702 93820 364708 93832
rect 364567 93792 364708 93820
rect 364567 93789 364579 93792
rect 364521 93783 364579 93789
rect 364702 93780 364708 93792
rect 364760 93780 364766 93832
rect 294156 93693 294184 93780
rect 294141 93687 294199 93693
rect 294141 93653 294153 93687
rect 294187 93653 294199 93687
rect 294141 93647 294199 93653
rect 375558 93548 375564 93560
rect 375519 93520 375564 93548
rect 375558 93508 375564 93520
rect 375616 93508 375622 93560
rect 266446 92528 266452 92540
rect 266407 92500 266452 92528
rect 266446 92488 266452 92500
rect 266504 92488 266510 92540
rect 242986 91740 242992 91792
rect 243044 91780 243050 91792
rect 243446 91780 243452 91792
rect 243044 91752 243452 91780
rect 243044 91740 243050 91752
rect 243446 91740 243452 91752
rect 243504 91740 243510 91792
rect 342438 89768 342444 89820
rect 342496 89768 342502 89820
rect 380989 89811 381047 89817
rect 380989 89777 381001 89811
rect 381035 89808 381047 89811
rect 381078 89808 381084 89820
rect 381035 89780 381084 89808
rect 381035 89777 381047 89780
rect 380989 89771 381047 89777
rect 381078 89768 381084 89780
rect 381136 89768 381142 89820
rect 233326 89700 233332 89752
rect 233384 89740 233390 89752
rect 233510 89740 233516 89752
rect 233384 89712 233516 89740
rect 233384 89700 233390 89712
rect 233510 89700 233516 89712
rect 233568 89700 233574 89752
rect 259638 89700 259644 89752
rect 259696 89700 259702 89752
rect 259656 89604 259684 89700
rect 342456 89684 342484 89768
rect 356422 89700 356428 89752
rect 356480 89700 356486 89752
rect 422294 89700 422300 89752
rect 422352 89740 422358 89752
rect 422478 89740 422484 89752
rect 422352 89712 422484 89740
rect 422352 89700 422358 89712
rect 422478 89700 422484 89712
rect 422536 89700 422542 89752
rect 427814 89700 427820 89752
rect 427872 89740 427878 89752
rect 427998 89740 428004 89752
rect 427872 89712 428004 89740
rect 427872 89700 427878 89712
rect 427998 89700 428004 89712
rect 428056 89700 428062 89752
rect 309229 89675 309287 89681
rect 309229 89641 309241 89675
rect 309275 89672 309287 89675
rect 309318 89672 309324 89684
rect 309275 89644 309324 89672
rect 309275 89641 309287 89644
rect 309229 89635 309287 89641
rect 309318 89632 309324 89644
rect 309376 89632 309382 89684
rect 342438 89632 342444 89684
rect 342496 89632 342502 89684
rect 259730 89604 259736 89616
rect 259656 89576 259736 89604
rect 259730 89564 259736 89576
rect 259788 89564 259794 89616
rect 356440 89604 356468 89700
rect 358998 89632 359004 89684
rect 359056 89672 359062 89684
rect 359182 89672 359188 89684
rect 359056 89644 359188 89672
rect 359056 89632 359062 89644
rect 359182 89632 359188 89644
rect 359240 89632 359246 89684
rect 408770 89672 408776 89684
rect 408731 89644 408776 89672
rect 408770 89632 408776 89644
rect 408828 89632 408834 89684
rect 356514 89604 356520 89616
rect 356440 89576 356520 89604
rect 356514 89564 356520 89576
rect 356572 89564 356578 89616
rect 298370 88952 298376 89004
rect 298428 88992 298434 89004
rect 298557 88995 298615 89001
rect 298557 88992 298569 88995
rect 298428 88964 298569 88992
rect 298428 88952 298434 88964
rect 298557 88961 298569 88964
rect 298603 88961 298615 88995
rect 298557 88955 298615 88961
rect 365622 87184 365628 87236
rect 365680 87224 365686 87236
rect 373902 87224 373908 87236
rect 365680 87196 373908 87224
rect 365680 87184 365686 87196
rect 373902 87184 373908 87196
rect 373960 87184 373966 87236
rect 267734 87116 267740 87168
rect 267792 87156 267798 87168
rect 273714 87156 273720 87168
rect 267792 87128 273720 87156
rect 267792 87116 267798 87128
rect 273714 87116 273720 87128
rect 273772 87116 273778 87168
rect 328546 87116 328552 87168
rect 328604 87156 328610 87168
rect 338022 87156 338028 87168
rect 328604 87128 338028 87156
rect 328604 87116 328610 87128
rect 338022 87116 338028 87128
rect 338080 87116 338086 87168
rect 340782 87116 340788 87168
rect 340840 87156 340846 87168
rect 354582 87156 354588 87168
rect 340840 87128 354588 87156
rect 340840 87116 340846 87128
rect 354582 87116 354588 87128
rect 354640 87116 354646 87168
rect 415394 87048 415400 87100
rect 415452 87088 415458 87100
rect 424778 87088 424784 87100
rect 415452 87060 424784 87088
rect 415452 87048 415458 87060
rect 424778 87048 424784 87060
rect 424836 87048 424842 87100
rect 475930 87048 475936 87100
rect 475988 87088 475994 87100
rect 476114 87088 476120 87100
rect 475988 87060 476120 87088
rect 475988 87048 475994 87060
rect 476114 87048 476120 87060
rect 476172 87048 476178 87100
rect 572622 87048 572628 87100
rect 572680 87088 572686 87100
rect 576762 87088 576768 87100
rect 572680 87060 576768 87088
rect 572680 87048 572686 87060
rect 576762 87048 576768 87060
rect 576820 87048 576826 87100
rect 267090 87020 267096 87032
rect 267016 86992 267096 87020
rect 267016 86964 267044 86992
rect 267090 86980 267096 86992
rect 267148 86980 267154 87032
rect 331306 86980 331312 87032
rect 331364 87020 331370 87032
rect 331398 87020 331404 87032
rect 331364 86992 331404 87020
rect 331364 86980 331370 86992
rect 331398 86980 331404 86992
rect 331456 86980 331462 87032
rect 334250 86980 334256 87032
rect 334308 87020 334314 87032
rect 334434 87020 334440 87032
rect 334308 86992 334440 87020
rect 334308 86980 334314 86992
rect 334434 86980 334440 86992
rect 334492 86980 334498 87032
rect 380986 87020 380992 87032
rect 380947 86992 380992 87020
rect 380986 86980 380992 86992
rect 381044 86980 381050 87032
rect 407761 87023 407819 87029
rect 407761 86989 407773 87023
rect 407807 87020 407819 87023
rect 407850 87020 407856 87032
rect 407807 86992 407856 87020
rect 407807 86989 407819 86992
rect 407761 86983 407819 86989
rect 407850 86980 407856 86992
rect 407908 86980 407914 87032
rect 425054 86980 425060 87032
rect 425112 87020 425118 87032
rect 434530 87020 434536 87032
rect 425112 86992 434536 87020
rect 425112 86980 425118 86992
rect 434530 86980 434536 86992
rect 434588 86980 434594 87032
rect 466546 86980 466552 87032
rect 466604 87020 466610 87032
rect 466638 87020 466644 87032
rect 466604 86992 466644 87020
rect 466604 86980 466610 86992
rect 466638 86980 466644 86992
rect 466696 86980 466702 87032
rect 241790 86952 241796 86964
rect 241751 86924 241796 86952
rect 241790 86912 241796 86924
rect 241848 86912 241854 86964
rect 266998 86912 267004 86964
rect 267056 86912 267062 86964
rect 288618 86952 288624 86964
rect 288579 86924 288624 86952
rect 288618 86912 288624 86924
rect 288676 86912 288682 86964
rect 305178 86952 305184 86964
rect 305139 86924 305184 86952
rect 305178 86912 305184 86924
rect 305236 86912 305242 86964
rect 308122 86952 308128 86964
rect 308083 86924 308128 86952
rect 308122 86912 308128 86924
rect 308180 86912 308186 86964
rect 310698 86952 310704 86964
rect 310659 86924 310704 86952
rect 310698 86912 310704 86924
rect 310756 86912 310762 86964
rect 324498 86912 324504 86964
rect 324556 86952 324562 86964
rect 324590 86952 324596 86964
rect 324556 86924 324596 86952
rect 324556 86912 324562 86924
rect 324590 86912 324596 86924
rect 324648 86912 324654 86964
rect 342530 86952 342536 86964
rect 342491 86924 342536 86952
rect 342530 86912 342536 86924
rect 342588 86912 342594 86964
rect 346578 86952 346584 86964
rect 346539 86924 346584 86952
rect 346578 86912 346584 86924
rect 346636 86912 346642 86964
rect 382458 86952 382464 86964
rect 382419 86924 382464 86952
rect 382458 86912 382464 86924
rect 382516 86912 382522 86964
rect 422386 86952 422392 86964
rect 422347 86924 422392 86952
rect 422386 86912 422392 86924
rect 422444 86912 422450 86964
rect 270586 86844 270592 86896
rect 270644 86884 270650 86896
rect 270862 86884 270868 86896
rect 270644 86856 270868 86884
rect 270644 86844 270650 86856
rect 270862 86844 270868 86856
rect 270920 86844 270926 86896
rect 357526 86844 357532 86896
rect 357584 86884 357590 86896
rect 357710 86884 357716 86896
rect 357584 86856 357716 86884
rect 357584 86844 357590 86856
rect 357710 86844 357716 86856
rect 357768 86844 357774 86896
rect 240137 85663 240195 85669
rect 240137 85629 240149 85663
rect 240183 85660 240195 85663
rect 240226 85660 240232 85672
rect 240183 85632 240232 85660
rect 240183 85629 240195 85632
rect 240137 85623 240195 85629
rect 240226 85620 240232 85632
rect 240284 85620 240290 85672
rect 287146 85660 287152 85672
rect 287107 85632 287152 85660
rect 287146 85620 287152 85632
rect 287204 85620 287210 85672
rect 236270 85592 236276 85604
rect 236231 85564 236276 85592
rect 236270 85552 236276 85564
rect 236328 85552 236334 85604
rect 295518 85552 295524 85604
rect 295576 85592 295582 85604
rect 295610 85592 295616 85604
rect 295576 85564 295616 85592
rect 295576 85552 295582 85564
rect 295610 85552 295616 85564
rect 295668 85552 295674 85604
rect 327166 85552 327172 85604
rect 327224 85592 327230 85604
rect 327258 85592 327264 85604
rect 327224 85564 327264 85592
rect 327224 85552 327230 85564
rect 327258 85552 327264 85564
rect 327316 85552 327322 85604
rect 347866 85552 347872 85604
rect 347924 85592 347930 85604
rect 348050 85592 348056 85604
rect 347924 85564 348056 85592
rect 347924 85552 347930 85564
rect 348050 85552 348056 85564
rect 348108 85552 348114 85604
rect 352098 85552 352104 85604
rect 352156 85592 352162 85604
rect 352190 85592 352196 85604
rect 352156 85564 352196 85592
rect 352156 85552 352162 85564
rect 352190 85552 352196 85564
rect 352248 85552 352254 85604
rect 375561 85595 375619 85601
rect 375561 85561 375573 85595
rect 375607 85592 375619 85595
rect 375650 85592 375656 85604
rect 375607 85564 375656 85592
rect 375607 85561 375619 85564
rect 375561 85555 375619 85561
rect 375650 85552 375656 85564
rect 375708 85552 375714 85604
rect 249978 85524 249984 85536
rect 249939 85496 249984 85524
rect 249978 85484 249984 85496
rect 250036 85484 250042 85536
rect 254121 85527 254179 85533
rect 254121 85493 254133 85527
rect 254167 85524 254179 85527
rect 254210 85524 254216 85536
rect 254167 85496 254216 85524
rect 254167 85493 254179 85496
rect 254121 85487 254179 85493
rect 254210 85484 254216 85496
rect 254268 85484 254274 85536
rect 287146 85484 287152 85536
rect 287204 85524 287210 85536
rect 287241 85527 287299 85533
rect 287241 85524 287253 85527
rect 287204 85496 287253 85524
rect 287204 85484 287210 85496
rect 287241 85493 287253 85496
rect 287287 85493 287299 85527
rect 334250 85524 334256 85536
rect 334211 85496 334256 85524
rect 287241 85487 287299 85493
rect 334250 85484 334256 85496
rect 334308 85484 334314 85536
rect 380986 85524 380992 85536
rect 380947 85496 380992 85524
rect 380986 85484 380992 85496
rect 381044 85484 381050 85536
rect 407758 85524 407764 85536
rect 407719 85496 407764 85524
rect 407758 85484 407764 85496
rect 407816 85484 407822 85536
rect 408681 85527 408739 85533
rect 408681 85493 408693 85527
rect 408727 85524 408739 85527
rect 408862 85524 408868 85536
rect 408727 85496 408868 85524
rect 408727 85493 408739 85496
rect 408681 85487 408739 85493
rect 408862 85484 408868 85496
rect 408920 85484 408926 85536
rect 466454 85524 466460 85536
rect 466415 85496 466460 85524
rect 466454 85484 466460 85496
rect 466512 85484 466518 85536
rect 472066 85524 472072 85536
rect 472027 85496 472072 85524
rect 472066 85484 472072 85496
rect 472124 85484 472130 85536
rect 480438 85524 480444 85536
rect 480399 85496 480444 85524
rect 480438 85484 480444 85496
rect 480496 85484 480502 85536
rect 236270 85456 236276 85468
rect 236231 85428 236276 85456
rect 236270 85416 236276 85428
rect 236328 85416 236334 85468
rect 272058 84300 272064 84312
rect 271984 84272 272064 84300
rect 271984 84244 272012 84272
rect 272058 84260 272064 84272
rect 272116 84260 272122 84312
rect 271966 84192 271972 84244
rect 272024 84192 272030 84244
rect 294138 84232 294144 84244
rect 294099 84204 294144 84232
rect 294138 84192 294144 84204
rect 294196 84192 294202 84244
rect 298554 84192 298560 84244
rect 298612 84232 298618 84244
rect 364518 84232 364524 84244
rect 298612 84204 298657 84232
rect 364479 84204 364524 84232
rect 298612 84192 298618 84204
rect 364518 84192 364524 84204
rect 364576 84192 364582 84244
rect 259641 84167 259699 84173
rect 259641 84133 259653 84167
rect 259687 84164 259699 84167
rect 259730 84164 259736 84176
rect 259687 84136 259736 84164
rect 259687 84133 259699 84136
rect 259641 84127 259699 84133
rect 259730 84124 259736 84136
rect 259788 84124 259794 84176
rect 353478 84124 353484 84176
rect 353536 84124 353542 84176
rect 356514 84124 356520 84176
rect 356572 84124 356578 84176
rect 357710 84164 357716 84176
rect 357671 84136 357716 84164
rect 357710 84124 357716 84136
rect 357768 84124 357774 84176
rect 358998 84164 359004 84176
rect 358959 84136 359004 84164
rect 358998 84124 359004 84136
rect 359056 84124 359062 84176
rect 353386 84056 353392 84108
rect 353444 84096 353450 84108
rect 353496 84096 353524 84124
rect 353444 84068 353524 84096
rect 353444 84056 353450 84068
rect 356532 84040 356560 84124
rect 356514 83988 356520 84040
rect 356572 83988 356578 84040
rect 271966 82804 271972 82816
rect 271927 82776 271972 82804
rect 271966 82764 271972 82776
rect 272024 82764 272030 82816
rect 356425 82807 356483 82813
rect 356425 82773 356437 82807
rect 356471 82804 356483 82807
rect 356514 82804 356520 82816
rect 356471 82776 356520 82804
rect 356471 82773 356483 82776
rect 356425 82767 356483 82773
rect 356514 82764 356520 82776
rect 356572 82764 356578 82816
rect 243173 80767 243231 80773
rect 243173 80733 243185 80767
rect 243219 80764 243231 80767
rect 243354 80764 243360 80776
rect 243219 80736 243360 80764
rect 243219 80733 243231 80736
rect 243173 80727 243231 80733
rect 243354 80724 243360 80736
rect 243412 80724 243418 80776
rect 433613 80223 433671 80229
rect 433613 80189 433625 80223
rect 433659 80220 433671 80223
rect 433702 80220 433708 80232
rect 433659 80192 433708 80220
rect 433659 80189 433671 80192
rect 433613 80183 433671 80189
rect 433702 80180 433708 80192
rect 433760 80180 433766 80232
rect 309318 80084 309324 80096
rect 309279 80056 309324 80084
rect 309318 80044 309324 80056
rect 309376 80044 309382 80096
rect 332778 80044 332784 80096
rect 332836 80044 332842 80096
rect 336826 80044 336832 80096
rect 336884 80044 336890 80096
rect 365898 80044 365904 80096
rect 365956 80044 365962 80096
rect 376938 80044 376944 80096
rect 376996 80044 377002 80096
rect 387978 80044 387984 80096
rect 388036 80044 388042 80096
rect 255498 80016 255504 80028
rect 255459 79988 255504 80016
rect 255498 79976 255504 79988
rect 255556 79976 255562 80028
rect 332796 79960 332824 80044
rect 336844 79960 336872 80044
rect 342530 80016 342536 80028
rect 342491 79988 342536 80016
rect 342530 79976 342536 79988
rect 342588 79976 342594 80028
rect 346578 80016 346584 80028
rect 346539 79988 346584 80016
rect 346578 79976 346584 79988
rect 346636 79976 346642 80028
rect 365916 79960 365944 80044
rect 376956 79960 376984 80044
rect 387996 79960 388024 80044
rect 332778 79908 332784 79960
rect 332836 79908 332842 79960
rect 336826 79908 336832 79960
rect 336884 79908 336890 79960
rect 365898 79908 365904 79960
rect 365956 79908 365962 79960
rect 376938 79908 376944 79960
rect 376996 79908 377002 79960
rect 387978 79908 387984 79960
rect 388036 79908 388042 79960
rect 249978 79336 249984 79348
rect 249939 79308 249984 79336
rect 249978 79296 249984 79308
rect 250036 79296 250042 79348
rect 334253 79339 334311 79345
rect 334253 79305 334265 79339
rect 334299 79336 334311 79339
rect 334434 79336 334440 79348
rect 334299 79308 334440 79336
rect 334299 79305 334311 79308
rect 334253 79299 334311 79305
rect 334434 79296 334440 79308
rect 334492 79296 334498 79348
rect 3326 79160 3332 79212
rect 3384 79200 3390 79212
rect 7650 79200 7656 79212
rect 3384 79172 7656 79200
rect 3384 79160 3390 79172
rect 7650 79160 7656 79172
rect 7708 79160 7714 79212
rect 266449 77979 266507 77985
rect 266449 77945 266461 77979
rect 266495 77976 266507 77979
rect 266630 77976 266636 77988
rect 266495 77948 266636 77976
rect 266495 77945 266507 77948
rect 266449 77939 266507 77945
rect 266630 77936 266636 77948
rect 266688 77936 266694 77988
rect 359001 77979 359059 77985
rect 359001 77945 359013 77979
rect 359047 77976 359059 77979
rect 359274 77976 359280 77988
rect 359047 77948 359280 77976
rect 359047 77945 359059 77948
rect 359001 77939 359059 77945
rect 359274 77936 359280 77948
rect 359332 77936 359338 77988
rect 386598 77392 386604 77444
rect 386656 77392 386662 77444
rect 348050 77364 348056 77376
rect 347976 77336 348056 77364
rect 347976 77308 348004 77336
rect 348050 77324 348056 77336
rect 348108 77324 348114 77376
rect 352009 77367 352067 77373
rect 352009 77333 352021 77367
rect 352055 77364 352067 77367
rect 352098 77364 352104 77376
rect 352055 77336 352104 77364
rect 352055 77333 352067 77336
rect 352009 77327 352067 77333
rect 352098 77324 352104 77336
rect 352156 77324 352162 77376
rect 386616 77308 386644 77392
rect 392210 77364 392216 77376
rect 392136 77336 392216 77364
rect 392136 77308 392164 77336
rect 392210 77324 392216 77336
rect 392268 77324 392274 77376
rect 416866 77324 416872 77376
rect 416924 77364 416930 77376
rect 416958 77364 416964 77376
rect 416924 77336 416964 77364
rect 416924 77324 416930 77336
rect 416958 77324 416964 77336
rect 417016 77324 417022 77376
rect 232038 77256 232044 77308
rect 232096 77256 232102 77308
rect 241790 77296 241796 77308
rect 241751 77268 241796 77296
rect 241790 77256 241796 77268
rect 241848 77256 241854 77308
rect 270678 77256 270684 77308
rect 270736 77296 270742 77308
rect 270862 77296 270868 77308
rect 270736 77268 270868 77296
rect 270736 77256 270742 77268
rect 270862 77256 270868 77268
rect 270920 77256 270926 77308
rect 281718 77296 281724 77308
rect 281679 77268 281724 77296
rect 281718 77256 281724 77268
rect 281776 77256 281782 77308
rect 288618 77296 288624 77308
rect 288579 77268 288624 77296
rect 288618 77256 288624 77268
rect 288676 77256 288682 77308
rect 305178 77296 305184 77308
rect 305139 77268 305184 77296
rect 305178 77256 305184 77268
rect 305236 77256 305242 77308
rect 308122 77296 308128 77308
rect 308083 77268 308128 77296
rect 308122 77256 308128 77268
rect 308180 77256 308186 77308
rect 309226 77256 309232 77308
rect 309284 77296 309290 77308
rect 309321 77299 309379 77305
rect 309321 77296 309333 77299
rect 309284 77268 309333 77296
rect 309284 77256 309290 77268
rect 309321 77265 309333 77268
rect 309367 77265 309379 77299
rect 310698 77296 310704 77308
rect 310659 77268 310704 77296
rect 309321 77259 309379 77265
rect 310698 77256 310704 77268
rect 310756 77256 310762 77308
rect 347958 77256 347964 77308
rect 348016 77256 348022 77308
rect 386598 77256 386604 77308
rect 386656 77256 386662 77308
rect 392118 77256 392124 77308
rect 392176 77256 392182 77308
rect 422389 77299 422447 77305
rect 422389 77265 422401 77299
rect 422435 77296 422447 77299
rect 422478 77296 422484 77308
rect 422435 77268 422484 77296
rect 422435 77265 422447 77268
rect 422389 77259 422447 77265
rect 422478 77256 422484 77268
rect 422536 77256 422542 77308
rect 433610 77296 433616 77308
rect 433571 77268 433616 77296
rect 433610 77256 433616 77268
rect 433668 77256 433674 77308
rect 232056 77172 232084 77256
rect 232038 77120 232044 77172
rect 232096 77120 232102 77172
rect 466457 77163 466515 77169
rect 466457 77129 466469 77163
rect 466503 77160 466515 77163
rect 466546 77160 466552 77172
rect 466503 77132 466552 77160
rect 466503 77129 466515 77132
rect 466457 77123 466515 77129
rect 466546 77120 466552 77132
rect 466604 77120 466610 77172
rect 480441 77163 480499 77169
rect 480441 77129 480453 77163
rect 480487 77160 480499 77163
rect 480530 77160 480536 77172
rect 480487 77132 480536 77160
rect 480487 77129 480499 77132
rect 480441 77123 480499 77129
rect 480530 77120 480536 77132
rect 480588 77120 480594 77172
rect 427906 76344 427912 76356
rect 427867 76316 427912 76344
rect 427906 76304 427912 76316
rect 427964 76304 427970 76356
rect 398742 76236 398748 76288
rect 398800 76276 398806 76288
rect 405642 76276 405648 76288
rect 398800 76248 405648 76276
rect 398800 76236 398806 76248
rect 405642 76236 405648 76248
rect 405700 76236 405706 76288
rect 309042 76168 309048 76220
rect 309100 76208 309106 76220
rect 317322 76208 317328 76220
rect 309100 76180 317328 76208
rect 309100 76168 309106 76180
rect 317322 76168 317328 76180
rect 317380 76168 317386 76220
rect 514570 76100 514576 76152
rect 514628 76140 514634 76152
rect 516870 76140 516876 76152
rect 514628 76112 516876 76140
rect 514628 76100 514634 76112
rect 516870 76100 516876 76112
rect 516928 76100 516934 76152
rect 475930 76032 475936 76084
rect 475988 76072 475994 76084
rect 478138 76072 478144 76084
rect 475988 76044 478144 76072
rect 475988 76032 475994 76044
rect 478138 76032 478144 76044
rect 478196 76032 478202 76084
rect 283466 75964 283472 76016
rect 283524 76004 283530 76016
rect 290550 76004 290556 76016
rect 283524 75976 290556 76004
rect 283524 75964 283530 75976
rect 290550 75964 290556 75976
rect 290608 75964 290614 76016
rect 346210 75964 346216 76016
rect 346268 76004 346274 76016
rect 346268 75976 346348 76004
rect 346268 75964 346274 75976
rect 346320 75948 346348 75976
rect 370038 75964 370044 76016
rect 370096 76004 370102 76016
rect 370314 76004 370320 76016
rect 370096 75976 370320 76004
rect 370096 75964 370102 75976
rect 370314 75964 370320 75976
rect 370372 75964 370378 76016
rect 408678 76004 408684 76016
rect 408639 75976 408684 76004
rect 408678 75964 408684 75976
rect 408736 75964 408742 76016
rect 524230 75964 524236 76016
rect 524288 76004 524294 76016
rect 526438 76004 526444 76016
rect 524288 75976 526444 76004
rect 524288 75964 524294 75976
rect 526438 75964 526444 75976
rect 526496 75964 526502 76016
rect 236273 75939 236331 75945
rect 236273 75905 236285 75939
rect 236319 75936 236331 75939
rect 236362 75936 236368 75948
rect 236319 75908 236368 75936
rect 236319 75905 236331 75908
rect 236273 75899 236331 75905
rect 236362 75896 236368 75908
rect 236420 75896 236426 75948
rect 240226 75896 240232 75948
rect 240284 75936 240290 75948
rect 240410 75936 240416 75948
rect 240284 75908 240416 75936
rect 240284 75896 240290 75908
rect 240410 75896 240416 75908
rect 240468 75896 240474 75948
rect 281718 75936 281724 75948
rect 281679 75908 281724 75936
rect 281718 75896 281724 75908
rect 281776 75896 281782 75948
rect 287238 75936 287244 75948
rect 287199 75908 287244 75936
rect 287238 75896 287244 75908
rect 287296 75896 287302 75948
rect 319070 75896 319076 75948
rect 319128 75936 319134 75948
rect 319162 75936 319168 75948
rect 319128 75908 319168 75936
rect 319128 75896 319134 75908
rect 319162 75896 319168 75908
rect 319220 75896 319226 75948
rect 327166 75896 327172 75948
rect 327224 75936 327230 75948
rect 327258 75936 327264 75948
rect 327224 75908 327264 75936
rect 327224 75896 327230 75908
rect 327258 75896 327264 75908
rect 327316 75896 327322 75948
rect 346302 75896 346308 75948
rect 346360 75896 346366 75948
rect 380989 75939 381047 75945
rect 380989 75905 381001 75939
rect 381035 75936 381047 75939
rect 381078 75936 381084 75948
rect 381035 75908 381084 75936
rect 381035 75905 381047 75908
rect 380989 75899 381047 75905
rect 381078 75896 381084 75908
rect 381136 75896 381142 75948
rect 382458 75936 382464 75948
rect 382419 75908 382464 75936
rect 382458 75896 382464 75908
rect 382516 75896 382522 75948
rect 407758 75936 407764 75948
rect 407719 75908 407764 75936
rect 407758 75896 407764 75908
rect 407816 75896 407822 75948
rect 270678 75868 270684 75880
rect 270639 75840 270684 75868
rect 270678 75828 270684 75840
rect 270736 75828 270742 75880
rect 375558 75868 375564 75880
rect 375519 75840 375564 75868
rect 375558 75828 375564 75840
rect 375616 75828 375622 75880
rect 408678 75868 408684 75880
rect 408639 75840 408684 75868
rect 408678 75828 408684 75840
rect 408736 75828 408742 75880
rect 266998 74604 267004 74656
rect 267056 74644 267062 74656
rect 267056 74616 267228 74644
rect 267056 74604 267062 74616
rect 255498 74576 255504 74588
rect 255459 74548 255504 74576
rect 255498 74536 255504 74548
rect 255556 74536 255562 74588
rect 266814 74468 266820 74520
rect 266872 74508 266878 74520
rect 267200 74508 267228 74616
rect 357710 74576 357716 74588
rect 357671 74548 357716 74576
rect 357710 74536 357716 74548
rect 357768 74536 357774 74588
rect 266872 74480 267228 74508
rect 334345 74511 334403 74517
rect 266872 74468 266878 74480
rect 334345 74477 334357 74511
rect 334391 74508 334403 74511
rect 334434 74508 334440 74520
rect 334391 74480 334440 74508
rect 334391 74477 334403 74480
rect 334345 74471 334403 74477
rect 334434 74468 334440 74480
rect 334492 74468 334498 74520
rect 364518 74508 364524 74520
rect 364479 74480 364524 74508
rect 364518 74468 364524 74480
rect 364576 74468 364582 74520
rect 271966 73216 271972 73228
rect 271927 73188 271972 73216
rect 271966 73176 271972 73188
rect 272024 73176 272030 73228
rect 356422 73216 356428 73228
rect 356383 73188 356428 73216
rect 356422 73176 356428 73188
rect 356480 73176 356486 73228
rect 359182 73108 359188 73160
rect 359240 73148 359246 73160
rect 359274 73148 359280 73160
rect 359240 73120 359280 73148
rect 359240 73108 359246 73120
rect 359274 73108 359280 73120
rect 359332 73108 359338 73160
rect 294046 72428 294052 72480
rect 294104 72468 294110 72480
rect 294230 72468 294236 72480
rect 294104 72440 294236 72468
rect 294104 72428 294110 72440
rect 294230 72428 294236 72440
rect 294288 72428 294294 72480
rect 259638 71108 259644 71120
rect 259599 71080 259644 71108
rect 259638 71068 259644 71080
rect 259696 71068 259702 71120
rect 244458 70496 244464 70508
rect 244419 70468 244464 70496
rect 244458 70456 244464 70468
rect 244516 70456 244522 70508
rect 277578 70456 277584 70508
rect 277636 70456 277642 70508
rect 305178 70496 305184 70508
rect 305139 70468 305184 70496
rect 305178 70456 305184 70468
rect 305236 70456 305242 70508
rect 416958 70496 416964 70508
rect 416884 70468 416964 70496
rect 277596 70372 277624 70456
rect 416884 70372 416912 70468
rect 416958 70456 416964 70468
rect 417016 70456 417022 70508
rect 277578 70320 277584 70372
rect 277636 70320 277642 70372
rect 416866 70320 416872 70372
rect 416924 70320 416930 70372
rect 236362 67844 236368 67856
rect 236288 67816 236368 67844
rect 236288 67584 236316 67816
rect 236362 67804 236368 67816
rect 236420 67804 236426 67856
rect 331398 67736 331404 67788
rect 331456 67736 331462 67788
rect 309226 67668 309232 67720
rect 309284 67668 309290 67720
rect 240134 67600 240140 67652
rect 240192 67640 240198 67652
rect 240318 67640 240324 67652
rect 240192 67612 240324 67640
rect 240192 67600 240198 67612
rect 240318 67600 240324 67612
rect 240376 67600 240382 67652
rect 243170 67640 243176 67652
rect 243131 67612 243176 67640
rect 243170 67600 243176 67612
rect 243228 67600 243234 67652
rect 244458 67640 244464 67652
rect 244419 67612 244464 67640
rect 244458 67600 244464 67612
rect 244516 67600 244522 67652
rect 254118 67640 254124 67652
rect 254079 67612 254124 67640
rect 254118 67600 254124 67612
rect 254176 67600 254182 67652
rect 292758 67600 292764 67652
rect 292816 67640 292822 67652
rect 292850 67640 292856 67652
rect 292816 67612 292856 67640
rect 292816 67600 292822 67612
rect 292850 67600 292856 67612
rect 292908 67600 292914 67652
rect 305178 67640 305184 67652
rect 305139 67612 305184 67640
rect 305178 67600 305184 67612
rect 305236 67600 305242 67652
rect 309244 67640 309272 67668
rect 331416 67652 331444 67736
rect 376938 67708 376944 67720
rect 376864 67680 376944 67708
rect 376864 67652 376892 67680
rect 376938 67668 376944 67680
rect 376996 67668 377002 67720
rect 309318 67640 309324 67652
rect 309244 67612 309324 67640
rect 309318 67600 309324 67612
rect 309376 67600 309382 67652
rect 310606 67600 310612 67652
rect 310664 67640 310670 67652
rect 310698 67640 310704 67652
rect 310664 67612 310704 67640
rect 310664 67600 310670 67612
rect 310698 67600 310704 67612
rect 310756 67600 310762 67652
rect 318978 67600 318984 67652
rect 319036 67640 319042 67652
rect 319070 67640 319076 67652
rect 319036 67612 319076 67640
rect 319036 67600 319042 67612
rect 319070 67600 319076 67612
rect 319128 67600 319134 67652
rect 331398 67600 331404 67652
rect 331456 67600 331462 67652
rect 376846 67600 376852 67652
rect 376904 67600 376910 67652
rect 400490 67600 400496 67652
rect 400548 67640 400554 67652
rect 400582 67640 400588 67652
rect 400548 67612 400588 67640
rect 400548 67600 400554 67612
rect 400582 67600 400588 67612
rect 400640 67600 400646 67652
rect 422386 67600 422392 67652
rect 422444 67640 422450 67652
rect 422478 67640 422484 67652
rect 422444 67612 422484 67640
rect 422444 67600 422450 67612
rect 422478 67600 422484 67612
rect 422536 67600 422542 67652
rect 427909 67643 427967 67649
rect 427909 67609 427921 67643
rect 427955 67640 427967 67643
rect 427998 67640 428004 67652
rect 427955 67612 428004 67640
rect 427955 67609 427967 67612
rect 427909 67603 427967 67609
rect 427998 67600 428004 67612
rect 428056 67600 428062 67652
rect 472066 67640 472072 67652
rect 472027 67612 472072 67640
rect 472066 67600 472072 67612
rect 472124 67600 472130 67652
rect 231854 67532 231860 67584
rect 231912 67572 231918 67584
rect 232038 67572 232044 67584
rect 231912 67544 232044 67572
rect 231912 67532 231918 67544
rect 232038 67532 232044 67544
rect 232096 67532 232102 67584
rect 236270 67532 236276 67584
rect 236328 67532 236334 67584
rect 281718 67572 281724 67584
rect 281679 67544 281724 67572
rect 281718 67532 281724 67544
rect 281776 67532 281782 67584
rect 381078 67572 381084 67584
rect 381039 67544 381084 67572
rect 381078 67532 381084 67544
rect 381136 67532 381142 67584
rect 416866 67532 416872 67584
rect 416924 67572 416930 67584
rect 417050 67572 417056 67584
rect 416924 67544 417056 67572
rect 416924 67532 416930 67544
rect 417050 67532 417056 67544
rect 417108 67532 417114 67584
rect 480254 67532 480260 67584
rect 480312 67572 480318 67584
rect 480438 67572 480444 67584
rect 480312 67544 480444 67572
rect 480312 67532 480318 67544
rect 480438 67532 480444 67544
rect 480496 67532 480502 67584
rect 370038 66376 370044 66428
rect 370096 66376 370102 66428
rect 283190 66348 283196 66360
rect 283116 66320 283196 66348
rect 265158 66240 265164 66292
rect 265216 66280 265222 66292
rect 265250 66280 265256 66292
rect 265216 66252 265256 66280
rect 265216 66240 265222 66252
rect 265250 66240 265256 66252
rect 265308 66240 265314 66292
rect 270681 66283 270739 66289
rect 270681 66249 270693 66283
rect 270727 66280 270739 66283
rect 270770 66280 270776 66292
rect 270727 66252 270776 66280
rect 270727 66249 270739 66252
rect 270681 66243 270739 66249
rect 270770 66240 270776 66252
rect 270828 66240 270834 66292
rect 249886 66172 249892 66224
rect 249944 66212 249950 66224
rect 249978 66212 249984 66224
rect 249944 66184 249984 66212
rect 249944 66172 249950 66184
rect 249978 66172 249984 66184
rect 250036 66172 250042 66224
rect 283116 66221 283144 66320
rect 283190 66308 283196 66320
rect 283248 66308 283254 66360
rect 287238 66308 287244 66360
rect 287296 66308 287302 66360
rect 287256 66221 287284 66308
rect 370056 66292 370084 66376
rect 375561 66351 375619 66357
rect 375561 66348 375573 66351
rect 375484 66320 375573 66348
rect 352006 66280 352012 66292
rect 351967 66252 352012 66280
rect 352006 66240 352012 66252
rect 352064 66240 352070 66292
rect 370038 66240 370044 66292
rect 370096 66240 370102 66292
rect 283101 66215 283159 66221
rect 283101 66181 283113 66215
rect 283147 66181 283159 66215
rect 283101 66175 283159 66181
rect 287241 66215 287299 66221
rect 287241 66181 287253 66215
rect 287287 66181 287299 66215
rect 292758 66212 292764 66224
rect 292719 66184 292764 66212
rect 287241 66175 287299 66181
rect 292758 66172 292764 66184
rect 292816 66172 292822 66224
rect 293954 66172 293960 66224
rect 294012 66212 294018 66224
rect 294230 66212 294236 66224
rect 294012 66184 294236 66212
rect 294012 66172 294018 66184
rect 294230 66172 294236 66184
rect 294288 66172 294294 66224
rect 324498 66212 324504 66224
rect 324459 66184 324504 66212
rect 324498 66172 324504 66184
rect 324556 66172 324562 66224
rect 346578 66172 346584 66224
rect 346636 66212 346642 66224
rect 346670 66212 346676 66224
rect 346636 66184 346676 66212
rect 346636 66172 346642 66184
rect 346670 66172 346676 66184
rect 346728 66172 346734 66224
rect 375484 66221 375512 66320
rect 375561 66317 375573 66320
rect 375607 66317 375619 66351
rect 375561 66311 375619 66317
rect 408681 66283 408739 66289
rect 408681 66249 408693 66283
rect 408727 66280 408739 66283
rect 408770 66280 408776 66292
rect 408727 66252 408776 66280
rect 408727 66249 408739 66252
rect 408681 66243 408739 66249
rect 408770 66240 408776 66252
rect 408828 66240 408834 66292
rect 375469 66215 375527 66221
rect 375469 66181 375481 66215
rect 375515 66181 375527 66215
rect 393222 66212 393228 66224
rect 375469 66175 375527 66181
rect 393148 66184 393228 66212
rect 393148 66156 393176 66184
rect 393222 66172 393228 66184
rect 393280 66172 393286 66224
rect 407758 66212 407764 66224
rect 407719 66184 407764 66212
rect 407758 66172 407764 66184
rect 407816 66172 407822 66224
rect 393130 66104 393136 66156
rect 393188 66104 393194 66156
rect 334342 64988 334348 65000
rect 334303 64960 334348 64988
rect 334342 64948 334348 64960
rect 334400 64948 334406 65000
rect 266446 64920 266452 64932
rect 266407 64892 266452 64920
rect 266446 64880 266452 64892
rect 266504 64880 266510 64932
rect 357618 64880 357624 64932
rect 357676 64920 357682 64932
rect 357710 64920 357716 64932
rect 357676 64892 357716 64920
rect 357676 64880 357682 64892
rect 357710 64880 357716 64892
rect 357768 64880 357774 64932
rect 364518 64920 364524 64932
rect 364479 64892 364524 64920
rect 364518 64880 364524 64892
rect 364576 64880 364582 64932
rect 249886 64852 249892 64864
rect 249847 64824 249892 64852
rect 249886 64812 249892 64824
rect 249944 64812 249950 64864
rect 255498 64852 255504 64864
rect 255459 64824 255504 64852
rect 255498 64812 255504 64824
rect 255556 64812 255562 64864
rect 271966 64812 271972 64864
rect 272024 64852 272030 64864
rect 272058 64852 272064 64864
rect 272024 64824 272064 64852
rect 272024 64812 272030 64824
rect 272058 64812 272064 64824
rect 272116 64812 272122 64864
rect 310606 64852 310612 64864
rect 310567 64824 310612 64852
rect 310606 64812 310612 64824
rect 310664 64812 310670 64864
rect 331398 64852 331404 64864
rect 331359 64824 331404 64852
rect 331398 64812 331404 64824
rect 331456 64812 331462 64864
rect 334342 64852 334348 64864
rect 334303 64824 334348 64852
rect 334342 64812 334348 64824
rect 334400 64812 334406 64864
rect 356422 64812 356428 64864
rect 356480 64852 356486 64864
rect 356606 64852 356612 64864
rect 356480 64824 356612 64852
rect 356480 64812 356486 64824
rect 356606 64812 356612 64824
rect 356664 64812 356670 64864
rect 240042 64472 240048 64524
rect 240100 64512 240106 64524
rect 248322 64512 248328 64524
rect 240100 64484 248328 64512
rect 240100 64472 240106 64484
rect 248322 64472 248328 64484
rect 248380 64472 248386 64524
rect 267642 63860 267648 63912
rect 267700 63900 267706 63912
rect 275922 63900 275928 63912
rect 267700 63872 275928 63900
rect 267700 63860 267706 63872
rect 275922 63860 275928 63872
rect 275980 63860 275986 63912
rect 355502 63792 355508 63844
rect 355560 63832 355566 63844
rect 360378 63832 360384 63844
rect 355560 63804 360384 63832
rect 355560 63792 355566 63804
rect 360378 63792 360384 63804
rect 360436 63792 360442 63844
rect 393314 63792 393320 63844
rect 393372 63832 393378 63844
rect 405642 63832 405648 63844
rect 393372 63804 405648 63832
rect 393372 63792 393378 63804
rect 405642 63792 405648 63804
rect 405700 63792 405706 63844
rect 346210 63588 346216 63640
rect 346268 63628 346274 63640
rect 346486 63628 346492 63640
rect 346268 63600 346492 63628
rect 346268 63588 346274 63600
rect 346486 63588 346492 63600
rect 346544 63588 346550 63640
rect 521654 63588 521660 63640
rect 521712 63628 521718 63640
rect 526438 63628 526444 63640
rect 521712 63600 526444 63628
rect 521712 63588 521718 63600
rect 526438 63588 526444 63600
rect 526496 63588 526502 63640
rect 337470 63520 337476 63572
rect 337528 63560 337534 63572
rect 344922 63560 344928 63572
rect 337528 63532 344928 63560
rect 337528 63520 337534 63532
rect 344922 63520 344928 63532
rect 344980 63520 344986 63572
rect 356517 63495 356575 63501
rect 356517 63461 356529 63495
rect 356563 63492 356575 63495
rect 356606 63492 356612 63504
rect 356563 63464 356612 63492
rect 356563 63461 356575 63464
rect 356517 63455 356575 63461
rect 356606 63452 356612 63464
rect 356664 63452 356670 63504
rect 359182 63492 359188 63504
rect 359143 63464 359188 63492
rect 359182 63452 359188 63464
rect 359240 63452 359246 63504
rect 281718 61452 281724 61464
rect 281679 61424 281724 61452
rect 281718 61412 281724 61424
rect 281776 61412 281782 61464
rect 386598 61412 386604 61464
rect 386656 61452 386662 61464
rect 386782 61452 386788 61464
rect 386656 61424 386788 61452
rect 386656 61412 386662 61424
rect 386782 61412 386788 61424
rect 386840 61412 386846 61464
rect 259638 60800 259644 60852
rect 259696 60800 259702 60852
rect 270770 60840 270776 60852
rect 270696 60812 270776 60840
rect 259656 60716 259684 60800
rect 270696 60716 270724 60812
rect 270770 60800 270776 60812
rect 270828 60800 270834 60852
rect 347958 60800 347964 60852
rect 348016 60800 348022 60852
rect 347976 60716 348004 60800
rect 259638 60664 259644 60716
rect 259696 60664 259702 60716
rect 270678 60664 270684 60716
rect 270736 60664 270742 60716
rect 347958 60664 347964 60716
rect 348016 60664 348022 60716
rect 433518 60664 433524 60716
rect 433576 60704 433582 60716
rect 433702 60704 433708 60716
rect 433576 60676 433708 60704
rect 433576 60664 433582 60676
rect 433702 60664 433708 60676
rect 433760 60664 433766 60716
rect 471974 60664 471980 60716
rect 472032 60704 472038 60716
rect 472158 60704 472164 60716
rect 472032 60676 472164 60704
rect 472032 60664 472038 60676
rect 472158 60664 472164 60676
rect 472216 60664 472222 60716
rect 240134 57944 240140 57996
rect 240192 57984 240198 57996
rect 240226 57984 240232 57996
rect 240192 57956 240232 57984
rect 240192 57944 240198 57956
rect 240226 57944 240232 57956
rect 240284 57944 240290 57996
rect 244366 57944 244372 57996
rect 244424 57984 244430 57996
rect 244550 57984 244556 57996
rect 244424 57956 244556 57984
rect 244424 57944 244430 57956
rect 244550 57944 244556 57956
rect 244608 57944 244614 57996
rect 298278 57944 298284 57996
rect 298336 57944 298342 57996
rect 308030 57944 308036 57996
rect 308088 57984 308094 57996
rect 308122 57984 308128 57996
rect 308088 57956 308128 57984
rect 308088 57944 308094 57956
rect 308122 57944 308128 57956
rect 308180 57944 308186 57996
rect 381078 57984 381084 57996
rect 381039 57956 381084 57984
rect 381078 57944 381084 57956
rect 381136 57944 381142 57996
rect 298296 57848 298324 57944
rect 387886 57876 387892 57928
rect 387944 57916 387950 57928
rect 387978 57916 387984 57928
rect 387944 57888 387984 57916
rect 387944 57876 387950 57888
rect 387978 57876 387984 57888
rect 388036 57876 388042 57928
rect 416869 57919 416927 57925
rect 416869 57885 416881 57919
rect 416915 57916 416927 57919
rect 416958 57916 416964 57928
rect 416915 57888 416964 57916
rect 416915 57885 416927 57888
rect 416869 57879 416927 57885
rect 416958 57876 416964 57888
rect 417016 57876 417022 57928
rect 433613 57919 433671 57925
rect 433613 57885 433625 57919
rect 433659 57916 433671 57919
rect 433702 57916 433708 57928
rect 433659 57888 433708 57916
rect 433659 57885 433671 57888
rect 433613 57879 433671 57885
rect 433702 57876 433708 57888
rect 433760 57876 433766 57928
rect 466549 57919 466607 57925
rect 466549 57885 466561 57919
rect 466595 57916 466607 57919
rect 466638 57916 466644 57928
rect 466595 57888 466644 57916
rect 466595 57885 466607 57888
rect 466549 57879 466607 57885
rect 466638 57876 466644 57888
rect 466696 57876 466702 57928
rect 472069 57919 472127 57925
rect 472069 57885 472081 57919
rect 472115 57916 472127 57919
rect 472158 57916 472164 57928
rect 472115 57888 472164 57916
rect 472115 57885 472127 57888
rect 472069 57879 472127 57885
rect 472158 57876 472164 57888
rect 472216 57876 472222 57928
rect 480346 57876 480352 57928
rect 480404 57916 480410 57928
rect 480530 57916 480536 57928
rect 480404 57888 480536 57916
rect 480404 57876 480410 57888
rect 480530 57876 480536 57888
rect 480588 57876 480594 57928
rect 298370 57848 298376 57860
rect 298296 57820 298376 57848
rect 298370 57808 298376 57820
rect 298428 57808 298434 57860
rect 287238 56692 287244 56704
rect 287199 56664 287244 56692
rect 287238 56652 287244 56664
rect 287296 56652 287302 56704
rect 283098 56624 283104 56636
rect 283059 56596 283104 56624
rect 283098 56584 283104 56596
rect 283156 56584 283162 56636
rect 324498 56624 324504 56636
rect 324459 56596 324504 56624
rect 324498 56584 324504 56596
rect 324556 56584 324562 56636
rect 375469 56627 375527 56633
rect 375469 56593 375481 56627
rect 375515 56624 375527 56627
rect 375558 56624 375564 56636
rect 375515 56596 375564 56624
rect 375515 56593 375527 56596
rect 375469 56587 375527 56593
rect 375558 56584 375564 56596
rect 375616 56584 375622 56636
rect 407758 56624 407764 56636
rect 407719 56596 407764 56624
rect 407758 56584 407764 56596
rect 407816 56584 407822 56636
rect 240226 56556 240232 56568
rect 240187 56528 240232 56556
rect 240226 56516 240232 56528
rect 240284 56516 240290 56568
rect 249886 56556 249892 56568
rect 249847 56528 249892 56556
rect 249886 56516 249892 56528
rect 249944 56516 249950 56568
rect 281629 56559 281687 56565
rect 281629 56525 281641 56559
rect 281675 56556 281687 56559
rect 281718 56556 281724 56568
rect 281675 56528 281724 56556
rect 281675 56525 281687 56528
rect 281629 56519 281687 56525
rect 281718 56516 281724 56528
rect 281776 56516 281782 56568
rect 287238 56556 287244 56568
rect 287199 56528 287244 56556
rect 287238 56516 287244 56528
rect 287296 56516 287302 56568
rect 329926 56516 329932 56568
rect 329984 56556 329990 56568
rect 330018 56556 330024 56568
rect 329984 56528 330024 56556
rect 329984 56516 329990 56528
rect 330018 56516 330024 56528
rect 330076 56516 330082 56568
rect 353478 56516 353484 56568
rect 353536 56556 353542 56568
rect 353662 56556 353668 56568
rect 353536 56528 353668 56556
rect 353536 56516 353542 56528
rect 353662 56516 353668 56528
rect 353720 56516 353726 56568
rect 397733 56559 397791 56565
rect 397733 56525 397745 56559
rect 397779 56556 397791 56559
rect 397822 56556 397828 56568
rect 397779 56528 397828 56556
rect 397779 56525 397791 56528
rect 397733 56519 397791 56525
rect 397822 56516 397828 56528
rect 397880 56516 397886 56568
rect 375558 56488 375564 56500
rect 375519 56460 375564 56488
rect 375558 56448 375564 56460
rect 375616 56448 375622 56500
rect 255498 55264 255504 55276
rect 255459 55236 255504 55264
rect 255498 55224 255504 55236
rect 255556 55224 255562 55276
rect 266814 55224 266820 55276
rect 266872 55264 266878 55276
rect 266998 55264 267004 55276
rect 266872 55236 267004 55264
rect 266872 55224 266878 55236
rect 266998 55224 267004 55236
rect 267056 55224 267062 55276
rect 310609 55267 310667 55273
rect 310609 55233 310621 55267
rect 310655 55264 310667 55267
rect 310882 55264 310888 55276
rect 310655 55236 310888 55264
rect 310655 55233 310667 55236
rect 310609 55227 310667 55233
rect 310882 55224 310888 55236
rect 310940 55224 310946 55276
rect 298370 55156 298376 55208
rect 298428 55196 298434 55208
rect 298462 55196 298468 55208
rect 298428 55168 298468 55196
rect 298428 55156 298434 55168
rect 298462 55156 298468 55168
rect 298520 55156 298526 55208
rect 329926 55196 329932 55208
rect 329887 55168 329932 55196
rect 329926 55156 329932 55168
rect 329984 55156 329990 55208
rect 342441 55199 342499 55205
rect 342441 55165 342453 55199
rect 342487 55196 342499 55199
rect 342530 55196 342536 55208
rect 342487 55168 342536 55196
rect 342487 55165 342499 55168
rect 342441 55159 342499 55165
rect 342530 55156 342536 55168
rect 342588 55156 342594 55208
rect 367278 55156 367284 55208
rect 367336 55196 367342 55208
rect 367370 55196 367376 55208
rect 367336 55168 367376 55196
rect 367336 55156 367342 55168
rect 367370 55156 367376 55168
rect 367428 55156 367434 55208
rect 266998 55128 267004 55140
rect 266959 55100 267004 55128
rect 266998 55088 267004 55100
rect 267056 55088 267062 55140
rect 359182 53836 359188 53848
rect 359143 53808 359188 53836
rect 359182 53796 359188 53808
rect 359240 53796 359246 53848
rect 271969 51799 272027 51805
rect 271969 51765 271981 51799
rect 272015 51796 272027 51799
rect 272058 51796 272064 51808
rect 272015 51768 272064 51796
rect 272015 51765 272027 51768
rect 271969 51759 272027 51765
rect 272058 51756 272064 51768
rect 272116 51756 272122 51808
rect 375561 51731 375619 51737
rect 375561 51697 375573 51731
rect 375607 51728 375619 51731
rect 375650 51728 375656 51740
rect 375607 51700 375656 51728
rect 375607 51697 375619 51700
rect 375561 51691 375619 51697
rect 375650 51688 375656 51700
rect 375708 51688 375714 51740
rect 249886 51184 249892 51196
rect 249847 51156 249892 51184
rect 249886 51144 249892 51156
rect 249944 51144 249950 51196
rect 305178 51184 305184 51196
rect 305104 51156 305184 51184
rect 261018 51076 261024 51128
rect 261076 51076 261082 51128
rect 261036 50992 261064 51076
rect 305104 51060 305132 51156
rect 305178 51144 305184 51156
rect 305236 51144 305242 51196
rect 321738 51184 321744 51196
rect 321699 51156 321744 51184
rect 321738 51144 321744 51156
rect 321796 51144 321802 51196
rect 309318 51076 309324 51128
rect 309376 51076 309382 51128
rect 327258 51076 327264 51128
rect 327316 51076 327322 51128
rect 382369 51119 382427 51125
rect 382369 51085 382381 51119
rect 382415 51116 382427 51119
rect 382458 51116 382464 51128
rect 382415 51088 382464 51116
rect 382415 51085 382427 51088
rect 382369 51079 382427 51085
rect 382458 51076 382464 51088
rect 382516 51076 382522 51128
rect 392210 51116 392216 51128
rect 392136 51088 392216 51116
rect 305086 51008 305092 51060
rect 305144 51008 305150 51060
rect 261018 50940 261024 50992
rect 261076 50940 261082 50992
rect 309336 50980 309364 51076
rect 327276 50992 327304 51076
rect 392136 51060 392164 51088
rect 392210 51076 392216 51088
rect 392268 51076 392274 51128
rect 408678 51076 408684 51128
rect 408736 51116 408742 51128
rect 408736 51088 408816 51116
rect 408736 51076 408742 51088
rect 408788 51060 408816 51088
rect 392118 51008 392124 51060
rect 392176 51008 392182 51060
rect 408770 51008 408776 51060
rect 408828 51008 408834 51060
rect 309410 50980 309416 50992
rect 309336 50952 309416 50980
rect 309410 50940 309416 50952
rect 309468 50940 309474 50992
rect 327258 50940 327264 50992
rect 327316 50940 327322 50992
rect 236362 48396 236368 48408
rect 236288 48368 236368 48396
rect 236288 48340 236316 48368
rect 236362 48356 236368 48368
rect 236420 48356 236426 48408
rect 332778 48396 332784 48408
rect 332704 48368 332784 48396
rect 233418 48288 233424 48340
rect 233476 48328 233482 48340
rect 233510 48328 233516 48340
rect 233476 48300 233516 48328
rect 233476 48288 233482 48300
rect 233510 48288 233516 48300
rect 233568 48288 233574 48340
rect 236270 48288 236276 48340
rect 236328 48288 236334 48340
rect 331401 48331 331459 48337
rect 331401 48297 331413 48331
rect 331447 48328 331459 48331
rect 331490 48328 331496 48340
rect 331447 48300 331496 48328
rect 331447 48297 331459 48300
rect 331401 48291 331459 48297
rect 331490 48288 331496 48300
rect 331548 48288 331554 48340
rect 332704 48272 332732 48368
rect 332778 48356 332784 48368
rect 332836 48356 332842 48408
rect 352098 48396 352104 48408
rect 352024 48368 352104 48396
rect 352024 48340 352052 48368
rect 352098 48356 352104 48368
rect 352156 48356 352162 48408
rect 359093 48399 359151 48405
rect 359093 48365 359105 48399
rect 359139 48396 359151 48399
rect 359182 48396 359188 48408
rect 359139 48368 359188 48396
rect 359139 48365 359151 48368
rect 359093 48359 359151 48365
rect 359182 48356 359188 48368
rect 359240 48356 359246 48408
rect 416866 48396 416872 48408
rect 416827 48368 416872 48396
rect 416866 48356 416872 48368
rect 416924 48356 416930 48408
rect 334345 48331 334403 48337
rect 334345 48297 334357 48331
rect 334391 48328 334403 48331
rect 334434 48328 334440 48340
rect 334391 48300 334440 48328
rect 334391 48297 334403 48300
rect 334345 48291 334403 48297
rect 334434 48288 334440 48300
rect 334492 48288 334498 48340
rect 352006 48288 352012 48340
rect 352064 48288 352070 48340
rect 382366 48328 382372 48340
rect 382327 48300 382372 48328
rect 382366 48288 382372 48300
rect 382424 48288 382430 48340
rect 393130 48288 393136 48340
rect 393188 48328 393194 48340
rect 393222 48328 393228 48340
rect 393188 48300 393228 48328
rect 393188 48288 393194 48300
rect 393222 48288 393228 48300
rect 393280 48288 393286 48340
rect 422386 48288 422392 48340
rect 422444 48328 422450 48340
rect 422478 48328 422484 48340
rect 422444 48300 422484 48328
rect 422444 48288 422450 48300
rect 422478 48288 422484 48300
rect 422536 48288 422542 48340
rect 433610 48328 433616 48340
rect 433571 48300 433616 48328
rect 433610 48288 433616 48300
rect 433668 48288 433674 48340
rect 466546 48328 466552 48340
rect 466507 48300 466552 48328
rect 466546 48288 466552 48300
rect 466604 48288 466610 48340
rect 472066 48328 472072 48340
rect 472027 48300 472072 48328
rect 472066 48288 472072 48300
rect 472124 48288 472130 48340
rect 332686 48220 332692 48272
rect 332744 48220 332750 48272
rect 380986 48220 380992 48272
rect 381044 48260 381050 48272
rect 381170 48260 381176 48272
rect 381044 48232 381176 48260
rect 381044 48220 381050 48232
rect 381170 48220 381176 48232
rect 381228 48220 381234 48272
rect 386690 48220 386696 48272
rect 386748 48260 386754 48272
rect 386782 48260 386788 48272
rect 386748 48232 386788 48260
rect 386748 48220 386754 48232
rect 386782 48220 386788 48232
rect 386840 48220 386846 48272
rect 392118 48260 392124 48272
rect 392079 48232 392124 48260
rect 392118 48220 392124 48232
rect 392176 48220 392182 48272
rect 416866 48220 416872 48272
rect 416924 48260 416930 48272
rect 417050 48260 417056 48272
rect 416924 48232 417056 48260
rect 416924 48220 416930 48232
rect 417050 48220 417056 48232
rect 417108 48220 417114 48272
rect 400582 47172 400588 47184
rect 400543 47144 400588 47172
rect 400582 47132 400588 47144
rect 400640 47132 400646 47184
rect 249886 47036 249892 47048
rect 249847 47008 249892 47036
rect 249886 46996 249892 47008
rect 249944 46996 249950 47048
rect 270678 47036 270684 47048
rect 270604 47008 270684 47036
rect 270604 46980 270632 47008
rect 270678 46996 270684 47008
rect 270736 46996 270742 47048
rect 287238 47036 287244 47048
rect 287199 47008 287244 47036
rect 287238 46996 287244 47008
rect 287296 46996 287302 47048
rect 292761 47039 292819 47045
rect 292761 47005 292773 47039
rect 292807 47036 292819 47039
rect 292850 47036 292856 47048
rect 292807 47008 292856 47036
rect 292807 47005 292819 47008
rect 292761 46999 292819 47005
rect 292850 46996 292856 47008
rect 292908 46996 292914 47048
rect 321738 47036 321744 47048
rect 321699 47008 321744 47036
rect 321738 46996 321744 47008
rect 321796 46996 321802 47048
rect 240226 46968 240232 46980
rect 240187 46940 240232 46968
rect 240226 46928 240232 46940
rect 240284 46928 240290 46980
rect 270586 46928 270592 46980
rect 270644 46928 270650 46980
rect 271966 46968 271972 46980
rect 271927 46940 271972 46968
rect 271966 46928 271972 46940
rect 272024 46928 272030 46980
rect 281626 46968 281632 46980
rect 281587 46940 281632 46968
rect 281626 46928 281632 46940
rect 281684 46928 281690 46980
rect 329929 46971 329987 46977
rect 329929 46937 329941 46971
rect 329975 46968 329987 46971
rect 330018 46968 330024 46980
rect 329975 46940 330024 46968
rect 329975 46937 329987 46940
rect 329929 46931 329987 46937
rect 330018 46928 330024 46940
rect 330076 46928 330082 46980
rect 347958 46928 347964 46980
rect 348016 46968 348022 46980
rect 348142 46968 348148 46980
rect 348016 46940 348148 46968
rect 348016 46928 348022 46940
rect 348142 46928 348148 46940
rect 348200 46928 348206 46980
rect 370038 46928 370044 46980
rect 370096 46968 370102 46980
rect 370130 46968 370136 46980
rect 370096 46940 370136 46968
rect 370096 46928 370102 46940
rect 370130 46928 370136 46940
rect 370188 46928 370194 46980
rect 397730 46968 397736 46980
rect 397691 46940 397736 46968
rect 397730 46928 397736 46940
rect 397788 46928 397794 46980
rect 451366 46928 451372 46980
rect 451424 46968 451430 46980
rect 451642 46968 451648 46980
rect 451424 46940 451648 46968
rect 451424 46928 451430 46940
rect 451642 46928 451648 46940
rect 451700 46928 451706 46980
rect 231946 46900 231952 46912
rect 231907 46872 231952 46900
rect 231946 46860 231952 46872
rect 232004 46860 232010 46912
rect 236270 46900 236276 46912
rect 236231 46872 236276 46900
rect 236270 46860 236276 46872
rect 236328 46860 236334 46912
rect 244458 46900 244464 46912
rect 244419 46872 244464 46900
rect 244458 46860 244464 46872
rect 244516 46860 244522 46912
rect 249886 46900 249892 46912
rect 249847 46872 249892 46900
rect 249886 46860 249892 46872
rect 249944 46860 249950 46912
rect 288526 46860 288532 46912
rect 288584 46900 288590 46912
rect 288618 46900 288624 46912
rect 288584 46872 288624 46900
rect 288584 46860 288590 46872
rect 288618 46860 288624 46872
rect 288676 46860 288682 46912
rect 309321 46903 309379 46909
rect 309321 46869 309333 46903
rect 309367 46900 309379 46903
rect 309410 46900 309416 46912
rect 309367 46872 309416 46900
rect 309367 46869 309379 46872
rect 309321 46863 309379 46869
rect 309410 46860 309416 46872
rect 309468 46860 309474 46912
rect 321646 46860 321652 46912
rect 321704 46900 321710 46912
rect 321738 46900 321744 46912
rect 321704 46872 321744 46900
rect 321704 46860 321710 46872
rect 321738 46860 321744 46872
rect 321796 46860 321802 46912
rect 407758 46900 407764 46912
rect 407719 46872 407764 46900
rect 407758 46860 407764 46872
rect 407816 46860 407822 46912
rect 255590 45568 255596 45620
rect 255648 45608 255654 45620
rect 255774 45608 255780 45620
rect 255648 45580 255780 45608
rect 255648 45568 255654 45580
rect 255774 45568 255780 45580
rect 255832 45568 255838 45620
rect 267001 45611 267059 45617
rect 267001 45577 267013 45611
rect 267047 45608 267059 45611
rect 267090 45608 267096 45620
rect 267047 45580 267096 45608
rect 267047 45577 267059 45580
rect 267001 45571 267059 45577
rect 267090 45568 267096 45580
rect 267148 45568 267154 45620
rect 342438 45608 342444 45620
rect 342399 45580 342444 45608
rect 342438 45568 342444 45580
rect 342496 45568 342502 45620
rect 356514 45608 356520 45620
rect 356475 45580 356520 45608
rect 356514 45568 356520 45580
rect 356572 45568 356578 45620
rect 359090 45608 359096 45620
rect 359051 45580 359096 45608
rect 359090 45568 359096 45580
rect 359148 45568 359154 45620
rect 400582 45608 400588 45620
rect 400543 45580 400588 45608
rect 400582 45568 400588 45580
rect 400640 45568 400646 45620
rect 282917 45543 282975 45549
rect 282917 45509 282929 45543
rect 282963 45540 282975 45543
rect 283190 45540 283196 45552
rect 282963 45512 283196 45540
rect 282963 45509 282975 45512
rect 282917 45503 282975 45509
rect 283190 45500 283196 45512
rect 283248 45500 283254 45552
rect 292850 45540 292856 45552
rect 292811 45512 292856 45540
rect 292850 45500 292856 45512
rect 292908 45500 292914 45552
rect 353570 45540 353576 45552
rect 353531 45512 353576 45540
rect 353570 45500 353576 45512
rect 353628 45500 353634 45552
rect 408678 45500 408684 45552
rect 408736 45540 408742 45552
rect 408770 45540 408776 45552
rect 408736 45512 408776 45540
rect 408736 45500 408742 45512
rect 408770 45500 408776 45512
rect 408828 45500 408834 45552
rect 400674 45472 400680 45484
rect 400635 45444 400680 45472
rect 400674 45432 400680 45444
rect 400732 45432 400738 45484
rect 330018 44112 330024 44124
rect 329979 44084 330024 44112
rect 330018 44072 330024 44084
rect 330076 44072 330082 44124
rect 271966 42916 271972 42968
rect 272024 42956 272030 42968
rect 272061 42959 272119 42965
rect 272061 42956 272073 42959
rect 272024 42928 272073 42956
rect 272024 42916 272030 42928
rect 272061 42925 272073 42928
rect 272107 42925 272119 42959
rect 272061 42919 272119 42925
rect 267090 42072 267096 42084
rect 267051 42044 267096 42072
rect 267090 42032 267096 42044
rect 267148 42032 267154 42084
rect 332686 42032 332692 42084
rect 332744 42072 332750 42084
rect 332870 42072 332876 42084
rect 332744 42044 332876 42072
rect 332744 42032 332750 42044
rect 332870 42032 332876 42044
rect 332928 42032 332934 42084
rect 357529 41463 357587 41469
rect 357529 41429 357541 41463
rect 357575 41460 357587 41463
rect 357618 41460 357624 41472
rect 357575 41432 357624 41460
rect 357575 41429 357587 41432
rect 357529 41423 357587 41429
rect 357618 41420 357624 41432
rect 357676 41420 357682 41472
rect 471974 41352 471980 41404
rect 472032 41392 472038 41404
rect 472158 41392 472164 41404
rect 472032 41364 472164 41392
rect 472032 41352 472038 41364
rect 472158 41352 472164 41364
rect 472216 41352 472222 41404
rect 451366 41284 451372 41336
rect 451424 41324 451430 41336
rect 451734 41324 451740 41336
rect 451424 41296 451740 41324
rect 451424 41284 451430 41296
rect 451734 41284 451740 41296
rect 451792 41284 451798 41336
rect 356514 40740 356520 40792
rect 356572 40780 356578 40792
rect 356609 40783 356667 40789
rect 356609 40780 356621 40783
rect 356572 40752 356621 40780
rect 356572 40740 356578 40752
rect 356609 40749 356621 40752
rect 356655 40749 356667 40783
rect 356609 40743 356667 40749
rect 267734 40332 267740 40384
rect 267792 40372 267798 40384
rect 277302 40372 277308 40384
rect 267792 40344 277308 40372
rect 267792 40332 267798 40344
rect 277302 40332 277308 40344
rect 277360 40332 277366 40384
rect 402974 40332 402980 40384
rect 403032 40372 403038 40384
rect 412450 40372 412456 40384
rect 403032 40344 412456 40372
rect 403032 40332 403038 40344
rect 412450 40332 412456 40344
rect 412508 40332 412514 40384
rect 252738 40168 252744 40180
rect 252699 40140 252744 40168
rect 252738 40128 252744 40140
rect 252796 40128 252802 40180
rect 324498 40168 324504 40180
rect 324459 40140 324504 40168
rect 324498 40128 324504 40140
rect 324556 40128 324562 40180
rect 311802 40060 311808 40112
rect 311860 40100 311866 40112
rect 317322 40100 317328 40112
rect 311860 40072 317328 40100
rect 311860 40060 311866 40072
rect 317322 40060 317328 40072
rect 317380 40060 317386 40112
rect 521654 40060 521660 40112
rect 521712 40100 521718 40112
rect 526438 40100 526444 40112
rect 521712 40072 526444 40100
rect 521712 40060 521718 40072
rect 526438 40060 526444 40072
rect 526496 40060 526502 40112
rect 480254 38700 480260 38752
rect 480312 38740 480318 38752
rect 480530 38740 480536 38752
rect 480312 38712 480536 38740
rect 480312 38700 480318 38712
rect 480530 38700 480536 38712
rect 480588 38700 480594 38752
rect 376846 38632 376852 38684
rect 376904 38672 376910 38684
rect 376938 38672 376944 38684
rect 376904 38644 376944 38672
rect 376904 38632 376910 38644
rect 376938 38632 376944 38644
rect 376996 38632 377002 38684
rect 382366 38632 382372 38684
rect 382424 38672 382430 38684
rect 382458 38672 382464 38684
rect 382424 38644 382464 38672
rect 382424 38632 382430 38644
rect 382458 38632 382464 38644
rect 382516 38632 382522 38684
rect 472158 38604 472164 38616
rect 472119 38576 472164 38604
rect 472158 38564 472164 38576
rect 472216 38564 472222 38616
rect 231949 37315 232007 37321
rect 231949 37281 231961 37315
rect 231995 37312 232007 37315
rect 232038 37312 232044 37324
rect 231995 37284 232044 37312
rect 231995 37281 232007 37284
rect 231949 37275 232007 37281
rect 232038 37272 232044 37284
rect 232096 37272 232102 37324
rect 236273 37315 236331 37321
rect 236273 37281 236285 37315
rect 236319 37312 236331 37315
rect 236362 37312 236368 37324
rect 236319 37284 236368 37312
rect 236319 37281 236331 37284
rect 236273 37275 236331 37281
rect 236362 37272 236368 37284
rect 236420 37272 236426 37324
rect 244461 37315 244519 37321
rect 244461 37281 244473 37315
rect 244507 37312 244519 37315
rect 244550 37312 244556 37324
rect 244507 37284 244556 37312
rect 244507 37281 244519 37284
rect 244461 37275 244519 37281
rect 244550 37272 244556 37284
rect 244608 37272 244614 37324
rect 249886 37312 249892 37324
rect 249847 37284 249892 37312
rect 249886 37272 249892 37284
rect 249944 37272 249950 37324
rect 287238 37272 287244 37324
rect 287296 37312 287302 37324
rect 287330 37312 287336 37324
rect 287296 37284 287336 37312
rect 287296 37272 287302 37284
rect 287330 37272 287336 37284
rect 287388 37272 287394 37324
rect 295518 37272 295524 37324
rect 295576 37312 295582 37324
rect 295702 37312 295708 37324
rect 295576 37284 295708 37312
rect 295576 37272 295582 37284
rect 295702 37272 295708 37284
rect 295760 37272 295766 37324
rect 309318 37312 309324 37324
rect 309279 37284 309324 37312
rect 309318 37272 309324 37284
rect 309376 37272 309382 37324
rect 310606 37272 310612 37324
rect 310664 37312 310670 37324
rect 310790 37312 310796 37324
rect 310664 37284 310796 37312
rect 310664 37272 310670 37284
rect 310790 37272 310796 37284
rect 310848 37272 310854 37324
rect 331398 37272 331404 37324
rect 331456 37312 331462 37324
rect 331490 37312 331496 37324
rect 331456 37284 331496 37312
rect 331456 37272 331462 37284
rect 331490 37272 331496 37284
rect 331548 37272 331554 37324
rect 334342 37272 334348 37324
rect 334400 37312 334406 37324
rect 334434 37312 334440 37324
rect 334400 37284 334440 37312
rect 334400 37272 334406 37284
rect 334434 37272 334440 37284
rect 334492 37272 334498 37324
rect 352006 37272 352012 37324
rect 352064 37312 352070 37324
rect 352098 37312 352104 37324
rect 352064 37284 352104 37312
rect 352064 37272 352070 37284
rect 352098 37272 352104 37284
rect 352156 37272 352162 37324
rect 407758 37312 407764 37324
rect 407719 37284 407764 37312
rect 407758 37272 407764 37284
rect 407816 37272 407822 37324
rect 353570 37244 353576 37256
rect 353531 37216 353576 37244
rect 353570 37204 353576 37216
rect 353628 37204 353634 37256
rect 400674 37176 400680 37188
rect 400635 37148 400680 37176
rect 400674 37136 400680 37148
rect 400732 37136 400738 37188
rect 364610 36020 364616 36032
rect 364536 35992 364616 36020
rect 364536 35964 364564 35992
rect 364610 35980 364616 35992
rect 364668 35980 364674 36032
rect 282914 35952 282920 35964
rect 282875 35924 282920 35952
rect 282914 35912 282920 35924
rect 282972 35912 282978 35964
rect 292850 35952 292856 35964
rect 292811 35924 292856 35952
rect 292850 35912 292856 35924
rect 292908 35912 292914 35964
rect 347866 35912 347872 35964
rect 347924 35952 347930 35964
rect 348142 35952 348148 35964
rect 347924 35924 348148 35952
rect 347924 35912 347930 35924
rect 348142 35912 348148 35924
rect 348200 35912 348206 35964
rect 356606 35952 356612 35964
rect 356567 35924 356612 35952
rect 356606 35912 356612 35924
rect 356664 35912 356670 35964
rect 357526 35952 357532 35964
rect 357487 35924 357532 35952
rect 357526 35912 357532 35924
rect 357584 35912 357590 35964
rect 364518 35912 364524 35964
rect 364576 35912 364582 35964
rect 367370 35912 367376 35964
rect 367428 35952 367434 35964
rect 367462 35952 367468 35964
rect 367428 35924 367468 35952
rect 367428 35912 367434 35924
rect 367462 35912 367468 35924
rect 367520 35912 367526 35964
rect 370038 35912 370044 35964
rect 370096 35952 370102 35964
rect 370130 35952 370136 35964
rect 370096 35924 370136 35952
rect 370096 35912 370102 35924
rect 370130 35912 370136 35924
rect 370188 35912 370194 35964
rect 392121 35955 392179 35961
rect 392121 35921 392133 35955
rect 392167 35952 392179 35955
rect 392210 35952 392216 35964
rect 392167 35924 392216 35952
rect 392167 35921 392179 35924
rect 392121 35915 392179 35921
rect 392210 35912 392216 35924
rect 392268 35912 392274 35964
rect 3510 35844 3516 35896
rect 3568 35884 3574 35896
rect 7558 35884 7564 35896
rect 3568 35856 7564 35884
rect 3568 35844 3574 35856
rect 7558 35844 7564 35856
rect 7616 35844 7622 35896
rect 231857 35887 231915 35893
rect 231857 35853 231869 35887
rect 231903 35884 231915 35887
rect 232038 35884 232044 35896
rect 231903 35856 232044 35884
rect 231903 35853 231915 35856
rect 231857 35847 231915 35853
rect 232038 35844 232044 35856
rect 232096 35844 232102 35896
rect 358906 35844 358912 35896
rect 358964 35884 358970 35896
rect 359090 35884 359096 35896
rect 358964 35856 359096 35884
rect 358964 35844 358970 35856
rect 359090 35844 359096 35856
rect 359148 35844 359154 35896
rect 375558 35844 375564 35896
rect 375616 35884 375622 35896
rect 375742 35884 375748 35896
rect 375616 35856 375748 35884
rect 375616 35844 375622 35856
rect 375742 35844 375748 35856
rect 375800 35844 375806 35896
rect 342349 32419 342407 32425
rect 342349 32385 342361 32419
rect 342395 32416 342407 32419
rect 342438 32416 342444 32428
rect 342395 32388 342444 32416
rect 342395 32385 342407 32388
rect 342349 32379 342407 32385
rect 342438 32376 342444 32388
rect 342496 32376 342502 32428
rect 240226 31872 240232 31884
rect 240187 31844 240232 31872
rect 240226 31832 240232 31844
rect 240284 31832 240290 31884
rect 408770 31804 408776 31816
rect 408696 31776 408776 31804
rect 408696 31748 408724 31776
rect 408770 31764 408776 31776
rect 408828 31764 408834 31816
rect 416958 31804 416964 31816
rect 416884 31776 416964 31804
rect 416884 31748 416912 31776
rect 416958 31764 416964 31776
rect 417016 31764 417022 31816
rect 451734 31804 451740 31816
rect 451660 31776 451740 31804
rect 451660 31748 451688 31776
rect 451734 31764 451740 31776
rect 451792 31764 451798 31816
rect 480254 31764 480260 31816
rect 480312 31764 480318 31816
rect 408678 31696 408684 31748
rect 408736 31696 408742 31748
rect 416866 31696 416872 31748
rect 416924 31696 416930 31748
rect 451642 31696 451648 31748
rect 451700 31696 451706 31748
rect 252741 31671 252799 31677
rect 252741 31637 252753 31671
rect 252787 31668 252799 31671
rect 252830 31668 252836 31680
rect 252787 31640 252836 31668
rect 252787 31637 252799 31640
rect 252741 31631 252799 31637
rect 252830 31628 252836 31640
rect 252888 31628 252894 31680
rect 480272 31668 480300 31764
rect 480346 31668 480352 31680
rect 480272 31640 480352 31668
rect 480346 31628 480352 31640
rect 480404 31628 480410 31680
rect 472158 31192 472164 31204
rect 472119 31164 472164 31192
rect 472158 31152 472164 31164
rect 472216 31152 472222 31204
rect 356517 31127 356575 31133
rect 356517 31093 356529 31127
rect 356563 31124 356575 31127
rect 356606 31124 356612 31136
rect 356563 31096 356612 31124
rect 356563 31093 356575 31096
rect 356517 31087 356575 31093
rect 356606 31084 356612 31096
rect 356664 31084 356670 31136
rect 278774 29180 278780 29232
rect 278832 29220 278838 29232
rect 283098 29220 283104 29232
rect 278832 29192 283104 29220
rect 278832 29180 278838 29192
rect 283098 29180 283104 29192
rect 283156 29180 283162 29232
rect 466270 29180 466276 29232
rect 466328 29220 466334 29232
rect 473262 29220 473268 29232
rect 466328 29192 473268 29220
rect 466328 29180 466334 29192
rect 473262 29180 473268 29192
rect 473320 29180 473326 29232
rect 572622 29180 572628 29232
rect 572680 29220 572686 29232
rect 576762 29220 576768 29232
rect 572680 29192 576768 29220
rect 572680 29180 572686 29192
rect 576762 29180 576768 29192
rect 576820 29180 576826 29232
rect 261018 29084 261024 29096
rect 260944 29056 261024 29084
rect 260944 29028 260972 29056
rect 261018 29044 261024 29056
rect 261076 29044 261082 29096
rect 386782 29084 386788 29096
rect 386708 29056 386788 29084
rect 386708 29028 386736 29056
rect 386782 29044 386788 29056
rect 386840 29044 386846 29096
rect 521654 29044 521660 29096
rect 521712 29084 521718 29096
rect 525886 29084 525892 29096
rect 521712 29056 525892 29084
rect 521712 29044 521718 29056
rect 525886 29044 525892 29056
rect 525944 29044 525950 29096
rect 244366 28976 244372 29028
rect 244424 29016 244430 29028
rect 244550 29016 244556 29028
rect 244424 28988 244556 29016
rect 244424 28976 244430 28988
rect 244550 28976 244556 28988
rect 244608 28976 244614 29028
rect 249886 28976 249892 29028
rect 249944 29016 249950 29028
rect 249978 29016 249984 29028
rect 249944 28988 249984 29016
rect 249944 28976 249950 28988
rect 249978 28976 249984 28988
rect 250036 28976 250042 29028
rect 260926 28976 260932 29028
rect 260984 28976 260990 29028
rect 267090 29016 267096 29028
rect 267051 28988 267096 29016
rect 267090 28976 267096 28988
rect 267148 28976 267154 29028
rect 270678 28976 270684 29028
rect 270736 29016 270742 29028
rect 270770 29016 270776 29028
rect 270736 28988 270776 29016
rect 270736 28976 270742 28988
rect 270770 28976 270776 28988
rect 270828 28976 270834 29028
rect 272058 29016 272064 29028
rect 272019 28988 272064 29016
rect 272058 28976 272064 28988
rect 272116 28976 272122 29028
rect 321646 28976 321652 29028
rect 321704 29016 321710 29028
rect 321738 29016 321744 29028
rect 321704 28988 321744 29016
rect 321704 28976 321710 28988
rect 321738 28976 321744 28988
rect 321796 28976 321802 29028
rect 324498 29016 324504 29028
rect 324459 28988 324504 29016
rect 324498 28976 324504 28988
rect 324556 28976 324562 29028
rect 381078 28976 381084 29028
rect 381136 29016 381142 29028
rect 381170 29016 381176 29028
rect 381136 28988 381176 29016
rect 381136 28976 381142 28988
rect 381170 28976 381176 28988
rect 381228 28976 381234 29028
rect 386690 28976 386696 29028
rect 386748 28976 386754 29028
rect 387886 28976 387892 29028
rect 387944 29016 387950 29028
rect 388070 29016 388076 29028
rect 387944 28988 388076 29016
rect 387944 28976 387950 28988
rect 388070 28976 388076 28988
rect 388128 28976 388134 29028
rect 393130 28976 393136 29028
rect 393188 29016 393194 29028
rect 393222 29016 393228 29028
rect 393188 28988 393228 29016
rect 393188 28976 393194 28988
rect 393222 28976 393228 28988
rect 393280 28976 393286 29028
rect 243078 28908 243084 28960
rect 243136 28948 243142 28960
rect 243170 28948 243176 28960
rect 243136 28920 243176 28948
rect 243136 28908 243142 28920
rect 243170 28908 243176 28920
rect 243228 28908 243234 28960
rect 252830 28948 252836 28960
rect 252791 28920 252836 28948
rect 252830 28908 252836 28920
rect 252888 28908 252894 28960
rect 254210 28908 254216 28960
rect 254268 28948 254274 28960
rect 254302 28948 254308 28960
rect 254268 28920 254308 28948
rect 254268 28908 254274 28920
rect 254302 28908 254308 28920
rect 254360 28908 254366 28960
rect 259546 28908 259552 28960
rect 259604 28948 259610 28960
rect 259730 28948 259736 28960
rect 259604 28920 259736 28948
rect 259604 28908 259610 28920
rect 259730 28908 259736 28920
rect 259788 28908 259794 28960
rect 265158 28908 265164 28960
rect 265216 28948 265222 28960
rect 265250 28948 265256 28960
rect 265216 28920 265256 28948
rect 265216 28908 265222 28920
rect 265250 28908 265256 28920
rect 265308 28908 265314 28960
rect 266538 28908 266544 28960
rect 266596 28948 266602 28960
rect 266630 28948 266636 28960
rect 266596 28920 266636 28948
rect 266596 28908 266602 28920
rect 266630 28908 266636 28920
rect 266688 28908 266694 28960
rect 281718 28948 281724 28960
rect 281679 28920 281724 28948
rect 281718 28908 281724 28920
rect 281776 28908 281782 28960
rect 288434 28908 288440 28960
rect 288492 28948 288498 28960
rect 288618 28948 288624 28960
rect 288492 28920 288624 28948
rect 288492 28908 288498 28920
rect 288618 28908 288624 28920
rect 288676 28908 288682 28960
rect 293954 28908 293960 28960
rect 294012 28948 294018 28960
rect 294138 28948 294144 28960
rect 294012 28920 294144 28948
rect 294012 28908 294018 28920
rect 294138 28908 294144 28920
rect 294196 28908 294202 28960
rect 371234 28908 371240 28960
rect 371292 28948 371298 28960
rect 371418 28948 371424 28960
rect 371292 28920 371424 28948
rect 371292 28908 371298 28920
rect 371418 28908 371424 28920
rect 371476 28908 371482 28960
rect 427817 28951 427875 28957
rect 427817 28917 427829 28951
rect 427863 28948 427875 28951
rect 427906 28948 427912 28960
rect 427863 28920 427912 28948
rect 427863 28917 427875 28920
rect 427817 28911 427875 28917
rect 427906 28908 427912 28920
rect 427964 28908 427970 28960
rect 400490 28840 400496 28892
rect 400548 28880 400554 28892
rect 400674 28880 400680 28892
rect 400548 28852 400680 28880
rect 400548 28840 400554 28852
rect 400674 28840 400680 28852
rect 400732 28840 400738 28892
rect 422386 27616 422392 27668
rect 422444 27656 422450 27668
rect 422478 27656 422484 27668
rect 422444 27628 422484 27656
rect 422444 27616 422450 27628
rect 422478 27616 422484 27628
rect 422536 27616 422542 27668
rect 266630 27588 266636 27600
rect 266591 27560 266636 27588
rect 266630 27548 266636 27560
rect 266688 27548 266694 27600
rect 270681 27591 270739 27597
rect 270681 27557 270693 27591
rect 270727 27588 270739 27591
rect 270770 27588 270776 27600
rect 270727 27560 270776 27588
rect 270727 27557 270739 27560
rect 270681 27551 270739 27557
rect 270770 27548 270776 27560
rect 270828 27548 270834 27600
rect 318978 27588 318984 27600
rect 318939 27560 318984 27588
rect 318978 27548 318984 27560
rect 319036 27548 319042 27600
rect 324409 27591 324467 27597
rect 324409 27557 324421 27591
rect 324455 27588 324467 27591
rect 324498 27588 324504 27600
rect 324455 27560 324504 27588
rect 324455 27557 324467 27560
rect 324409 27551 324467 27557
rect 324498 27548 324504 27560
rect 324556 27548 324562 27600
rect 327166 27548 327172 27600
rect 327224 27588 327230 27600
rect 327258 27588 327264 27600
rect 327224 27560 327264 27588
rect 327224 27548 327230 27560
rect 327258 27548 327264 27560
rect 327316 27548 327322 27600
rect 331306 27548 331312 27600
rect 331364 27588 331370 27600
rect 331398 27588 331404 27600
rect 331364 27560 331404 27588
rect 331364 27548 331370 27560
rect 331398 27548 331404 27560
rect 331456 27548 331462 27600
rect 346486 27588 346492 27600
rect 346447 27560 346492 27588
rect 346486 27548 346492 27560
rect 346544 27548 346550 27600
rect 376846 27548 376852 27600
rect 376904 27588 376910 27600
rect 377030 27588 377036 27600
rect 376904 27560 377036 27588
rect 376904 27548 376910 27560
rect 377030 27548 377036 27560
rect 377088 27548 377094 27600
rect 382366 27548 382372 27600
rect 382424 27588 382430 27600
rect 382642 27588 382648 27600
rect 382424 27560 382648 27588
rect 382424 27548 382430 27560
rect 382642 27548 382648 27560
rect 382700 27548 382706 27600
rect 393222 27588 393228 27600
rect 393183 27560 393228 27588
rect 393222 27548 393228 27560
rect 393280 27548 393286 27600
rect 407758 27588 407764 27600
rect 407719 27560 407764 27588
rect 407758 27548 407764 27560
rect 407816 27548 407822 27600
rect 480346 27588 480352 27600
rect 480307 27560 480352 27588
rect 480346 27548 480352 27560
rect 480404 27548 480410 27600
rect 240226 26364 240232 26376
rect 240187 26336 240232 26364
rect 240226 26324 240232 26336
rect 240284 26324 240290 26376
rect 356514 26364 356520 26376
rect 356475 26336 356520 26364
rect 356514 26324 356520 26336
rect 356572 26324 356578 26376
rect 231854 26296 231860 26308
rect 231815 26268 231860 26296
rect 231854 26256 231860 26268
rect 231912 26256 231918 26308
rect 330021 26299 330079 26305
rect 330021 26265 330033 26299
rect 330067 26296 330079 26299
rect 330110 26296 330116 26308
rect 330067 26268 330116 26296
rect 330067 26265 330079 26268
rect 330021 26259 330079 26265
rect 330110 26256 330116 26268
rect 330168 26256 330174 26308
rect 236362 26228 236368 26240
rect 236323 26200 236368 26228
rect 236362 26188 236368 26200
rect 236420 26188 236426 26240
rect 240226 26188 240232 26240
rect 240284 26188 240290 26240
rect 347866 26228 347872 26240
rect 347827 26200 347872 26228
rect 347866 26188 347872 26200
rect 347924 26188 347930 26240
rect 357526 26228 357532 26240
rect 357487 26200 357532 26228
rect 357526 26188 357532 26200
rect 357584 26188 357590 26240
rect 358906 26188 358912 26240
rect 358964 26188 358970 26240
rect 364794 26228 364800 26240
rect 364755 26200 364800 26228
rect 364794 26188 364800 26200
rect 364852 26188 364858 26240
rect 392210 26228 392216 26240
rect 392171 26200 392216 26228
rect 392210 26188 392216 26200
rect 392268 26188 392274 26240
rect 231762 26120 231768 26172
rect 231820 26160 231826 26172
rect 231854 26160 231860 26172
rect 231820 26132 231860 26160
rect 231820 26120 231826 26132
rect 231854 26120 231860 26132
rect 231912 26120 231918 26172
rect 240244 26160 240272 26188
rect 240318 26160 240324 26172
rect 240244 26132 240324 26160
rect 240318 26120 240324 26132
rect 240376 26120 240382 26172
rect 358924 26160 358952 26188
rect 358998 26160 359004 26172
rect 358924 26132 359004 26160
rect 358998 26120 359004 26132
rect 359056 26120 359062 26172
rect 365714 22720 365720 22772
rect 365772 22760 365778 22772
rect 365990 22760 365996 22772
rect 365772 22732 365996 22760
rect 365772 22720 365778 22732
rect 365990 22720 365996 22732
rect 366048 22720 366054 22772
rect 422110 22516 422116 22568
rect 422168 22556 422174 22568
rect 422386 22556 422392 22568
rect 422168 22528 422392 22556
rect 422168 22516 422174 22528
rect 422386 22516 422392 22528
rect 422444 22516 422450 22568
rect 472158 22284 472164 22296
rect 472119 22256 472164 22284
rect 472158 22244 472164 22256
rect 472216 22244 472222 22296
rect 380802 22176 380808 22228
rect 380860 22216 380866 22228
rect 381170 22216 381176 22228
rect 380860 22188 381176 22216
rect 380860 22176 380866 22188
rect 381170 22176 381176 22188
rect 381228 22176 381234 22228
rect 277578 22148 277584 22160
rect 277504 22120 277584 22148
rect 277504 22092 277532 22120
rect 277578 22108 277584 22120
rect 277636 22108 277642 22160
rect 277486 22040 277492 22092
rect 277544 22040 277550 22092
rect 416774 22040 416780 22092
rect 416832 22080 416838 22092
rect 416958 22080 416964 22092
rect 416832 22052 416964 22080
rect 416832 22040 416838 22052
rect 416958 22040 416964 22052
rect 417016 22040 417022 22092
rect 244277 19431 244335 19437
rect 244277 19397 244289 19431
rect 244323 19428 244335 19431
rect 244366 19428 244372 19440
rect 244323 19400 244372 19428
rect 244323 19397 244335 19400
rect 244277 19391 244335 19397
rect 244366 19388 244372 19400
rect 244424 19388 244430 19440
rect 347869 19431 347927 19437
rect 347869 19397 347881 19431
rect 347915 19428 347927 19431
rect 347958 19428 347964 19440
rect 347915 19400 347964 19428
rect 347915 19397 347927 19400
rect 347869 19391 347927 19397
rect 347958 19388 347964 19400
rect 348016 19388 348022 19440
rect 427814 19428 427820 19440
rect 427775 19400 427820 19428
rect 427814 19388 427820 19400
rect 427872 19388 427878 19440
rect 252830 19360 252836 19372
rect 252791 19332 252836 19360
rect 252830 19320 252836 19332
rect 252888 19320 252894 19372
rect 260926 19320 260932 19372
rect 260984 19360 260990 19372
rect 261018 19360 261024 19372
rect 260984 19332 261024 19360
rect 260984 19320 260990 19332
rect 261018 19320 261024 19332
rect 261076 19320 261082 19372
rect 281718 19360 281724 19372
rect 281679 19332 281724 19360
rect 281718 19320 281724 19332
rect 281776 19320 281782 19372
rect 342346 19360 342352 19372
rect 342307 19332 342352 19360
rect 342346 19320 342352 19332
rect 342404 19320 342410 19372
rect 472158 19360 472164 19372
rect 472119 19332 472164 19360
rect 472158 19320 472164 19332
rect 472216 19320 472222 19372
rect 254302 19252 254308 19304
rect 254360 19252 254366 19304
rect 255590 19252 255596 19304
rect 255648 19252 255654 19304
rect 288526 19292 288532 19304
rect 288487 19264 288532 19292
rect 288526 19252 288532 19264
rect 288584 19252 288590 19304
rect 305086 19292 305092 19304
rect 305047 19264 305092 19292
rect 305086 19252 305092 19264
rect 305144 19252 305150 19304
rect 308030 19292 308036 19304
rect 307991 19264 308036 19292
rect 308030 19252 308036 19264
rect 308088 19252 308094 19304
rect 397549 19295 397607 19301
rect 397549 19261 397561 19295
rect 397595 19292 397607 19295
rect 397638 19292 397644 19304
rect 397595 19264 397644 19292
rect 397595 19261 397607 19264
rect 397549 19255 397607 19261
rect 397638 19252 397644 19264
rect 397696 19252 397702 19304
rect 427814 19292 427820 19304
rect 427775 19264 427820 19292
rect 427814 19252 427820 19264
rect 427872 19252 427878 19304
rect 254320 19168 254348 19252
rect 255608 19168 255636 19252
rect 266630 19224 266636 19236
rect 266591 19196 266636 19224
rect 266630 19184 266636 19196
rect 266688 19184 266694 19236
rect 254302 19116 254308 19168
rect 254360 19116 254366 19168
rect 255590 19116 255596 19168
rect 255648 19116 255654 19168
rect 272058 18068 272064 18080
rect 271984 18040 272064 18068
rect 271984 18012 272012 18040
rect 272058 18028 272064 18040
rect 272116 18028 272122 18080
rect 270678 18000 270684 18012
rect 270639 17972 270684 18000
rect 270678 17960 270684 17972
rect 270736 17960 270742 18012
rect 271966 17960 271972 18012
rect 272024 17960 272030 18012
rect 318978 18000 318984 18012
rect 318939 17972 318984 18000
rect 318978 17960 318984 17972
rect 319036 17960 319042 18012
rect 324406 18000 324412 18012
rect 324367 17972 324412 18000
rect 324406 17960 324412 17972
rect 324464 17960 324470 18012
rect 346486 18000 346492 18012
rect 346447 17972 346492 18000
rect 346486 17960 346492 17972
rect 346544 17960 346550 18012
rect 393222 18000 393228 18012
rect 393183 17972 393228 18000
rect 393222 17960 393228 17972
rect 393280 17960 393286 18012
rect 480346 18000 480352 18012
rect 480307 17972 480352 18000
rect 480346 17960 480352 17972
rect 480404 17960 480410 18012
rect 330110 17932 330116 17944
rect 330071 17904 330116 17932
rect 330110 17892 330116 17904
rect 330168 17892 330174 17944
rect 334342 17932 334348 17944
rect 334303 17904 334348 17932
rect 334342 17892 334348 17904
rect 334400 17892 334406 17944
rect 364794 17456 364800 17468
rect 364755 17428 364800 17456
rect 364794 17416 364800 17428
rect 364852 17416 364858 17468
rect 347682 16804 347688 16856
rect 347740 16844 347746 16856
rect 355962 16844 355968 16856
rect 347740 16816 355968 16844
rect 347740 16804 347746 16816
rect 355962 16804 355968 16816
rect 356020 16804 356026 16856
rect 514570 16736 514576 16788
rect 514628 16776 514634 16788
rect 516042 16776 516048 16788
rect 514628 16748 516048 16776
rect 514628 16736 514634 16748
rect 516042 16736 516048 16748
rect 516100 16736 516106 16788
rect 318702 16668 318708 16720
rect 318760 16708 318766 16720
rect 319622 16708 319628 16720
rect 318760 16680 319628 16708
rect 318760 16668 318766 16680
rect 319622 16668 319628 16680
rect 319680 16668 319686 16720
rect 334066 16668 334072 16720
rect 334124 16708 334130 16720
rect 338114 16708 338120 16720
rect 334124 16680 338120 16708
rect 334124 16668 334130 16680
rect 338114 16668 338120 16680
rect 338172 16668 338178 16720
rect 524230 16668 524236 16720
rect 524288 16708 524294 16720
rect 526438 16708 526444 16720
rect 524288 16680 526444 16708
rect 524288 16668 524294 16680
rect 526438 16668 526444 16680
rect 526496 16668 526502 16720
rect 236362 16640 236368 16652
rect 236323 16612 236368 16640
rect 236362 16600 236368 16612
rect 236420 16600 236426 16652
rect 244274 16640 244280 16652
rect 244235 16612 244280 16640
rect 244274 16600 244280 16612
rect 244332 16600 244338 16652
rect 392210 16640 392216 16652
rect 392171 16612 392216 16640
rect 392210 16600 392216 16612
rect 392268 16600 392274 16652
rect 125410 16328 125416 16380
rect 125468 16368 125474 16380
rect 292758 16368 292764 16380
rect 125468 16340 292764 16368
rect 125468 16328 125474 16340
rect 292758 16328 292764 16340
rect 292816 16328 292822 16380
rect 121362 16260 121368 16312
rect 121420 16300 121426 16312
rect 291286 16300 291292 16312
rect 121420 16272 291292 16300
rect 121420 16260 121426 16272
rect 291286 16260 291292 16272
rect 291344 16260 291350 16312
rect 114462 16192 114468 16244
rect 114520 16232 114526 16244
rect 287238 16232 287244 16244
rect 114520 16204 287244 16232
rect 114520 16192 114526 16204
rect 287238 16192 287244 16204
rect 287296 16192 287302 16244
rect 110322 16124 110328 16176
rect 110380 16164 110386 16176
rect 285766 16164 285772 16176
rect 110380 16136 285772 16164
rect 110380 16124 110386 16136
rect 285766 16124 285772 16136
rect 285824 16124 285830 16176
rect 107562 16056 107568 16108
rect 107620 16096 107626 16108
rect 284386 16096 284392 16108
rect 107620 16068 284392 16096
rect 107620 16056 107626 16068
rect 284386 16056 284392 16068
rect 284444 16056 284450 16108
rect 103422 15988 103428 16040
rect 103480 16028 103486 16040
rect 281718 16028 281724 16040
rect 103480 16000 281724 16028
rect 103480 15988 103486 16000
rect 281718 15988 281724 16000
rect 281776 15988 281782 16040
rect 31662 15920 31668 15972
rect 31720 15960 31726 15972
rect 245746 15960 245752 15972
rect 31720 15932 245752 15960
rect 31720 15920 31726 15932
rect 245746 15920 245752 15932
rect 245804 15920 245810 15972
rect 28902 15852 28908 15904
rect 28960 15892 28966 15904
rect 243078 15892 243084 15904
rect 28960 15864 243084 15892
rect 28960 15852 28966 15864
rect 243078 15852 243084 15864
rect 243136 15852 243142 15904
rect 336550 15172 336556 15224
rect 336608 15212 336614 15224
rect 336826 15212 336832 15224
rect 336608 15184 336832 15212
rect 336608 15172 336614 15184
rect 336826 15172 336832 15184
rect 336884 15172 336890 15224
rect 356330 15172 356336 15224
rect 356388 15212 356394 15224
rect 356422 15212 356428 15224
rect 356388 15184 356428 15212
rect 356388 15172 356394 15184
rect 356422 15172 356428 15184
rect 356480 15172 356486 15224
rect 129642 15104 129648 15156
rect 129700 15144 129706 15156
rect 295518 15144 295524 15156
rect 129700 15116 295524 15144
rect 129700 15104 129706 15116
rect 295518 15104 295524 15116
rect 295576 15104 295582 15156
rect 99282 15036 99288 15088
rect 99340 15076 99346 15088
rect 280246 15076 280252 15088
rect 99340 15048 280252 15076
rect 99340 15036 99346 15048
rect 280246 15036 280252 15048
rect 280304 15036 280310 15088
rect 96522 14968 96528 15020
rect 96580 15008 96586 15020
rect 278866 15008 278872 15020
rect 96580 14980 278872 15008
rect 96580 14968 96586 14980
rect 278866 14968 278872 14980
rect 278924 14968 278930 15020
rect 92382 14900 92388 14952
rect 92440 14940 92446 14952
rect 276106 14940 276112 14952
rect 92440 14912 276112 14940
rect 92440 14900 92446 14912
rect 276106 14900 276112 14912
rect 276164 14900 276170 14952
rect 89622 14832 89628 14884
rect 89680 14872 89686 14884
rect 274726 14872 274732 14884
rect 89680 14844 274732 14872
rect 89680 14832 89686 14844
rect 274726 14832 274732 14844
rect 274784 14832 274790 14884
rect 85482 14764 85488 14816
rect 85540 14804 85546 14816
rect 273346 14804 273352 14816
rect 85540 14776 273352 14804
rect 85540 14764 85546 14776
rect 273346 14764 273352 14776
rect 273404 14764 273410 14816
rect 82722 14696 82728 14748
rect 82780 14736 82786 14748
rect 270678 14736 270684 14748
rect 82780 14708 270684 14736
rect 82780 14696 82786 14708
rect 270678 14696 270684 14708
rect 270736 14696 270742 14748
rect 78582 14628 78588 14680
rect 78640 14668 78646 14680
rect 269206 14668 269212 14680
rect 78640 14640 269212 14668
rect 78640 14628 78646 14640
rect 269206 14628 269212 14640
rect 269264 14628 269270 14680
rect 392026 14628 392032 14680
rect 392084 14668 392090 14680
rect 392210 14668 392216 14680
rect 392084 14640 392216 14668
rect 392084 14628 392090 14640
rect 392210 14628 392216 14640
rect 392268 14628 392274 14680
rect 74442 14560 74448 14612
rect 74500 14600 74506 14612
rect 267826 14600 267832 14612
rect 74500 14572 267832 14600
rect 74500 14560 74506 14572
rect 267826 14560 267832 14572
rect 267884 14560 267890 14612
rect 71682 14492 71688 14544
rect 71740 14532 71746 14544
rect 265158 14532 265164 14544
rect 71740 14504 265164 14532
rect 71740 14492 71746 14504
rect 265158 14492 265164 14504
rect 265216 14492 265222 14544
rect 23382 14424 23388 14476
rect 23440 14464 23446 14476
rect 241698 14464 241704 14476
rect 23440 14436 241704 14464
rect 23440 14424 23446 14436
rect 241698 14424 241704 14436
rect 241756 14424 241762 14476
rect 244182 14424 244188 14476
rect 244240 14464 244246 14476
rect 354766 14464 354772 14476
rect 244240 14436 354772 14464
rect 244240 14424 244246 14436
rect 354766 14424 354772 14436
rect 354824 14424 354830 14476
rect 160002 14356 160008 14408
rect 160060 14396 160066 14408
rect 311986 14396 311992 14408
rect 160060 14368 311992 14396
rect 160060 14356 160066 14368
rect 311986 14356 311992 14368
rect 312044 14356 312050 14408
rect 157242 14288 157248 14340
rect 157300 14328 157306 14340
rect 309318 14328 309324 14340
rect 157300 14300 309324 14328
rect 157300 14288 157306 14300
rect 309318 14288 309324 14300
rect 309376 14288 309382 14340
rect 165522 14220 165528 14272
rect 165580 14260 165586 14272
rect 313458 14260 313464 14272
rect 165580 14232 313464 14260
rect 165580 14220 165586 14232
rect 313458 14220 313464 14232
rect 313516 14220 313522 14272
rect 168282 14152 168288 14204
rect 168340 14192 168346 14204
rect 316126 14192 316132 14204
rect 168340 14164 316132 14192
rect 168340 14152 168346 14164
rect 316126 14152 316132 14164
rect 316184 14152 316190 14204
rect 117222 14084 117228 14136
rect 117280 14124 117286 14136
rect 246298 14124 246304 14136
rect 117280 14096 246304 14124
rect 117280 14084 117286 14096
rect 246298 14084 246304 14096
rect 246356 14084 246362 14136
rect 240042 14016 240048 14068
rect 240100 14056 240106 14068
rect 352190 14056 352196 14068
rect 240100 14028 352196 14056
rect 240100 14016 240106 14028
rect 352190 14016 352196 14028
rect 352248 14016 352254 14068
rect 202782 13744 202788 13796
rect 202840 13784 202846 13796
rect 334158 13784 334164 13796
rect 202840 13756 334164 13784
rect 202840 13744 202846 13756
rect 334158 13744 334164 13756
rect 334216 13744 334222 13796
rect 159910 13676 159916 13728
rect 159968 13716 159974 13728
rect 310698 13716 310704 13728
rect 159968 13688 310704 13716
rect 159968 13676 159974 13688
rect 310698 13676 310704 13688
rect 310756 13676 310762 13728
rect 155862 13608 155868 13660
rect 155920 13648 155926 13660
rect 309134 13648 309140 13660
rect 155920 13620 309140 13648
rect 155920 13608 155926 13620
rect 309134 13608 309140 13620
rect 309192 13608 309198 13660
rect 153102 13540 153108 13592
rect 153160 13580 153166 13592
rect 307846 13580 307852 13592
rect 153160 13552 307852 13580
rect 153160 13540 153166 13552
rect 307846 13540 307852 13552
rect 307904 13540 307910 13592
rect 150342 13472 150348 13524
rect 150400 13512 150406 13524
rect 306466 13512 306472 13524
rect 150400 13484 306472 13512
rect 150400 13472 150406 13484
rect 306466 13472 306472 13484
rect 306524 13472 306530 13524
rect 148962 13404 148968 13456
rect 149020 13444 149026 13456
rect 305089 13447 305147 13453
rect 305089 13444 305101 13447
rect 149020 13416 305101 13444
rect 149020 13404 149026 13416
rect 305089 13413 305101 13416
rect 305135 13413 305147 13447
rect 305089 13407 305147 13413
rect 151722 13336 151728 13388
rect 151780 13376 151786 13388
rect 307938 13376 307944 13388
rect 151780 13348 307944 13376
rect 151780 13336 151786 13348
rect 307938 13336 307944 13348
rect 307996 13336 308002 13388
rect 146202 13268 146208 13320
rect 146260 13308 146266 13320
rect 303614 13308 303620 13320
rect 146260 13280 303620 13308
rect 146260 13268 146266 13280
rect 303614 13268 303620 13280
rect 303672 13268 303678 13320
rect 144822 13200 144828 13252
rect 144880 13240 144886 13252
rect 303706 13240 303712 13252
rect 144880 13212 303712 13240
rect 144880 13200 144886 13212
rect 303706 13200 303712 13212
rect 303764 13200 303770 13252
rect 132402 13132 132408 13184
rect 132460 13172 132466 13184
rect 296898 13172 296904 13184
rect 132460 13144 296904 13172
rect 132460 13132 132466 13144
rect 296898 13132 296904 13144
rect 296956 13132 296962 13184
rect 19242 13064 19248 13116
rect 19300 13104 19306 13116
rect 238846 13104 238852 13116
rect 19300 13076 238852 13104
rect 19300 13064 19306 13076
rect 238846 13064 238852 13076
rect 238904 13064 238910 13116
rect 382369 13107 382427 13113
rect 382369 13073 382381 13107
rect 382415 13104 382427 13107
rect 382642 13104 382648 13116
rect 382415 13076 382648 13104
rect 382415 13073 382427 13076
rect 382369 13067 382427 13073
rect 382642 13064 382648 13076
rect 382700 13064 382706 13116
rect 200022 12996 200028 13048
rect 200080 13036 200086 13048
rect 331306 13036 331312 13048
rect 200080 13008 331312 13036
rect 200080 12996 200086 13008
rect 331306 12996 331312 13008
rect 331364 12996 331370 13048
rect 206922 12928 206928 12980
rect 206980 12968 206986 12980
rect 335446 12968 335452 12980
rect 206980 12940 335452 12968
rect 206980 12928 206986 12940
rect 335446 12928 335452 12940
rect 335504 12928 335510 12980
rect 213822 12860 213828 12912
rect 213880 12900 213886 12912
rect 339678 12900 339684 12912
rect 213880 12872 339684 12900
rect 213880 12860 213886 12872
rect 339678 12860 339684 12872
rect 339736 12860 339742 12912
rect 211062 12792 211068 12844
rect 211120 12832 211126 12844
rect 336826 12832 336832 12844
rect 211120 12804 336832 12832
rect 211120 12792 211126 12804
rect 336826 12792 336832 12804
rect 336884 12792 336890 12844
rect 217962 12724 217968 12776
rect 218020 12764 218026 12776
rect 340966 12764 340972 12776
rect 218020 12736 340972 12764
rect 218020 12724 218026 12736
rect 340966 12724 340972 12736
rect 341024 12724 341030 12776
rect 220722 12656 220728 12708
rect 220780 12696 220786 12708
rect 342346 12696 342352 12708
rect 220780 12668 342352 12696
rect 220780 12656 220786 12668
rect 342346 12656 342352 12668
rect 342404 12656 342410 12708
rect 252741 12563 252799 12569
rect 252741 12529 252753 12563
rect 252787 12560 252799 12563
rect 252830 12560 252836 12572
rect 252787 12532 252836 12560
rect 252787 12529 252799 12532
rect 252741 12523 252799 12529
rect 252830 12520 252836 12532
rect 252888 12520 252894 12572
rect 293954 12492 293960 12504
rect 293915 12464 293960 12492
rect 293954 12452 293960 12464
rect 294012 12452 294018 12504
rect 347958 12492 347964 12504
rect 347884 12464 347964 12492
rect 347884 12436 347912 12464
rect 347958 12452 347964 12464
rect 348016 12452 348022 12504
rect 370038 12492 370044 12504
rect 369964 12464 370044 12492
rect 369964 12436 369992 12464
rect 370038 12452 370044 12464
rect 370096 12452 370102 12504
rect 393222 12492 393228 12504
rect 393056 12464 393228 12492
rect 393056 12436 393084 12464
rect 393222 12452 393228 12464
rect 393280 12452 393286 12504
rect 400490 12492 400496 12504
rect 400416 12464 400496 12492
rect 400416 12436 400444 12464
rect 400490 12452 400496 12464
rect 400548 12452 400554 12504
rect 184842 12384 184848 12436
rect 184900 12424 184906 12436
rect 323118 12424 323124 12436
rect 184900 12396 323124 12424
rect 184900 12384 184906 12396
rect 323118 12384 323124 12396
rect 323176 12384 323182 12436
rect 347866 12384 347872 12436
rect 347924 12384 347930 12436
rect 369946 12384 369952 12436
rect 370004 12384 370010 12436
rect 393038 12384 393044 12436
rect 393096 12384 393102 12436
rect 400398 12384 400404 12436
rect 400456 12384 400462 12436
rect 180702 12316 180708 12368
rect 180760 12356 180766 12368
rect 321738 12356 321744 12368
rect 180760 12328 321744 12356
rect 180760 12316 180766 12328
rect 321738 12316 321744 12328
rect 321796 12316 321802 12368
rect 176562 12248 176568 12300
rect 176620 12288 176626 12300
rect 320266 12288 320272 12300
rect 176620 12260 320272 12288
rect 176620 12248 176626 12260
rect 320266 12248 320272 12260
rect 320324 12248 320330 12300
rect 173802 12180 173808 12232
rect 173860 12220 173866 12232
rect 317598 12220 317604 12232
rect 173860 12192 317604 12220
rect 173860 12180 173866 12192
rect 317598 12180 317604 12192
rect 317656 12180 317662 12232
rect 169662 12112 169668 12164
rect 169720 12152 169726 12164
rect 316034 12152 316040 12164
rect 169720 12124 316040 12152
rect 169720 12112 169726 12124
rect 316034 12112 316040 12124
rect 316092 12112 316098 12164
rect 166902 12044 166908 12096
rect 166960 12084 166966 12096
rect 314746 12084 314752 12096
rect 166960 12056 314752 12084
rect 166960 12044 166966 12056
rect 314746 12044 314752 12056
rect 314804 12044 314810 12096
rect 162762 11976 162768 12028
rect 162820 12016 162826 12028
rect 313366 12016 313372 12028
rect 162820 11988 313372 12016
rect 162820 11976 162826 11988
rect 313366 11976 313372 11988
rect 313424 11976 313430 12028
rect 142062 11908 142068 11960
rect 142120 11948 142126 11960
rect 302418 11948 302424 11960
rect 142120 11920 302424 11948
rect 142120 11908 142126 11920
rect 302418 11908 302424 11920
rect 302476 11908 302482 11960
rect 416958 11908 416964 11960
rect 417016 11908 417022 11960
rect 126882 11840 126888 11892
rect 126940 11880 126946 11892
rect 293957 11883 294015 11889
rect 293957 11880 293969 11883
rect 126940 11852 293969 11880
rect 126940 11840 126946 11852
rect 293957 11849 293969 11852
rect 294003 11849 294015 11883
rect 293957 11843 294015 11849
rect 416976 11824 417004 11908
rect 128262 11772 128268 11824
rect 128320 11812 128326 11824
rect 295334 11812 295340 11824
rect 128320 11784 295340 11812
rect 128320 11772 128326 11784
rect 295334 11772 295340 11784
rect 295392 11772 295398 11824
rect 416958 11772 416964 11824
rect 417016 11772 417022 11824
rect 13630 11704 13636 11756
rect 13688 11744 13694 11756
rect 236178 11744 236184 11756
rect 13688 11716 236184 11744
rect 13688 11704 13694 11716
rect 236178 11704 236184 11716
rect 236236 11704 236242 11756
rect 252738 11744 252744 11756
rect 252699 11716 252744 11744
rect 252738 11704 252744 11716
rect 252796 11704 252802 11756
rect 187602 11636 187608 11688
rect 187660 11676 187666 11688
rect 325786 11676 325792 11688
rect 187660 11648 325792 11676
rect 187660 11636 187666 11648
rect 325786 11636 325792 11648
rect 325844 11636 325850 11688
rect 191742 11568 191748 11620
rect 191800 11608 191806 11620
rect 327258 11608 327264 11620
rect 191800 11580 327264 11608
rect 191800 11568 191806 11580
rect 327258 11568 327264 11580
rect 327316 11568 327322 11620
rect 194502 11500 194508 11552
rect 194560 11540 194566 11552
rect 328638 11540 328644 11552
rect 194560 11512 328644 11540
rect 194560 11500 194566 11512
rect 328638 11500 328644 11512
rect 328696 11500 328702 11552
rect 198642 11432 198648 11484
rect 198700 11472 198706 11484
rect 331214 11472 331220 11484
rect 198700 11444 331220 11472
rect 198700 11432 198706 11444
rect 331214 11432 331220 11444
rect 331272 11432 331278 11484
rect 201494 11364 201500 11416
rect 201552 11404 201558 11416
rect 332870 11404 332876 11416
rect 201552 11376 332876 11404
rect 201552 11364 201558 11376
rect 332870 11364 332876 11376
rect 332928 11364 332934 11416
rect 205542 11296 205548 11348
rect 205600 11336 205606 11348
rect 334345 11339 334403 11345
rect 334345 11336 334357 11339
rect 205600 11308 334357 11336
rect 205600 11296 205606 11308
rect 334345 11305 334357 11308
rect 334391 11305 334403 11339
rect 334345 11299 334403 11305
rect 143442 10956 143448 11008
rect 143500 10996 143506 11008
rect 302326 10996 302332 11008
rect 143500 10968 302332 10996
rect 143500 10956 143506 10968
rect 302326 10956 302332 10968
rect 302384 10956 302390 11008
rect 140682 10888 140688 10940
rect 140740 10928 140746 10940
rect 301038 10928 301044 10940
rect 140740 10900 301044 10928
rect 140740 10888 140746 10900
rect 301038 10888 301044 10900
rect 301096 10888 301102 10940
rect 124122 10820 124128 10872
rect 124180 10860 124186 10872
rect 292574 10860 292580 10872
rect 124180 10832 292580 10860
rect 124180 10820 124186 10832
rect 292574 10820 292580 10832
rect 292632 10820 292638 10872
rect 119982 10752 119988 10804
rect 120040 10792 120046 10804
rect 291194 10792 291200 10804
rect 120040 10764 291200 10792
rect 120040 10752 120046 10764
rect 291194 10752 291200 10764
rect 291252 10752 291258 10804
rect 117130 10684 117136 10736
rect 117188 10724 117194 10736
rect 288529 10727 288587 10733
rect 288529 10724 288541 10727
rect 117188 10696 288541 10724
rect 117188 10684 117194 10696
rect 288529 10693 288541 10696
rect 288575 10693 288587 10727
rect 288529 10687 288587 10693
rect 113082 10616 113088 10668
rect 113140 10656 113146 10668
rect 287054 10656 287060 10668
rect 113140 10628 287060 10656
rect 113140 10616 113146 10628
rect 287054 10616 287060 10628
rect 287112 10616 287118 10668
rect 289906 10616 289912 10668
rect 289964 10656 289970 10668
rect 367186 10656 367192 10668
rect 289964 10628 367192 10656
rect 289964 10616 289970 10628
rect 367186 10616 367192 10628
rect 367244 10616 367250 10668
rect 105170 10548 105176 10600
rect 105228 10588 105234 10600
rect 283006 10588 283012 10600
rect 105228 10560 283012 10588
rect 105228 10548 105234 10560
rect 283006 10548 283012 10560
rect 283064 10548 283070 10600
rect 289814 10548 289820 10600
rect 289872 10588 289878 10600
rect 367370 10588 367376 10600
rect 289872 10560 367376 10588
rect 289872 10548 289878 10560
rect 367370 10548 367376 10560
rect 367428 10548 367434 10600
rect 108758 10480 108764 10532
rect 108816 10520 108822 10532
rect 285674 10520 285680 10532
rect 108816 10492 285680 10520
rect 108816 10480 108822 10492
rect 285674 10480 285680 10492
rect 285732 10480 285738 10532
rect 287606 10480 287612 10532
rect 287664 10520 287670 10532
rect 365714 10520 365720 10532
rect 287664 10492 365720 10520
rect 287664 10480 287670 10492
rect 365714 10480 365720 10492
rect 365772 10480 365778 10532
rect 101582 10412 101588 10464
rect 101640 10452 101646 10464
rect 281534 10452 281540 10464
rect 101640 10424 281540 10452
rect 101640 10412 101646 10424
rect 281534 10412 281540 10424
rect 281592 10412 281598 10464
rect 299658 10412 299664 10464
rect 299716 10452 299722 10464
rect 379606 10452 379612 10464
rect 299716 10424 379612 10452
rect 299716 10412 299722 10424
rect 379606 10412 379612 10424
rect 379664 10412 379670 10464
rect 99190 10344 99196 10396
rect 99248 10384 99254 10396
rect 280154 10384 280160 10396
rect 99248 10356 280160 10384
rect 99248 10344 99254 10356
rect 280154 10344 280160 10356
rect 280212 10344 280218 10396
rect 300946 10344 300952 10396
rect 301004 10384 301010 10396
rect 383746 10384 383752 10396
rect 301004 10356 383752 10384
rect 301004 10344 301010 10356
rect 383746 10344 383752 10356
rect 383804 10344 383810 10396
rect 64782 10276 64788 10328
rect 64840 10316 64846 10328
rect 262306 10316 262312 10328
rect 64840 10288 262312 10316
rect 64840 10276 64846 10288
rect 262306 10276 262312 10288
rect 262364 10276 262370 10328
rect 292942 10276 292948 10328
rect 293000 10316 293006 10328
rect 378318 10316 378324 10328
rect 293000 10288 378324 10316
rect 293000 10276 293006 10288
rect 378318 10276 378324 10288
rect 378376 10276 378382 10328
rect 147582 10208 147588 10260
rect 147640 10248 147646 10260
rect 304994 10248 305000 10260
rect 147640 10220 305000 10248
rect 147640 10208 147646 10220
rect 304994 10208 305000 10220
rect 305052 10208 305058 10260
rect 151630 10140 151636 10192
rect 151688 10180 151694 10192
rect 306374 10180 306380 10192
rect 151688 10152 306380 10180
rect 151688 10140 151694 10152
rect 306374 10140 306380 10152
rect 306432 10140 306438 10192
rect 154482 10072 154488 10124
rect 154540 10112 154546 10124
rect 308033 10115 308091 10121
rect 308033 10112 308045 10115
rect 154540 10084 308045 10112
rect 154540 10072 154546 10084
rect 308033 10081 308045 10084
rect 308079 10081 308091 10115
rect 308033 10075 308091 10081
rect 158622 10004 158628 10056
rect 158680 10044 158686 10056
rect 310514 10044 310520 10056
rect 158680 10016 310520 10044
rect 158680 10004 158686 10016
rect 310514 10004 310520 10016
rect 310572 10004 310578 10056
rect 161382 9936 161388 9988
rect 161440 9976 161446 9988
rect 311894 9976 311900 9988
rect 161440 9948 311900 9976
rect 161440 9936 161446 9948
rect 311894 9936 311900 9948
rect 311952 9936 311958 9988
rect 376849 9979 376907 9985
rect 376849 9945 376861 9979
rect 376895 9976 376907 9979
rect 377030 9976 377036 9988
rect 376895 9948 377036 9976
rect 376895 9945 376907 9948
rect 376849 9939 376907 9945
rect 377030 9936 377036 9948
rect 377088 9936 377094 9988
rect 246758 9868 246764 9920
rect 246816 9908 246822 9920
rect 356238 9908 356244 9920
rect 246816 9880 356244 9908
rect 246816 9868 246822 9880
rect 356238 9868 356244 9880
rect 356296 9868 356302 9920
rect 250346 9800 250352 9852
rect 250404 9840 250410 9852
rect 357529 9843 357587 9849
rect 357529 9840 357541 9843
rect 250404 9812 357541 9840
rect 250404 9800 250410 9812
rect 357529 9809 357541 9812
rect 357575 9809 357587 9843
rect 357529 9803 357587 9809
rect 253842 9732 253848 9784
rect 253900 9772 253906 9784
rect 360286 9772 360292 9784
rect 253900 9744 360292 9772
rect 253900 9732 253906 9744
rect 360286 9732 360292 9744
rect 360344 9732 360350 9784
rect 249978 9664 249984 9716
rect 250036 9704 250042 9716
rect 250070 9704 250076 9716
rect 250036 9676 250076 9704
rect 250036 9664 250042 9676
rect 250070 9664 250076 9676
rect 250128 9664 250134 9716
rect 254026 9664 254032 9716
rect 254084 9704 254090 9716
rect 254302 9704 254308 9716
rect 254084 9676 254308 9704
rect 254084 9664 254090 9676
rect 254302 9664 254308 9676
rect 254360 9664 254366 9716
rect 255314 9664 255320 9716
rect 255372 9704 255378 9716
rect 255590 9704 255596 9716
rect 255372 9676 255596 9704
rect 255372 9664 255378 9676
rect 255590 9664 255596 9676
rect 255648 9664 255654 9716
rect 257430 9664 257436 9716
rect 257488 9704 257494 9716
rect 361758 9704 361764 9716
rect 257488 9676 361764 9704
rect 257488 9664 257494 9676
rect 361758 9664 361764 9676
rect 361816 9664 361822 9716
rect 375466 9664 375472 9716
rect 375524 9704 375530 9716
rect 375742 9704 375748 9716
rect 375524 9676 375748 9704
rect 375524 9664 375530 9676
rect 375742 9664 375748 9676
rect 375800 9664 375806 9716
rect 397546 9704 397552 9716
rect 397507 9676 397552 9704
rect 397546 9664 397552 9676
rect 397604 9664 397610 9716
rect 407761 9707 407819 9713
rect 407761 9673 407773 9707
rect 407807 9704 407819 9707
rect 407850 9704 407856 9716
rect 407807 9676 407856 9704
rect 407807 9673 407819 9676
rect 407761 9667 407819 9673
rect 407850 9664 407856 9676
rect 407908 9664 407914 9716
rect 422110 9664 422116 9716
rect 422168 9704 422174 9716
rect 422386 9704 422392 9716
rect 422168 9676 422392 9704
rect 422168 9664 422174 9676
rect 422386 9664 422392 9676
rect 422444 9664 422450 9716
rect 427817 9707 427875 9713
rect 427817 9673 427829 9707
rect 427863 9704 427875 9707
rect 427906 9704 427912 9716
rect 427863 9676 427912 9704
rect 427863 9673 427875 9676
rect 427817 9667 427875 9673
rect 427906 9664 427912 9676
rect 427964 9664 427970 9716
rect 203886 9596 203892 9648
rect 203944 9636 203950 9648
rect 333974 9636 333980 9648
rect 203944 9608 333980 9636
rect 203944 9596 203950 9608
rect 333974 9596 333980 9608
rect 334032 9596 334038 9648
rect 346486 9636 346492 9648
rect 346447 9608 346492 9636
rect 346486 9596 346492 9608
rect 346544 9596 346550 9648
rect 369946 9636 369952 9648
rect 369907 9608 369952 9636
rect 369946 9596 369952 9608
rect 370004 9596 370010 9648
rect 371234 9636 371240 9648
rect 371195 9608 371240 9636
rect 371234 9596 371240 9608
rect 371292 9596 371298 9648
rect 393038 9636 393044 9648
rect 392999 9608 393044 9636
rect 393038 9596 393044 9608
rect 393096 9596 393102 9648
rect 200390 9528 200396 9580
rect 200448 9568 200454 9580
rect 332594 9568 332600 9580
rect 200448 9540 332600 9568
rect 200448 9528 200454 9540
rect 332594 9528 332600 9540
rect 332652 9528 332658 9580
rect 196802 9460 196808 9512
rect 196860 9500 196866 9512
rect 330113 9503 330171 9509
rect 330113 9500 330125 9503
rect 196860 9472 330125 9500
rect 196860 9460 196866 9472
rect 330113 9469 330125 9472
rect 330159 9469 330171 9503
rect 330113 9463 330171 9469
rect 193214 9392 193220 9444
rect 193272 9432 193278 9444
rect 328730 9432 328736 9444
rect 193272 9404 328736 9432
rect 193272 9392 193278 9404
rect 328730 9392 328736 9404
rect 328788 9392 328794 9444
rect 189626 9324 189632 9376
rect 189684 9364 189690 9376
rect 327074 9364 327080 9376
rect 189684 9336 327080 9364
rect 189684 9324 189690 9336
rect 327074 9324 327080 9336
rect 327132 9324 327138 9376
rect 186038 9256 186044 9308
rect 186096 9296 186102 9308
rect 324406 9296 324412 9308
rect 186096 9268 324412 9296
rect 186096 9256 186102 9268
rect 324406 9256 324412 9268
rect 324464 9256 324470 9308
rect 361666 9296 361672 9308
rect 325344 9268 361672 9296
rect 182542 9188 182548 9240
rect 182600 9228 182606 9240
rect 323210 9228 323216 9240
rect 182600 9200 323216 9228
rect 182600 9188 182606 9200
rect 323210 9188 323216 9200
rect 323268 9188 323274 9240
rect 178954 9120 178960 9172
rect 179012 9160 179018 9172
rect 321554 9160 321560 9172
rect 179012 9132 321560 9160
rect 179012 9120 179018 9132
rect 321554 9120 321560 9132
rect 321612 9120 321618 9172
rect 322566 9120 322572 9172
rect 322624 9160 322630 9172
rect 325344 9160 325372 9268
rect 361666 9256 361672 9268
rect 361724 9256 361730 9308
rect 327074 9188 327080 9240
rect 327132 9228 327138 9240
rect 392026 9228 392032 9240
rect 327132 9200 392032 9228
rect 327132 9188 327138 9200
rect 392026 9188 392032 9200
rect 392084 9188 392090 9240
rect 322624 9132 325372 9160
rect 322624 9120 322630 9132
rect 325510 9120 325516 9172
rect 325568 9160 325574 9172
rect 390646 9160 390652 9172
rect 325568 9132 390652 9160
rect 325568 9120 325574 9132
rect 390646 9120 390652 9132
rect 390704 9120 390710 9172
rect 175366 9052 175372 9104
rect 175424 9092 175430 9104
rect 319070 9092 319076 9104
rect 175424 9064 319076 9092
rect 175424 9052 175430 9064
rect 319070 9052 319076 9064
rect 319128 9052 319134 9104
rect 328546 9052 328552 9104
rect 328604 9092 328610 9104
rect 394786 9092 394792 9104
rect 328604 9064 394792 9092
rect 328604 9052 328610 9064
rect 394786 9052 394792 9064
rect 394844 9052 394850 9104
rect 171778 8984 171784 9036
rect 171836 9024 171842 9036
rect 317690 9024 317696 9036
rect 171836 8996 317696 9024
rect 171836 8984 171842 8996
rect 317690 8984 317696 8996
rect 317748 8984 317754 9036
rect 323578 8984 323584 9036
rect 323636 9024 323642 9036
rect 389266 9024 389272 9036
rect 323636 8996 389272 9024
rect 323636 8984 323642 8996
rect 389266 8984 389272 8996
rect 389324 8984 389330 9036
rect 132586 8916 132592 8968
rect 132644 8956 132650 8968
rect 296806 8956 296812 8968
rect 132644 8928 296812 8956
rect 132644 8916 132650 8928
rect 296806 8916 296812 8928
rect 296864 8916 296870 8968
rect 334710 8916 334716 8968
rect 334768 8956 334774 8968
rect 401686 8956 401692 8968
rect 334768 8928 401692 8956
rect 334768 8916 334774 8928
rect 401686 8916 401692 8928
rect 401744 8916 401750 8968
rect 210970 8848 210976 8900
rect 211028 8888 211034 8900
rect 338206 8888 338212 8900
rect 211028 8860 338212 8888
rect 211028 8848 211034 8860
rect 338206 8848 338212 8860
rect 338264 8848 338270 8900
rect 207474 8780 207480 8832
rect 207532 8820 207538 8832
rect 335354 8820 335360 8832
rect 207532 8792 335360 8820
rect 207532 8780 207538 8792
rect 335354 8780 335360 8792
rect 335412 8780 335418 8832
rect 214650 8712 214656 8764
rect 214708 8752 214714 8764
rect 339770 8752 339776 8764
rect 214708 8724 339776 8752
rect 214708 8712 214714 8724
rect 339770 8712 339776 8724
rect 339828 8712 339834 8764
rect 221734 8644 221740 8696
rect 221792 8684 221798 8696
rect 343726 8684 343732 8696
rect 221792 8656 343732 8684
rect 221792 8644 221798 8656
rect 343726 8644 343732 8656
rect 343784 8644 343790 8696
rect 218146 8576 218152 8628
rect 218204 8616 218210 8628
rect 340874 8616 340880 8628
rect 218204 8588 340880 8616
rect 218204 8576 218210 8588
rect 340874 8576 340880 8588
rect 340932 8576 340938 8628
rect 225322 8508 225328 8560
rect 225380 8548 225386 8560
rect 345198 8548 345204 8560
rect 225380 8520 345204 8548
rect 225380 8508 225386 8520
rect 345198 8508 345204 8520
rect 345256 8508 345262 8560
rect 228910 8440 228916 8492
rect 228968 8480 228974 8492
rect 346489 8483 346547 8489
rect 346489 8480 346501 8483
rect 228968 8452 346501 8480
rect 228968 8440 228974 8452
rect 346489 8449 346501 8452
rect 346535 8449 346547 8483
rect 346489 8443 346547 8449
rect 232498 8372 232504 8424
rect 232556 8412 232562 8424
rect 349246 8412 349252 8424
rect 232556 8384 349252 8412
rect 232556 8372 232562 8384
rect 349246 8372 349252 8384
rect 349304 8372 349310 8424
rect 235994 8304 236000 8356
rect 236052 8344 236058 8356
rect 350718 8344 350724 8356
rect 236052 8316 350724 8344
rect 236052 8304 236058 8316
rect 350718 8304 350724 8316
rect 350776 8304 350782 8356
rect 358906 8304 358912 8356
rect 358964 8344 358970 8356
rect 358998 8344 359004 8356
rect 358964 8316 359004 8344
rect 358964 8304 358970 8316
rect 358998 8304 359004 8316
rect 359056 8304 359062 8356
rect 364426 8304 364432 8356
rect 364484 8344 364490 8356
rect 364794 8344 364800 8356
rect 364484 8316 364800 8344
rect 364484 8304 364490 8316
rect 364794 8304 364800 8316
rect 364852 8304 364858 8356
rect 56410 8236 56416 8288
rect 56468 8276 56474 8288
rect 258350 8276 258356 8288
rect 56468 8248 258356 8276
rect 56468 8236 56474 8248
rect 258350 8236 258356 8248
rect 258408 8236 258414 8288
rect 274082 8236 274088 8288
rect 274140 8276 274146 8288
rect 369949 8279 370007 8285
rect 369949 8276 369961 8279
rect 274140 8248 369961 8276
rect 274140 8236 274146 8248
rect 369949 8245 369961 8248
rect 369995 8245 370007 8279
rect 369949 8239 370007 8245
rect 52822 8168 52828 8220
rect 52880 8208 52886 8220
rect 256786 8208 256792 8220
rect 52880 8180 256792 8208
rect 52880 8168 52886 8180
rect 256786 8168 256792 8180
rect 256844 8168 256850 8220
rect 270494 8168 270500 8220
rect 270552 8208 270558 8220
rect 368566 8208 368572 8220
rect 270552 8180 368572 8208
rect 270552 8168 270558 8180
rect 368566 8168 368572 8180
rect 368624 8168 368630 8220
rect 49326 8100 49332 8152
rect 49384 8140 49390 8152
rect 254026 8140 254032 8152
rect 49384 8112 254032 8140
rect 49384 8100 49390 8112
rect 254026 8100 254032 8112
rect 254084 8100 254090 8152
rect 266998 8100 267004 8152
rect 267056 8140 267062 8152
rect 367094 8140 367100 8152
rect 267056 8112 367100 8140
rect 267056 8100 267062 8112
rect 367094 8100 367100 8112
rect 367152 8100 367158 8152
rect 44542 8032 44548 8084
rect 44600 8072 44606 8084
rect 252646 8072 252652 8084
rect 44600 8044 252652 8072
rect 44600 8032 44606 8044
rect 252646 8032 252652 8044
rect 252704 8032 252710 8084
rect 263410 8032 263416 8084
rect 263468 8072 263474 8084
rect 364426 8072 364432 8084
rect 263468 8044 364432 8072
rect 263468 8032 263474 8044
rect 364426 8032 364432 8044
rect 364484 8032 364490 8084
rect 40954 7964 40960 8016
rect 41012 8004 41018 8016
rect 249978 8004 249984 8016
rect 41012 7976 249984 8004
rect 41012 7964 41018 7976
rect 249978 7964 249984 7976
rect 250036 7964 250042 8016
rect 259822 7964 259828 8016
rect 259880 8004 259886 8016
rect 363046 8004 363052 8016
rect 259880 7976 363052 8004
rect 259880 7964 259886 7976
rect 363046 7964 363052 7976
rect 363104 7964 363110 8016
rect 37366 7896 37372 7948
rect 37424 7936 37430 7948
rect 248506 7936 248512 7948
rect 37424 7908 248512 7936
rect 37424 7896 37430 7908
rect 248506 7896 248512 7908
rect 248564 7896 248570 7948
rect 256234 7896 256240 7948
rect 256292 7936 256298 7948
rect 361574 7936 361580 7948
rect 256292 7908 361580 7936
rect 256292 7896 256298 7908
rect 361574 7896 361580 7908
rect 361632 7896 361638 7948
rect 33870 7828 33876 7880
rect 33928 7868 33934 7880
rect 247218 7868 247224 7880
rect 33928 7840 247224 7868
rect 33928 7828 33934 7840
rect 247218 7828 247224 7840
rect 247276 7828 247282 7880
rect 252646 7828 252652 7880
rect 252704 7868 252710 7880
rect 358906 7868 358912 7880
rect 252704 7840 358912 7868
rect 252704 7828 252710 7840
rect 358906 7828 358912 7840
rect 358964 7828 358970 7880
rect 30282 7760 30288 7812
rect 30340 7800 30346 7812
rect 244274 7800 244280 7812
rect 30340 7772 244280 7800
rect 30340 7760 30346 7772
rect 244274 7760 244280 7772
rect 244332 7760 244338 7812
rect 249150 7760 249156 7812
rect 249208 7800 249214 7812
rect 357434 7800 357440 7812
rect 249208 7772 357440 7800
rect 249208 7760 249214 7772
rect 357434 7760 357440 7772
rect 357492 7760 357498 7812
rect 26694 7692 26700 7744
rect 26752 7732 26758 7744
rect 242894 7732 242900 7744
rect 26752 7704 242900 7732
rect 26752 7692 26758 7704
rect 242894 7692 242900 7704
rect 242952 7692 242958 7744
rect 245562 7692 245568 7744
rect 245620 7732 245626 7744
rect 356146 7732 356152 7744
rect 245620 7704 356152 7732
rect 245620 7692 245626 7704
rect 356146 7692 356152 7704
rect 356204 7692 356210 7744
rect 8846 7624 8852 7676
rect 8904 7664 8910 7676
rect 233326 7664 233332 7676
rect 8904 7636 233332 7664
rect 8904 7624 8910 7636
rect 233326 7624 233332 7636
rect 233384 7624 233390 7676
rect 234798 7624 234804 7676
rect 234856 7664 234862 7676
rect 350626 7664 350632 7676
rect 234856 7636 350632 7664
rect 234856 7624 234862 7636
rect 350626 7624 350632 7636
rect 350684 7624 350690 7676
rect 4062 7556 4068 7608
rect 4120 7596 4126 7608
rect 230658 7596 230664 7608
rect 4120 7568 230664 7596
rect 4120 7556 4126 7568
rect 230658 7556 230664 7568
rect 230716 7556 230722 7608
rect 231302 7556 231308 7608
rect 231360 7596 231366 7608
rect 347866 7596 347872 7608
rect 231360 7568 347872 7596
rect 231360 7556 231366 7568
rect 347866 7556 347872 7568
rect 347924 7556 347930 7608
rect 351822 7556 351828 7608
rect 351880 7596 351886 7608
rect 405826 7596 405832 7608
rect 351880 7568 405832 7596
rect 351880 7556 351886 7568
rect 405826 7556 405832 7568
rect 405884 7556 405890 7608
rect 477586 7556 477592 7608
rect 477644 7596 477650 7608
rect 478690 7596 478696 7608
rect 477644 7568 478696 7596
rect 477644 7556 477650 7568
rect 478690 7556 478696 7568
rect 478748 7556 478754 7608
rect 87322 7488 87328 7540
rect 87380 7528 87386 7540
rect 274634 7528 274640 7540
rect 87380 7500 274640 7528
rect 87380 7488 87386 7500
rect 274634 7488 274640 7500
rect 274692 7488 274698 7540
rect 277670 7488 277676 7540
rect 277728 7528 277734 7540
rect 372706 7528 372712 7540
rect 277728 7500 372712 7528
rect 277728 7488 277734 7500
rect 372706 7488 372712 7500
rect 372764 7488 372770 7540
rect 90910 7420 90916 7472
rect 90968 7460 90974 7472
rect 276014 7460 276020 7472
rect 90968 7432 276020 7460
rect 90968 7420 90974 7432
rect 276014 7420 276020 7432
rect 276072 7420 276078 7472
rect 281258 7420 281264 7472
rect 281316 7460 281322 7472
rect 374086 7460 374092 7472
rect 281316 7432 374092 7460
rect 281316 7420 281322 7432
rect 374086 7420 374092 7432
rect 374144 7420 374150 7472
rect 94498 7352 94504 7404
rect 94556 7392 94562 7404
rect 277486 7392 277492 7404
rect 94556 7364 277492 7392
rect 94556 7352 94562 7364
rect 277486 7352 277492 7364
rect 277544 7352 277550 7404
rect 284754 7352 284760 7404
rect 284812 7392 284818 7404
rect 375466 7392 375472 7404
rect 284812 7364 375472 7392
rect 284812 7352 284818 7364
rect 375466 7352 375472 7364
rect 375524 7352 375530 7404
rect 138474 7284 138480 7336
rect 138532 7324 138538 7336
rect 300854 7324 300860 7336
rect 138532 7296 300860 7324
rect 138532 7284 138538 7296
rect 300854 7284 300860 7296
rect 300912 7284 300918 7336
rect 347958 7284 347964 7336
rect 348016 7324 348022 7336
rect 397546 7324 397552 7336
rect 348016 7296 397552 7324
rect 348016 7284 348022 7296
rect 397546 7284 397552 7296
rect 397604 7284 397610 7336
rect 141970 7216 141976 7268
rect 142028 7256 142034 7268
rect 302510 7256 302516 7268
rect 142028 7228 302516 7256
rect 142028 7216 142034 7228
rect 302510 7216 302516 7228
rect 302568 7216 302574 7268
rect 346486 7216 346492 7268
rect 346544 7256 346550 7268
rect 396166 7256 396172 7268
rect 346544 7228 396172 7256
rect 346544 7216 346550 7228
rect 396166 7216 396172 7228
rect 396224 7216 396230 7268
rect 224126 7148 224132 7200
rect 224184 7188 224190 7200
rect 345106 7188 345112 7200
rect 224184 7160 345112 7188
rect 224184 7148 224190 7160
rect 345106 7148 345112 7160
rect 345164 7148 345170 7200
rect 227714 7080 227720 7132
rect 227772 7120 227778 7132
rect 346394 7120 346400 7132
rect 227772 7092 346400 7120
rect 227772 7080 227778 7092
rect 346394 7080 346400 7092
rect 346452 7080 346458 7132
rect 238386 7012 238392 7064
rect 238444 7052 238450 7064
rect 351914 7052 351920 7064
rect 238444 7024 351920 7052
rect 238444 7012 238450 7024
rect 351914 7012 351920 7024
rect 351972 7012 351978 7064
rect 241974 6944 241980 6996
rect 242032 6984 242038 6996
rect 353386 6984 353392 6996
rect 242032 6956 353392 6984
rect 242032 6944 242038 6956
rect 353386 6944 353392 6956
rect 353444 6944 353450 6996
rect 163498 6808 163504 6860
rect 163556 6848 163562 6860
rect 313550 6848 313556 6860
rect 163556 6820 313556 6848
rect 163556 6808 163562 6820
rect 313550 6808 313556 6820
rect 313608 6808 313614 6860
rect 349062 6808 349068 6860
rect 349120 6848 349126 6860
rect 408770 6848 408776 6860
rect 349120 6820 408776 6848
rect 349120 6808 349126 6820
rect 408770 6808 408776 6820
rect 408828 6808 408834 6860
rect 83826 6740 83832 6792
rect 83884 6780 83890 6792
rect 271874 6780 271880 6792
rect 83884 6752 271880 6780
rect 83884 6740 83890 6752
rect 271874 6740 271880 6752
rect 271932 6740 271938 6792
rect 315209 6783 315267 6789
rect 315209 6749 315221 6783
rect 315255 6780 315267 6783
rect 320174 6780 320180 6792
rect 315255 6752 320180 6780
rect 315255 6749 315267 6752
rect 315209 6743 315267 6749
rect 320174 6740 320180 6752
rect 320232 6740 320238 6792
rect 325602 6740 325608 6792
rect 325660 6780 325666 6792
rect 386506 6780 386512 6792
rect 325660 6752 386512 6780
rect 325660 6740 325666 6752
rect 386506 6740 386512 6752
rect 386564 6740 386570 6792
rect 80238 6672 80244 6724
rect 80296 6712 80302 6724
rect 270586 6712 270592 6724
rect 80296 6684 270592 6712
rect 80296 6672 80302 6684
rect 270586 6672 270592 6684
rect 270644 6672 270650 6724
rect 318794 6672 318800 6724
rect 318852 6712 318858 6724
rect 380802 6712 380808 6724
rect 318852 6684 380808 6712
rect 318852 6672 318858 6684
rect 380802 6672 380808 6684
rect 380860 6672 380866 6724
rect 76650 6604 76656 6656
rect 76708 6644 76714 6656
rect 269114 6644 269120 6656
rect 76708 6616 269120 6644
rect 76708 6604 76714 6616
rect 269114 6604 269120 6616
rect 269172 6604 269178 6656
rect 320174 6604 320180 6656
rect 320232 6644 320238 6656
rect 385126 6644 385132 6656
rect 320232 6616 385132 6644
rect 320232 6604 320238 6616
rect 385126 6604 385132 6616
rect 385184 6604 385190 6656
rect 73062 6536 73068 6588
rect 73120 6576 73126 6588
rect 266354 6576 266360 6588
rect 73120 6548 266360 6576
rect 73120 6536 73126 6548
rect 266354 6536 266360 6548
rect 266412 6536 266418 6588
rect 312170 6536 312176 6588
rect 312228 6576 312234 6588
rect 389358 6576 389364 6588
rect 312228 6548 389364 6576
rect 312228 6536 312234 6548
rect 389358 6536 389364 6548
rect 389416 6536 389422 6588
rect 69474 6468 69480 6520
rect 69532 6508 69538 6520
rect 264974 6508 264980 6520
rect 69532 6480 264980 6508
rect 69532 6468 69538 6480
rect 264974 6468 264980 6480
rect 265032 6468 265038 6520
rect 308582 6468 308588 6520
rect 308640 6508 308646 6520
rect 387886 6508 387892 6520
rect 308640 6480 387892 6508
rect 308640 6468 308646 6480
rect 387886 6468 387892 6480
rect 387944 6468 387950 6520
rect 62390 6400 62396 6452
rect 62448 6440 62454 6452
rect 260926 6440 260932 6452
rect 62448 6412 260932 6440
rect 62448 6400 62454 6412
rect 260926 6400 260932 6412
rect 260984 6400 260990 6452
rect 304994 6400 305000 6452
rect 305052 6440 305058 6452
rect 386414 6440 386420 6452
rect 305052 6412 386420 6440
rect 305052 6400 305058 6412
rect 386414 6400 386420 6412
rect 386472 6400 386478 6452
rect 65978 6332 65984 6384
rect 66036 6372 66042 6384
rect 263686 6372 263692 6384
rect 66036 6344 263692 6372
rect 66036 6332 66042 6344
rect 263686 6332 263692 6344
rect 263744 6332 263750 6384
rect 290734 6332 290740 6384
rect 290792 6372 290798 6384
rect 378226 6372 378232 6384
rect 290792 6344 378232 6372
rect 290792 6332 290798 6344
rect 378226 6332 378232 6344
rect 378284 6332 378290 6384
rect 58802 6264 58808 6316
rect 58860 6304 58866 6316
rect 259454 6304 259460 6316
rect 58860 6276 259460 6304
rect 58860 6264 58866 6276
rect 259454 6264 259460 6276
rect 259512 6264 259518 6316
rect 287146 6264 287152 6316
rect 287204 6304 287210 6316
rect 376849 6307 376907 6313
rect 376849 6304 376861 6307
rect 287204 6276 376861 6304
rect 287204 6264 287210 6276
rect 376849 6273 376861 6276
rect 376895 6273 376907 6307
rect 376849 6267 376907 6273
rect 55214 6196 55220 6248
rect 55272 6236 55278 6248
rect 258258 6236 258264 6248
rect 55272 6208 258264 6236
rect 55272 6196 55278 6208
rect 258258 6196 258264 6208
rect 258316 6196 258322 6248
rect 283650 6196 283656 6248
rect 283708 6236 283714 6248
rect 375374 6236 375380 6248
rect 283708 6208 375380 6236
rect 283708 6196 283714 6208
rect 375374 6196 375380 6208
rect 375432 6196 375438 6248
rect 379974 6196 379980 6248
rect 380032 6236 380038 6248
rect 425146 6236 425152 6248
rect 380032 6208 425152 6236
rect 380032 6196 380038 6208
rect 425146 6196 425152 6208
rect 425204 6196 425210 6248
rect 51626 6128 51632 6180
rect 51684 6168 51690 6180
rect 255314 6168 255320 6180
rect 51684 6140 255320 6168
rect 51684 6128 51690 6140
rect 255314 6128 255320 6140
rect 255372 6128 255378 6180
rect 279970 6128 279976 6180
rect 280028 6168 280034 6180
rect 372798 6168 372804 6180
rect 280028 6140 372804 6168
rect 280028 6128 280034 6140
rect 372798 6128 372804 6140
rect 372856 6128 372862 6180
rect 372890 6128 372896 6180
rect 372948 6168 372954 6180
rect 421098 6168 421104 6180
rect 372948 6140 421104 6168
rect 372948 6128 372954 6140
rect 421098 6128 421104 6140
rect 421156 6128 421162 6180
rect 167086 6060 167092 6112
rect 167144 6100 167150 6112
rect 314562 6100 314568 6112
rect 167144 6072 314568 6100
rect 167144 6060 167150 6072
rect 314562 6060 314568 6072
rect 314620 6060 314626 6112
rect 314654 6060 314660 6112
rect 314712 6100 314718 6112
rect 371237 6103 371295 6109
rect 371237 6100 371249 6103
rect 314712 6072 371249 6100
rect 314712 6060 314718 6072
rect 371237 6069 371249 6072
rect 371283 6069 371295 6103
rect 371237 6063 371295 6069
rect 170582 5992 170588 6044
rect 170640 6032 170646 6044
rect 317414 6032 317420 6044
rect 170640 6004 317420 6032
rect 170640 5992 170646 6004
rect 317414 5992 317420 6004
rect 317472 5992 317478 6044
rect 322201 6035 322259 6041
rect 322201 6001 322213 6035
rect 322247 6032 322259 6035
rect 322934 6032 322940 6044
rect 322247 6004 322940 6032
rect 322247 6001 322259 6004
rect 322201 5995 322259 6001
rect 322934 5992 322940 6004
rect 322992 5992 322998 6044
rect 354950 5992 354956 6044
rect 355008 6032 355014 6044
rect 411346 6032 411352 6044
rect 355008 6004 411352 6032
rect 355008 5992 355014 6004
rect 411346 5992 411352 6004
rect 411404 5992 411410 6044
rect 174170 5924 174176 5976
rect 174228 5964 174234 5976
rect 174228 5936 315344 5964
rect 174228 5924 174234 5936
rect 177758 5856 177764 5908
rect 177816 5896 177822 5908
rect 315209 5899 315267 5905
rect 315209 5896 315221 5899
rect 177816 5868 315221 5896
rect 177816 5856 177822 5868
rect 315209 5865 315221 5868
rect 315255 5865 315267 5899
rect 315316 5896 315344 5936
rect 316586 5924 316592 5976
rect 316644 5964 316650 5976
rect 369854 5964 369860 5976
rect 316644 5936 369860 5964
rect 316644 5924 316650 5936
rect 369854 5924 369860 5936
rect 369912 5924 369918 5976
rect 318886 5896 318892 5908
rect 315316 5868 318892 5896
rect 315209 5859 315267 5865
rect 318886 5856 318892 5868
rect 318944 5856 318950 5908
rect 325326 5856 325332 5908
rect 325384 5896 325390 5908
rect 360194 5896 360200 5908
rect 325384 5868 360200 5896
rect 325384 5856 325390 5868
rect 360194 5856 360200 5868
rect 360252 5856 360258 5908
rect 362126 5856 362132 5908
rect 362184 5896 362190 5908
rect 415578 5896 415584 5908
rect 362184 5868 415584 5896
rect 362184 5856 362190 5868
rect 415578 5856 415584 5868
rect 415636 5856 415642 5908
rect 181346 5788 181352 5840
rect 181404 5828 181410 5840
rect 322201 5831 322259 5837
rect 322201 5828 322213 5831
rect 181404 5800 322213 5828
rect 181404 5788 181410 5800
rect 322201 5797 322213 5800
rect 322247 5797 322259 5831
rect 322201 5791 322259 5797
rect 322658 5788 322664 5840
rect 322716 5828 322722 5840
rect 364334 5828 364340 5840
rect 322716 5800 364340 5828
rect 322716 5788 322722 5800
rect 364334 5788 364340 5800
rect 364392 5788 364398 5840
rect 369210 5788 369216 5840
rect 369268 5828 369274 5840
rect 419626 5828 419632 5840
rect 369268 5800 419632 5828
rect 369268 5788 369274 5800
rect 419626 5788 419632 5800
rect 419684 5788 419690 5840
rect 184842 5720 184848 5772
rect 184900 5760 184906 5772
rect 324314 5760 324320 5772
rect 184900 5732 324320 5760
rect 184900 5720 184906 5732
rect 324314 5720 324320 5732
rect 324372 5720 324378 5772
rect 188430 5652 188436 5704
rect 188488 5692 188494 5704
rect 325694 5692 325700 5704
rect 188488 5664 325700 5692
rect 188488 5652 188494 5664
rect 325694 5652 325700 5664
rect 325752 5652 325758 5704
rect 192018 5584 192024 5636
rect 192076 5624 192082 5636
rect 328454 5624 328460 5636
rect 192076 5596 328460 5624
rect 192076 5584 192082 5596
rect 328454 5584 328460 5596
rect 328512 5584 328518 5636
rect 195606 5516 195612 5568
rect 195664 5556 195670 5568
rect 329834 5556 329840 5568
rect 195664 5528 329840 5556
rect 195664 5516 195670 5528
rect 329834 5516 329840 5528
rect 329892 5516 329898 5568
rect 137278 5448 137284 5500
rect 137336 5488 137342 5500
rect 299474 5488 299480 5500
rect 137336 5460 299480 5488
rect 137336 5448 137342 5460
rect 299474 5448 299480 5460
rect 299532 5448 299538 5500
rect 315758 5448 315764 5500
rect 315816 5488 315822 5500
rect 391934 5488 391940 5500
rect 315816 5460 391940 5488
rect 315816 5448 315822 5460
rect 391934 5448 391940 5460
rect 391992 5448 391998 5500
rect 401318 5448 401324 5500
rect 401376 5488 401382 5500
rect 436186 5488 436192 5500
rect 401376 5460 436192 5488
rect 401376 5448 401382 5460
rect 436186 5448 436192 5460
rect 436244 5448 436250 5500
rect 133782 5380 133788 5432
rect 133840 5420 133846 5432
rect 298094 5420 298100 5432
rect 133840 5392 298100 5420
rect 133840 5380 133846 5392
rect 298094 5380 298100 5392
rect 298152 5380 298158 5432
rect 301406 5380 301412 5432
rect 301464 5420 301470 5432
rect 383838 5420 383844 5432
rect 301464 5392 383844 5420
rect 301464 5380 301470 5392
rect 383838 5380 383844 5392
rect 383896 5380 383902 5432
rect 397822 5380 397828 5432
rect 397880 5420 397886 5432
rect 433610 5420 433616 5432
rect 397880 5392 433616 5420
rect 397880 5380 397886 5392
rect 433610 5380 433616 5392
rect 433668 5380 433674 5432
rect 130194 5312 130200 5364
rect 130252 5352 130258 5364
rect 296714 5352 296720 5364
rect 130252 5324 296720 5352
rect 130252 5312 130258 5324
rect 296714 5312 296720 5324
rect 296772 5312 296778 5364
rect 297910 5312 297916 5364
rect 297968 5352 297974 5364
rect 382369 5355 382427 5361
rect 382369 5352 382381 5355
rect 297968 5324 382381 5352
rect 297968 5312 297974 5324
rect 382369 5321 382381 5324
rect 382415 5321 382427 5355
rect 382369 5315 382427 5321
rect 394234 5312 394240 5364
rect 394292 5352 394298 5364
rect 432138 5352 432144 5364
rect 394292 5324 432144 5352
rect 394292 5312 394298 5324
rect 432138 5312 432144 5324
rect 432196 5312 432202 5364
rect 67174 5244 67180 5296
rect 67232 5284 67238 5296
rect 263778 5284 263784 5296
rect 67232 5256 263784 5284
rect 67232 5244 67238 5256
rect 263778 5244 263784 5256
rect 263836 5244 263842 5296
rect 294322 5244 294328 5296
rect 294380 5284 294386 5296
rect 380894 5284 380900 5296
rect 294380 5256 380900 5284
rect 294380 5244 294386 5256
rect 380894 5244 380900 5256
rect 380952 5244 380958 5296
rect 390646 5244 390652 5296
rect 390704 5284 390710 5296
rect 430666 5284 430672 5296
rect 390704 5256 430672 5284
rect 390704 5244 390710 5256
rect 430666 5244 430672 5256
rect 430724 5244 430730 5296
rect 21910 5176 21916 5228
rect 21968 5216 21974 5228
rect 240226 5216 240232 5228
rect 21968 5188 240232 5216
rect 21968 5176 21974 5188
rect 240226 5176 240232 5188
rect 240284 5176 240290 5228
rect 251450 5176 251456 5228
rect 251508 5216 251514 5228
rect 358814 5216 358820 5228
rect 251508 5188 358820 5216
rect 251508 5176 251514 5188
rect 358814 5176 358820 5188
rect 358872 5176 358878 5228
rect 387058 5176 387064 5228
rect 387116 5216 387122 5228
rect 427906 5216 427912 5228
rect 387116 5188 427912 5216
rect 387116 5176 387122 5188
rect 427906 5176 427912 5188
rect 427964 5176 427970 5228
rect 17310 5108 17316 5160
rect 17368 5148 17374 5160
rect 237466 5148 237472 5160
rect 17368 5120 237472 5148
rect 17368 5108 17374 5120
rect 237466 5108 237472 5120
rect 237524 5108 237530 5160
rect 247954 5108 247960 5160
rect 248012 5148 248018 5160
rect 356422 5148 356428 5160
rect 248012 5120 356428 5148
rect 248012 5108 248018 5120
rect 356422 5108 356428 5120
rect 356480 5108 356486 5160
rect 383562 5108 383568 5160
rect 383620 5148 383626 5160
rect 426710 5148 426716 5160
rect 383620 5120 426716 5148
rect 383620 5108 383626 5120
rect 426710 5108 426716 5120
rect 426768 5108 426774 5160
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 236086 5080 236092 5092
rect 12492 5052 236092 5080
rect 12492 5040 12498 5052
rect 236086 5040 236092 5052
rect 236144 5040 236150 5092
rect 244366 5040 244372 5092
rect 244424 5080 244430 5092
rect 354674 5080 354680 5092
rect 244424 5052 354680 5080
rect 244424 5040 244430 5052
rect 354674 5040 354680 5052
rect 354732 5040 354738 5092
rect 376386 5040 376392 5092
rect 376444 5080 376450 5092
rect 422386 5080 422392 5092
rect 376444 5052 422392 5080
rect 376444 5040 376450 5052
rect 422386 5040 422392 5052
rect 422444 5040 422450 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 233234 5012 233240 5024
rect 7708 4984 233240 5012
rect 7708 4972 7714 4984
rect 233234 4972 233240 4984
rect 233292 4972 233298 5024
rect 240778 4972 240784 5024
rect 240836 5012 240842 5024
rect 353294 5012 353300 5024
rect 240836 4984 353300 5012
rect 240836 4972 240842 4984
rect 353294 4972 353300 4984
rect 353352 4972 353358 5024
rect 365714 4972 365720 5024
rect 365772 5012 365778 5024
rect 416958 5012 416964 5024
rect 365772 4984 416964 5012
rect 365772 4972 365778 4984
rect 416958 4972 416964 4984
rect 417016 4972 417022 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 230750 4944 230756 4956
rect 2924 4916 230756 4944
rect 2924 4904 2930 4916
rect 230750 4904 230756 4916
rect 230808 4904 230814 4956
rect 237190 4904 237196 4956
rect 237248 4944 237254 4956
rect 350534 4944 350540 4956
rect 237248 4916 350540 4944
rect 237248 4904 237254 4916
rect 350534 4904 350540 4916
rect 350592 4904 350598 4956
rect 358538 4904 358544 4956
rect 358596 4944 358602 4956
rect 414106 4944 414112 4956
rect 358596 4916 414112 4944
rect 358596 4904 358602 4916
rect 414106 4904 414112 4916
rect 414164 4904 414170 4956
rect 503530 4904 503536 4956
rect 503588 4944 503594 4956
rect 529750 4944 529756 4956
rect 503588 4916 529756 4944
rect 503588 4904 503594 4916
rect 529750 4904 529756 4916
rect 529808 4904 529814 4956
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 230474 4876 230480 4888
rect 1728 4848 230480 4876
rect 1728 4836 1734 4848
rect 230474 4836 230480 4848
rect 230532 4836 230538 4888
rect 233694 4836 233700 4888
rect 233752 4876 233758 4888
rect 349154 4876 349160 4888
rect 233752 4848 349160 4876
rect 233752 4836 233758 4848
rect 349154 4836 349160 4848
rect 349212 4836 349218 4888
rect 351362 4836 351368 4888
rect 351420 4876 351426 4888
rect 410058 4876 410064 4888
rect 351420 4848 410064 4876
rect 351420 4836 351426 4848
rect 410058 4836 410064 4848
rect 410116 4836 410122 4888
rect 509142 4836 509148 4888
rect 509200 4876 509206 4888
rect 540514 4876 540520 4888
rect 509200 4848 540520 4876
rect 509200 4836 509206 4848
rect 540514 4836 540520 4848
rect 540572 4836 540578 4888
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 229094 4808 229100 4820
rect 624 4780 229100 4808
rect 624 4768 630 4780
rect 229094 4768 229100 4780
rect 229152 4768 229158 4820
rect 230106 4768 230112 4820
rect 230164 4808 230170 4820
rect 347774 4808 347780 4820
rect 230164 4780 347780 4808
rect 230164 4768 230170 4780
rect 347774 4768 347780 4780
rect 347832 4768 347838 4820
rect 347866 4768 347872 4820
rect 347924 4808 347930 4820
rect 408494 4808 408500 4820
rect 347924 4780 408500 4808
rect 347924 4768 347930 4780
rect 408494 4768 408500 4780
rect 408552 4768 408558 4820
rect 506290 4768 506296 4820
rect 506348 4808 506354 4820
rect 536926 4808 536932 4820
rect 506348 4780 536932 4808
rect 506348 4768 506354 4780
rect 536926 4768 536932 4780
rect 536984 4768 536990 4820
rect 215846 4700 215852 4752
rect 215904 4740 215910 4752
rect 339494 4740 339500 4752
rect 215904 4712 339500 4740
rect 215904 4700 215910 4712
rect 339494 4700 339500 4712
rect 339552 4700 339558 4752
rect 340690 4700 340696 4752
rect 340748 4740 340754 4752
rect 404538 4740 404544 4752
rect 340748 4712 404544 4740
rect 340748 4700 340754 4712
rect 404538 4700 404544 4712
rect 404596 4700 404602 4752
rect 404906 4700 404912 4752
rect 404964 4740 404970 4752
rect 437750 4740 437756 4752
rect 404964 4712 437756 4740
rect 404964 4700 404970 4712
rect 437750 4700 437756 4712
rect 437808 4700 437814 4752
rect 222930 4632 222936 4684
rect 222988 4672 222994 4684
rect 343634 4672 343640 4684
rect 222988 4644 343640 4672
rect 222988 4632 222994 4644
rect 343634 4632 343640 4644
rect 343692 4632 343698 4684
rect 344278 4632 344284 4684
rect 344336 4672 344342 4684
rect 405918 4672 405924 4684
rect 344336 4644 405924 4672
rect 344336 4632 344342 4644
rect 405918 4632 405924 4644
rect 405976 4632 405982 4684
rect 226518 4564 226524 4616
rect 226576 4604 226582 4616
rect 345014 4604 345020 4616
rect 226576 4576 345020 4604
rect 226576 4564 226582 4576
rect 345014 4564 345020 4576
rect 345072 4564 345078 4616
rect 356054 4564 356060 4616
rect 356112 4604 356118 4616
rect 362954 4604 362960 4616
rect 356112 4576 362960 4604
rect 356112 4564 356118 4576
rect 362954 4564 362960 4576
rect 363012 4564 363018 4616
rect 208670 4496 208676 4548
rect 208728 4536 208734 4548
rect 283558 4536 283564 4548
rect 208728 4508 283564 4536
rect 208728 4496 208734 4508
rect 283558 4496 283564 4508
rect 283616 4496 283622 4548
rect 319254 4496 319260 4548
rect 319312 4536 319318 4548
rect 393498 4536 393504 4548
rect 319312 4508 393504 4536
rect 319312 4496 319318 4508
rect 393498 4496 393504 4508
rect 393556 4496 393562 4548
rect 212258 4428 212264 4480
rect 212316 4468 212322 4480
rect 284938 4468 284944 4480
rect 212316 4440 284944 4468
rect 212316 4428 212322 4440
rect 284938 4428 284944 4440
rect 284996 4428 285002 4480
rect 322842 4428 322848 4480
rect 322900 4468 322906 4480
rect 394878 4468 394884 4480
rect 322900 4440 394884 4468
rect 322900 4428 322906 4440
rect 394878 4428 394884 4440
rect 394936 4428 394942 4480
rect 326430 4360 326436 4412
rect 326488 4400 326494 4412
rect 397454 4400 397460 4412
rect 326488 4372 397460 4400
rect 326488 4360 326494 4372
rect 397454 4360 397460 4372
rect 397512 4360 397518 4412
rect 330018 4292 330024 4344
rect 330076 4332 330082 4344
rect 399018 4332 399024 4344
rect 330076 4304 399024 4332
rect 330076 4292 330082 4304
rect 399018 4292 399024 4304
rect 399076 4292 399082 4344
rect 333606 4224 333612 4276
rect 333664 4264 333670 4276
rect 400398 4264 400404 4276
rect 333664 4236 400404 4264
rect 333664 4224 333670 4236
rect 400398 4224 400404 4236
rect 400456 4224 400462 4276
rect 406289 4267 406347 4273
rect 406289 4233 406301 4267
rect 406335 4264 406347 4267
rect 407850 4264 407856 4276
rect 406335 4236 407856 4264
rect 406335 4233 406347 4236
rect 406289 4227 406347 4233
rect 407850 4224 407856 4236
rect 407908 4224 407914 4276
rect 124214 4156 124220 4208
rect 124272 4196 124278 4208
rect 125410 4196 125416 4208
rect 124272 4168 125416 4196
rect 124272 4156 124278 4168
rect 125410 4156 125416 4168
rect 125468 4156 125474 4208
rect 140866 4156 140872 4208
rect 140924 4196 140930 4208
rect 142062 4196 142068 4208
rect 140924 4168 142068 4196
rect 140924 4156 140930 4168
rect 142062 4156 142068 4168
rect 142120 4156 142126 4208
rect 150434 4156 150440 4208
rect 150492 4196 150498 4208
rect 151630 4196 151636 4208
rect 150492 4168 151636 4196
rect 150492 4156 150498 4168
rect 151630 4156 151636 4168
rect 151688 4156 151694 4208
rect 158714 4156 158720 4208
rect 158772 4196 158778 4208
rect 159910 4196 159916 4208
rect 158772 4168 159916 4196
rect 158772 4156 158778 4168
rect 159910 4156 159916 4168
rect 159968 4156 159974 4208
rect 209866 4156 209872 4208
rect 209924 4196 209930 4208
rect 211062 4196 211068 4208
rect 209924 4168 211068 4196
rect 209924 4156 209930 4168
rect 211062 4156 211068 4168
rect 211120 4156 211126 4208
rect 314654 4196 314660 4208
rect 314488 4168 314660 4196
rect 42150 4088 42156 4140
rect 42208 4128 42214 4140
rect 50338 4128 50344 4140
rect 42208 4100 50344 4128
rect 42208 4088 42214 4100
rect 50338 4088 50344 4100
rect 50396 4088 50402 4140
rect 57606 4088 57612 4140
rect 57664 4128 57670 4140
rect 255958 4128 255964 4140
rect 57664 4100 255964 4128
rect 57664 4088 57670 4100
rect 255958 4088 255964 4100
rect 256016 4088 256022 4140
rect 276474 4088 276480 4140
rect 276532 4128 276538 4140
rect 314488 4128 314516 4168
rect 314654 4156 314660 4168
rect 314712 4156 314718 4208
rect 337102 4156 337108 4208
rect 337160 4196 337166 4208
rect 403066 4196 403072 4208
rect 337160 4168 403072 4196
rect 337160 4156 337166 4168
rect 403066 4156 403072 4168
rect 403124 4156 403130 4208
rect 404998 4196 405004 4208
rect 403452 4168 405004 4196
rect 276532 4100 314516 4128
rect 276532 4088 276538 4100
rect 314562 4088 314568 4140
rect 314620 4128 314626 4140
rect 316678 4128 316684 4140
rect 314620 4100 316684 4128
rect 314620 4088 314626 4100
rect 316678 4088 316684 4100
rect 316736 4088 316742 4140
rect 321646 4088 321652 4140
rect 321704 4128 321710 4140
rect 322750 4128 322756 4140
rect 321704 4100 322756 4128
rect 321704 4088 321710 4100
rect 322750 4088 322756 4100
rect 322808 4088 322814 4140
rect 331214 4088 331220 4140
rect 331272 4128 331278 4140
rect 332502 4128 332508 4140
rect 331272 4100 332508 4128
rect 331272 4088 331278 4100
rect 332502 4088 332508 4100
rect 332560 4088 332566 4140
rect 346670 4088 346676 4140
rect 346728 4128 346734 4140
rect 393961 4131 394019 4137
rect 393961 4128 393973 4131
rect 346728 4100 393973 4128
rect 346728 4088 346734 4100
rect 393961 4097 393973 4100
rect 394007 4097 394019 4131
rect 393961 4091 394019 4097
rect 50522 4020 50528 4072
rect 50580 4060 50586 4072
rect 253198 4060 253204 4072
rect 50580 4032 253204 4060
rect 50580 4020 50586 4032
rect 253198 4020 253204 4032
rect 253256 4020 253262 4072
rect 262214 4020 262220 4072
rect 262272 4060 262278 4072
rect 322658 4060 322664 4072
rect 262272 4032 322664 4060
rect 262272 4020 262278 4032
rect 322658 4020 322664 4032
rect 322716 4020 322722 4072
rect 339494 4020 339500 4072
rect 339552 4060 339558 4072
rect 392949 4063 393007 4069
rect 392949 4060 392961 4063
rect 339552 4032 392961 4060
rect 339552 4020 339558 4032
rect 392949 4029 392961 4032
rect 392995 4029 393007 4063
rect 392949 4023 393007 4029
rect 393869 4063 393927 4069
rect 393869 4029 393881 4063
rect 393915 4060 393927 4063
rect 403452 4060 403480 4168
rect 404998 4156 405004 4168
rect 405056 4156 405062 4208
rect 412008 4168 412680 4196
rect 403529 4131 403587 4137
rect 403529 4097 403541 4131
rect 403575 4128 403587 4131
rect 409233 4131 409291 4137
rect 409233 4128 409245 4131
rect 403575 4100 409245 4128
rect 403575 4097 403587 4100
rect 403529 4091 403587 4097
rect 409233 4097 409245 4100
rect 409279 4097 409291 4131
rect 412008 4128 412036 4168
rect 409233 4091 409291 4097
rect 410812 4100 412036 4128
rect 408313 4063 408371 4069
rect 408313 4060 408325 4063
rect 393915 4032 403480 4060
rect 403544 4032 408325 4060
rect 393915 4029 393927 4032
rect 393869 4023 393927 4029
rect 34974 3952 34980 4004
rect 35032 3992 35038 4004
rect 46198 3992 46204 4004
rect 35032 3964 46204 3992
rect 35032 3952 35038 3964
rect 46198 3952 46204 3964
rect 46256 3952 46262 4004
rect 46934 3952 46940 4004
rect 46992 3992 46998 4004
rect 252738 3992 252744 4004
rect 46992 3964 252744 3992
rect 46992 3952 46998 3964
rect 252738 3952 252744 3964
rect 252796 3952 252802 4004
rect 271690 3952 271696 4004
rect 271748 3992 271754 4004
rect 282181 3995 282239 4001
rect 282181 3992 282193 3995
rect 271748 3964 282193 3992
rect 271748 3952 271754 3964
rect 282181 3961 282193 3964
rect 282227 3961 282239 3995
rect 282181 3955 282239 3961
rect 282273 3995 282331 4001
rect 282273 3961 282285 3995
rect 282319 3992 282331 3995
rect 283466 3992 283472 4004
rect 282319 3964 283472 3992
rect 282319 3961 282331 3964
rect 282273 3955 282331 3961
rect 283466 3952 283472 3964
rect 283524 3952 283530 4004
rect 300302 3952 300308 4004
rect 300360 3992 300366 4004
rect 363690 3992 363696 4004
rect 300360 3964 363696 3992
rect 300360 3952 300366 3964
rect 363690 3952 363696 3964
rect 363748 3952 363754 4004
rect 364518 3952 364524 4004
rect 364576 3992 364582 4004
rect 366450 3992 366456 4004
rect 364576 3964 366456 3992
rect 364576 3952 364582 3964
rect 366450 3952 366456 3964
rect 366508 3952 366514 4004
rect 374641 3995 374699 4001
rect 374641 3961 374653 3995
rect 374687 3992 374699 3995
rect 403544 3992 403572 4032
rect 408313 4029 408325 4032
rect 408359 4029 408371 4063
rect 408313 4023 408371 4029
rect 408402 4020 408408 4072
rect 408460 4060 408466 4072
rect 410812 4060 410840 4100
rect 412082 4088 412088 4140
rect 412140 4128 412146 4140
rect 412542 4128 412548 4140
rect 412140 4100 412548 4128
rect 412140 4088 412146 4100
rect 412542 4088 412548 4100
rect 412600 4088 412606 4140
rect 412652 4128 412680 4168
rect 429856 4168 430620 4196
rect 414658 4128 414664 4140
rect 412652 4100 414664 4128
rect 414658 4088 414664 4100
rect 414716 4088 414722 4140
rect 415670 4088 415676 4140
rect 415728 4128 415734 4140
rect 416682 4128 416688 4140
rect 415728 4100 416688 4128
rect 415728 4088 415734 4100
rect 416682 4088 416688 4100
rect 416740 4088 416746 4140
rect 419166 4088 419172 4140
rect 419224 4128 419230 4140
rect 420270 4128 420276 4140
rect 419224 4100 420276 4128
rect 419224 4088 419230 4100
rect 420270 4088 420276 4100
rect 420328 4088 420334 4140
rect 420362 4088 420368 4140
rect 420420 4128 420426 4140
rect 420822 4128 420828 4140
rect 420420 4100 420828 4128
rect 420420 4088 420426 4100
rect 420822 4088 420828 4100
rect 420880 4088 420886 4140
rect 421558 4088 421564 4140
rect 421616 4128 421622 4140
rect 422202 4128 422208 4140
rect 421616 4100 422208 4128
rect 421616 4088 421622 4100
rect 422202 4088 422208 4100
rect 422260 4088 422266 4140
rect 422754 4088 422760 4140
rect 422812 4128 422818 4140
rect 423582 4128 423588 4140
rect 422812 4100 423588 4128
rect 422812 4088 422818 4100
rect 423582 4088 423588 4100
rect 423640 4088 423646 4140
rect 423677 4131 423735 4137
rect 423677 4097 423689 4131
rect 423723 4128 423735 4131
rect 429856 4128 429884 4168
rect 430592 4140 430620 4168
rect 423723 4100 429884 4128
rect 423723 4097 423735 4100
rect 423677 4091 423735 4097
rect 429930 4088 429936 4140
rect 429988 4128 429994 4140
rect 430482 4128 430488 4140
rect 429988 4100 430488 4128
rect 429988 4088 429994 4100
rect 430482 4088 430488 4100
rect 430540 4088 430546 4140
rect 430574 4088 430580 4140
rect 430632 4088 430638 4140
rect 431126 4088 431132 4140
rect 431184 4128 431190 4140
rect 431862 4128 431868 4140
rect 431184 4100 431868 4128
rect 431184 4088 431190 4100
rect 431862 4088 431868 4100
rect 431920 4088 431926 4140
rect 433518 4088 433524 4140
rect 433576 4128 433582 4140
rect 434622 4128 434628 4140
rect 433576 4100 434628 4128
rect 433576 4088 433582 4100
rect 434622 4088 434628 4100
rect 434680 4088 434686 4140
rect 437014 4088 437020 4140
rect 437072 4128 437078 4140
rect 442350 4128 442356 4140
rect 437072 4100 442356 4128
rect 437072 4088 437078 4100
rect 442350 4088 442356 4100
rect 442408 4088 442414 4140
rect 451274 4088 451280 4140
rect 451332 4128 451338 4140
rect 453390 4128 453396 4140
rect 451332 4100 453396 4128
rect 451332 4088 451338 4100
rect 453390 4088 453396 4100
rect 453448 4088 453454 4140
rect 469122 4088 469128 4140
rect 469180 4128 469186 4140
rect 469858 4128 469864 4140
rect 469180 4100 469864 4128
rect 469180 4088 469186 4100
rect 469858 4088 469864 4100
rect 469916 4088 469922 4140
rect 470318 4088 470324 4140
rect 470376 4128 470382 4140
rect 470778 4128 470784 4140
rect 470376 4100 470784 4128
rect 470376 4088 470382 4100
rect 470778 4088 470784 4100
rect 470836 4088 470842 4140
rect 472158 4088 472164 4140
rect 472216 4128 472222 4140
rect 472710 4128 472716 4140
rect 472216 4100 472716 4128
rect 472216 4088 472222 4100
rect 472710 4088 472716 4100
rect 472768 4088 472774 4140
rect 473354 4088 473360 4140
rect 473412 4128 473418 4140
rect 473906 4128 473912 4140
rect 473412 4100 473912 4128
rect 473412 4088 473418 4100
rect 473906 4088 473912 4100
rect 473964 4088 473970 4140
rect 474642 4088 474648 4140
rect 474700 4128 474706 4140
rect 475102 4128 475108 4140
rect 474700 4100 475108 4128
rect 474700 4088 474706 4100
rect 475102 4088 475108 4100
rect 475160 4088 475166 4140
rect 478782 4088 478788 4140
rect 478840 4128 478846 4140
rect 482278 4128 482284 4140
rect 478840 4100 482284 4128
rect 478840 4088 478846 4100
rect 482278 4088 482284 4100
rect 482336 4088 482342 4140
rect 493962 4088 493968 4140
rect 494020 4128 494026 4140
rect 513190 4128 513196 4140
rect 494020 4100 513196 4128
rect 494020 4088 494026 4100
rect 513190 4088 513196 4100
rect 513248 4088 513254 4140
rect 517422 4088 517428 4140
rect 517480 4128 517486 4140
rect 557166 4128 557172 4140
rect 517480 4100 557172 4128
rect 517480 4088 517486 4100
rect 557166 4088 557172 4100
rect 557224 4088 557230 4140
rect 558178 4088 558184 4140
rect 558236 4128 558242 4140
rect 576210 4128 576216 4140
rect 558236 4100 576216 4128
rect 558236 4088 558242 4100
rect 576210 4088 576216 4100
rect 576268 4088 576274 4140
rect 408460 4032 410840 4060
rect 408460 4020 408466 4032
rect 410886 4020 410892 4072
rect 410944 4060 410950 4072
rect 413370 4060 413376 4072
rect 410944 4032 413376 4060
rect 410944 4020 410950 4032
rect 413370 4020 413376 4032
rect 413428 4020 413434 4072
rect 414474 4020 414480 4072
rect 414532 4060 414538 4072
rect 416130 4060 416136 4072
rect 414532 4032 416136 4060
rect 414532 4020 414538 4032
rect 416130 4020 416136 4032
rect 416188 4020 416194 4072
rect 416225 4063 416283 4069
rect 416225 4029 416237 4063
rect 416271 4060 416283 4063
rect 438946 4060 438952 4072
rect 416271 4032 438952 4060
rect 416271 4029 416283 4032
rect 416225 4023 416283 4029
rect 438946 4020 438952 4032
rect 439004 4020 439010 4072
rect 440602 4020 440608 4072
rect 440660 4060 440666 4072
rect 445018 4060 445024 4072
rect 440660 4032 445024 4060
rect 440660 4020 440666 4032
rect 445018 4020 445024 4032
rect 445076 4020 445082 4072
rect 445386 4020 445392 4072
rect 445444 4060 445450 4072
rect 451918 4060 451924 4072
rect 445444 4032 451924 4060
rect 445444 4020 445450 4032
rect 451918 4020 451924 4032
rect 451976 4020 451982 4072
rect 454862 4020 454868 4072
rect 454920 4060 454926 4072
rect 456058 4060 456064 4072
rect 454920 4032 456064 4060
rect 454920 4020 454926 4032
rect 456058 4020 456064 4032
rect 456116 4020 456122 4072
rect 477402 4020 477408 4072
rect 477460 4060 477466 4072
rect 479886 4060 479892 4072
rect 477460 4032 479892 4060
rect 477460 4020 477466 4032
rect 479886 4020 479892 4032
rect 479944 4020 479950 4072
rect 492582 4020 492588 4072
rect 492640 4060 492646 4072
rect 509602 4060 509608 4072
rect 492640 4032 509608 4060
rect 492640 4020 492646 4032
rect 509602 4020 509608 4032
rect 509660 4020 509666 4072
rect 510522 4020 510528 4072
rect 510580 4060 510586 4072
rect 516965 4063 517023 4069
rect 516965 4060 516977 4063
rect 510580 4032 516977 4060
rect 510580 4020 510586 4032
rect 516965 4029 516977 4032
rect 517011 4029 517023 4063
rect 516965 4023 517023 4029
rect 518802 4020 518808 4072
rect 518860 4060 518866 4072
rect 559558 4060 559564 4072
rect 518860 4032 559564 4060
rect 518860 4020 518866 4032
rect 559558 4020 559564 4032
rect 559616 4020 559622 4072
rect 374687 3964 403572 3992
rect 403621 3995 403679 4001
rect 374687 3961 374699 3964
rect 374641 3955 374699 3961
rect 403621 3961 403633 3995
rect 403667 3992 403679 3995
rect 409138 3992 409144 4004
rect 403667 3964 409144 3992
rect 403667 3961 403679 3964
rect 403621 3955 403679 3961
rect 409138 3952 409144 3964
rect 409196 3952 409202 4004
rect 409233 3995 409291 4001
rect 409233 3961 409245 3995
rect 409279 3992 409291 3995
rect 424410 3992 424416 4004
rect 409279 3964 424416 3992
rect 409279 3961 409291 3964
rect 409233 3955 409291 3961
rect 424410 3952 424416 3964
rect 424468 3952 424474 4004
rect 427538 3952 427544 4004
rect 427596 3992 427602 4004
rect 432693 3995 432751 4001
rect 427596 3964 432644 3992
rect 427596 3952 427602 3964
rect 45738 3884 45744 3936
rect 45796 3924 45802 3936
rect 251818 3924 251824 3936
rect 45796 3896 251824 3924
rect 45796 3884 45802 3896
rect 251818 3884 251824 3896
rect 251876 3884 251882 3936
rect 258626 3884 258632 3936
rect 258684 3924 258690 3936
rect 322566 3924 322572 3936
rect 258684 3896 322572 3924
rect 258684 3884 258690 3896
rect 322566 3884 322572 3896
rect 322624 3884 322630 3936
rect 325234 3884 325240 3936
rect 325292 3924 325298 3936
rect 391198 3924 391204 3936
rect 325292 3896 391204 3924
rect 325292 3884 325298 3896
rect 391198 3884 391204 3896
rect 391256 3884 391262 3936
rect 392949 3927 393007 3933
rect 392949 3893 392961 3927
rect 392995 3924 393007 3927
rect 396718 3924 396724 3936
rect 392995 3896 396724 3924
rect 392995 3893 393007 3896
rect 392949 3887 393007 3893
rect 396718 3884 396724 3896
rect 396776 3884 396782 3936
rect 400214 3884 400220 3936
rect 400272 3924 400278 3936
rect 432414 3924 432420 3936
rect 400272 3896 432420 3924
rect 400272 3884 400278 3896
rect 432414 3884 432420 3896
rect 432472 3884 432478 3936
rect 432616 3924 432644 3964
rect 432693 3961 432705 3995
rect 432739 3992 432751 3995
rect 448514 3992 448520 4004
rect 432739 3964 448520 3992
rect 432739 3961 432751 3964
rect 432693 3955 432751 3961
rect 448514 3952 448520 3964
rect 448572 3952 448578 4004
rect 456150 3952 456156 4004
rect 456208 3992 456214 4004
rect 462958 3992 462964 4004
rect 456208 3964 462964 3992
rect 456208 3952 456214 3964
rect 462958 3952 462964 3964
rect 463016 3952 463022 4004
rect 493870 3952 493876 4004
rect 493928 3992 493934 4004
rect 511994 3992 512000 4004
rect 493928 3964 512000 3992
rect 493928 3952 493934 3964
rect 511994 3952 512000 3964
rect 512052 3952 512058 4004
rect 520090 3952 520096 4004
rect 520148 3992 520154 4004
rect 561950 3992 561956 4004
rect 520148 3964 561956 3992
rect 520148 3952 520154 3964
rect 561950 3952 561956 3964
rect 562008 3952 562014 4004
rect 442258 3924 442264 3936
rect 432616 3896 442264 3924
rect 442258 3884 442264 3896
rect 442316 3884 442322 3936
rect 496078 3884 496084 3936
rect 496136 3924 496142 3936
rect 515582 3924 515588 3936
rect 496136 3896 515588 3924
rect 496136 3884 496142 3896
rect 515582 3884 515588 3896
rect 515640 3884 515646 3936
rect 520182 3884 520188 3936
rect 520240 3924 520246 3936
rect 564342 3924 564348 3936
rect 520240 3896 564348 3924
rect 520240 3884 520246 3896
rect 564342 3884 564348 3896
rect 564400 3884 564406 3936
rect 565078 3884 565084 3936
rect 565136 3924 565142 3936
rect 579798 3924 579804 3936
rect 565136 3896 579804 3924
rect 565136 3884 565142 3896
rect 579798 3884 579804 3896
rect 579856 3884 579862 3936
rect 38562 3816 38568 3868
rect 38620 3856 38626 3868
rect 248414 3856 248420 3868
rect 38620 3828 248420 3856
rect 38620 3816 38626 3828
rect 248414 3816 248420 3828
rect 248472 3816 248478 3868
rect 255038 3816 255044 3868
rect 255096 3856 255102 3868
rect 255096 3828 316724 3856
rect 255096 3816 255102 3828
rect 39758 3748 39764 3800
rect 39816 3788 39822 3800
rect 249794 3788 249800 3800
rect 39816 3760 249800 3788
rect 39816 3748 39822 3760
rect 249794 3748 249800 3760
rect 249852 3748 249858 3800
rect 272886 3748 272892 3800
rect 272944 3788 272950 3800
rect 316586 3788 316592 3800
rect 272944 3760 316592 3788
rect 272944 3748 272950 3760
rect 316586 3748 316592 3760
rect 316644 3748 316650 3800
rect 32674 3680 32680 3732
rect 32732 3720 32738 3732
rect 245654 3720 245660 3732
rect 32732 3692 245660 3720
rect 32732 3680 32738 3692
rect 245654 3680 245660 3692
rect 245712 3680 245718 3732
rect 264606 3680 264612 3732
rect 264664 3720 264670 3732
rect 282089 3723 282147 3729
rect 282089 3720 282101 3723
rect 264664 3692 282101 3720
rect 264664 3680 264670 3692
rect 282089 3689 282101 3692
rect 282135 3689 282147 3723
rect 282089 3683 282147 3689
rect 282181 3723 282239 3729
rect 282181 3689 282193 3723
rect 282227 3720 282239 3723
rect 287698 3720 287704 3732
rect 282227 3692 287704 3720
rect 282227 3689 282239 3692
rect 282181 3683 282239 3689
rect 287698 3680 287704 3692
rect 287756 3680 287762 3732
rect 299106 3680 299112 3732
rect 299164 3720 299170 3732
rect 300946 3720 300952 3732
rect 299164 3692 300952 3720
rect 299164 3680 299170 3692
rect 300946 3680 300952 3692
rect 301004 3680 301010 3732
rect 307386 3680 307392 3732
rect 307444 3720 307450 3732
rect 309778 3720 309784 3732
rect 307444 3692 309784 3720
rect 307444 3680 307450 3692
rect 309778 3680 309784 3692
rect 309836 3680 309842 3732
rect 316696 3720 316724 3828
rect 316954 3816 316960 3868
rect 317012 3856 317018 3868
rect 327074 3856 327080 3868
rect 317012 3828 327080 3856
rect 317012 3816 317018 3828
rect 327074 3816 327080 3828
rect 327132 3816 327138 3868
rect 332410 3816 332416 3868
rect 332468 3856 332474 3868
rect 393961 3859 394019 3865
rect 332468 3828 392256 3856
rect 332468 3816 332474 3828
rect 318058 3748 318064 3800
rect 318116 3788 318122 3800
rect 389818 3788 389824 3800
rect 318116 3760 389824 3788
rect 318116 3748 318122 3760
rect 389818 3748 389824 3760
rect 389876 3748 389882 3800
rect 392228 3788 392256 3828
rect 393961 3825 393973 3859
rect 394007 3856 394019 3859
rect 400858 3856 400864 3868
rect 394007 3828 400864 3856
rect 394007 3825 394019 3828
rect 393961 3819 394019 3825
rect 400858 3816 400864 3828
rect 400916 3816 400922 3868
rect 402514 3816 402520 3868
rect 402572 3856 402578 3868
rect 403529 3859 403587 3865
rect 403529 3856 403541 3859
rect 402572 3828 403541 3856
rect 402572 3816 402578 3828
rect 403529 3825 403541 3828
rect 403575 3825 403587 3859
rect 403529 3819 403587 3825
rect 403710 3816 403716 3868
rect 403768 3856 403774 3868
rect 437658 3856 437664 3868
rect 403768 3828 437664 3856
rect 403768 3816 403774 3828
rect 437658 3816 437664 3828
rect 437716 3816 437722 3868
rect 448974 3816 448980 3868
rect 449032 3856 449038 3868
rect 453298 3856 453304 3868
rect 449032 3828 453304 3856
rect 449032 3816 449038 3828
rect 453298 3816 453304 3828
rect 453356 3816 453362 3868
rect 467926 3816 467932 3868
rect 467984 3856 467990 3868
rect 470686 3856 470692 3868
rect 467984 3828 470692 3856
rect 467984 3816 467990 3828
rect 470686 3816 470692 3828
rect 470744 3816 470750 3868
rect 482830 3816 482836 3868
rect 482888 3856 482894 3868
rect 490558 3856 490564 3868
rect 482888 3828 490564 3856
rect 482888 3816 482894 3828
rect 490558 3816 490564 3828
rect 490616 3816 490622 3868
rect 496722 3816 496728 3868
rect 496780 3856 496786 3868
rect 509789 3859 509847 3865
rect 509789 3856 509801 3859
rect 496780 3828 509801 3856
rect 496780 3816 496786 3828
rect 509789 3825 509801 3828
rect 509835 3825 509847 3859
rect 509789 3819 509847 3825
rect 509878 3816 509884 3868
rect 509936 3856 509942 3868
rect 520274 3856 520280 3868
rect 509936 3828 520280 3856
rect 509936 3816 509942 3828
rect 520274 3816 520280 3828
rect 520332 3816 520338 3868
rect 521562 3816 521568 3868
rect 521620 3856 521626 3868
rect 566734 3856 566740 3868
rect 521620 3828 566740 3856
rect 521620 3816 521626 3828
rect 566734 3816 566740 3828
rect 566792 3816 566798 3868
rect 395338 3788 395344 3800
rect 392228 3760 395344 3788
rect 395338 3748 395344 3760
rect 395396 3748 395402 3800
rect 399018 3748 399024 3800
rect 399076 3788 399082 3800
rect 434806 3788 434812 3800
rect 399076 3760 434812 3788
rect 399076 3748 399082 3760
rect 434806 3748 434812 3760
rect 434864 3748 434870 3800
rect 438210 3748 438216 3800
rect 438268 3788 438274 3800
rect 447778 3788 447784 3800
rect 438268 3760 447784 3788
rect 438268 3748 438274 3760
rect 447778 3748 447784 3760
rect 447836 3748 447842 3800
rect 459646 3748 459652 3800
rect 459704 3788 459710 3800
rect 464338 3788 464344 3800
rect 459704 3760 464344 3788
rect 459704 3748 459710 3760
rect 464338 3748 464344 3760
rect 464396 3748 464402 3800
rect 489178 3748 489184 3800
rect 489236 3788 489242 3800
rect 497734 3788 497740 3800
rect 489236 3760 497740 3788
rect 489236 3748 489242 3760
rect 497734 3748 497740 3760
rect 497792 3748 497798 3800
rect 500862 3748 500868 3800
rect 500920 3788 500926 3800
rect 525058 3788 525064 3800
rect 500920 3760 525064 3788
rect 500920 3748 500926 3760
rect 525058 3748 525064 3760
rect 525116 3748 525122 3800
rect 525610 3748 525616 3800
rect 525668 3788 525674 3800
rect 572622 3788 572628 3800
rect 525668 3760 572628 3788
rect 525668 3748 525674 3760
rect 572622 3748 572628 3760
rect 572680 3748 572686 3800
rect 325326 3720 325332 3732
rect 316696 3692 325332 3720
rect 325326 3680 325332 3692
rect 325384 3680 325390 3732
rect 352558 3680 352564 3732
rect 352616 3720 352622 3732
rect 353202 3720 353208 3732
rect 352616 3692 353208 3720
rect 352616 3680 352622 3692
rect 353202 3680 353208 3692
rect 353260 3680 353266 3732
rect 372801 3723 372859 3729
rect 372801 3689 372813 3723
rect 372847 3720 372859 3723
rect 378410 3720 378416 3732
rect 372847 3692 378416 3720
rect 372847 3689 372859 3692
rect 372801 3683 372859 3689
rect 378410 3680 378416 3692
rect 378468 3680 378474 3732
rect 385862 3680 385868 3732
rect 385920 3720 385926 3732
rect 403621 3723 403679 3729
rect 403621 3720 403633 3723
rect 385920 3692 403633 3720
rect 385920 3680 385926 3692
rect 403621 3689 403633 3692
rect 403667 3689 403679 3723
rect 403621 3683 403679 3689
rect 403713 3723 403771 3729
rect 403713 3689 403725 3723
rect 403759 3720 403771 3723
rect 433334 3720 433340 3732
rect 403759 3692 433340 3720
rect 403759 3689 403771 3692
rect 403713 3683 403771 3689
rect 433334 3680 433340 3692
rect 433392 3680 433398 3732
rect 434530 3680 434536 3732
rect 434588 3720 434594 3732
rect 446398 3720 446404 3732
rect 434588 3692 446404 3720
rect 434588 3680 434594 3692
rect 446398 3680 446404 3692
rect 446456 3680 446462 3732
rect 450170 3680 450176 3732
rect 450228 3720 450234 3732
rect 451182 3720 451188 3732
rect 450228 3692 451188 3720
rect 450228 3680 450234 3692
rect 451182 3680 451188 3692
rect 451240 3680 451246 3732
rect 466822 3680 466828 3732
rect 466880 3720 466886 3732
rect 467742 3720 467748 3732
rect 466880 3692 467748 3720
rect 466880 3680 466886 3692
rect 467742 3680 467748 3692
rect 467800 3680 467806 3732
rect 485682 3680 485688 3732
rect 485740 3720 485746 3732
rect 495342 3720 495348 3732
rect 485740 3692 495348 3720
rect 485740 3680 485746 3692
rect 495342 3680 495348 3692
rect 495400 3680 495406 3732
rect 498838 3680 498844 3732
rect 498896 3720 498902 3732
rect 519078 3720 519084 3732
rect 498896 3692 519084 3720
rect 498896 3680 498902 3692
rect 519078 3680 519084 3692
rect 519136 3680 519142 3732
rect 522942 3680 522948 3732
rect 523000 3720 523006 3732
rect 569034 3720 569040 3732
rect 523000 3692 569040 3720
rect 523000 3680 523006 3692
rect 569034 3680 569040 3692
rect 569092 3680 569098 3732
rect 25498 3612 25504 3664
rect 25556 3652 25562 3664
rect 238205 3655 238263 3661
rect 238205 3652 238217 3655
rect 25556 3624 238217 3652
rect 25556 3612 25562 3624
rect 238205 3621 238217 3624
rect 238251 3621 238263 3655
rect 238205 3615 238263 3621
rect 239582 3612 239588 3664
rect 239640 3652 239646 3664
rect 240042 3652 240048 3664
rect 239640 3624 240048 3652
rect 239640 3612 239646 3624
rect 240042 3612 240048 3624
rect 240100 3612 240106 3664
rect 243170 3612 243176 3664
rect 243228 3652 243234 3664
rect 244182 3652 244188 3664
rect 243228 3624 244188 3652
rect 243228 3612 243234 3624
rect 244182 3612 244188 3624
rect 244240 3612 244246 3664
rect 269298 3612 269304 3664
rect 269356 3652 269362 3664
rect 289814 3652 289820 3664
rect 269356 3624 289820 3652
rect 269356 3612 269362 3624
rect 289814 3612 289820 3624
rect 289872 3612 289878 3664
rect 291930 3612 291936 3664
rect 291988 3652 291994 3664
rect 299658 3652 299664 3664
rect 291988 3624 299664 3652
rect 291988 3612 291994 3624
rect 299658 3612 299664 3624
rect 299716 3612 299722 3664
rect 303798 3612 303804 3664
rect 303856 3652 303862 3664
rect 382918 3652 382924 3664
rect 303856 3624 382924 3652
rect 303856 3612 303862 3624
rect 382918 3612 382924 3624
rect 382976 3612 382982 3664
rect 388254 3612 388260 3664
rect 388312 3652 388318 3664
rect 389082 3652 389088 3664
rect 388312 3624 389088 3652
rect 388312 3612 388318 3624
rect 389082 3612 389088 3624
rect 389140 3612 389146 3664
rect 391842 3612 391848 3664
rect 391900 3652 391906 3664
rect 408310 3652 408316 3664
rect 391900 3624 408316 3652
rect 391900 3612 391906 3624
rect 408310 3612 408316 3624
rect 408368 3612 408374 3664
rect 408405 3655 408463 3661
rect 408405 3621 408417 3655
rect 408451 3652 408463 3655
rect 408497 3655 408555 3661
rect 408497 3652 408509 3655
rect 408451 3624 408509 3652
rect 408451 3621 408463 3624
rect 408405 3615 408463 3621
rect 408497 3621 408509 3624
rect 408543 3621 408555 3655
rect 408497 3615 408555 3621
rect 408586 3612 408592 3664
rect 408644 3652 408650 3664
rect 423677 3655 423735 3661
rect 423677 3652 423689 3655
rect 408644 3624 423689 3652
rect 408644 3612 408650 3624
rect 423677 3621 423689 3624
rect 423723 3621 423735 3655
rect 423677 3615 423735 3621
rect 423769 3655 423827 3661
rect 423769 3621 423781 3655
rect 423815 3652 423827 3655
rect 426618 3652 426624 3664
rect 423815 3624 426624 3652
rect 423815 3621 423827 3624
rect 423769 3615 423827 3621
rect 426618 3612 426624 3624
rect 426676 3612 426682 3664
rect 426713 3655 426771 3661
rect 426713 3621 426725 3655
rect 426759 3652 426771 3655
rect 429286 3652 429292 3664
rect 426759 3624 429292 3652
rect 426759 3621 426771 3624
rect 426713 3615 426771 3621
rect 429286 3612 429292 3624
rect 429344 3612 429350 3664
rect 442994 3612 443000 3664
rect 443052 3652 443058 3664
rect 456978 3652 456984 3664
rect 443052 3624 456984 3652
rect 443052 3612 443058 3624
rect 456978 3612 456984 3624
rect 457036 3612 457042 3664
rect 458450 3612 458456 3664
rect 458508 3652 458514 3664
rect 464430 3652 464436 3664
rect 458508 3624 464436 3652
rect 458508 3612 458514 3624
rect 464430 3612 464436 3624
rect 464488 3612 464494 3664
rect 484302 3612 484308 3664
rect 484360 3652 484366 3664
rect 492950 3652 492956 3664
rect 484360 3624 492956 3652
rect 484360 3612 484366 3624
rect 492950 3612 492956 3624
rect 493008 3612 493014 3664
rect 499482 3612 499488 3664
rect 499540 3652 499546 3664
rect 522666 3652 522672 3664
rect 499540 3624 522672 3652
rect 499540 3612 499546 3624
rect 522666 3612 522672 3624
rect 522724 3612 522730 3664
rect 524322 3612 524328 3664
rect 524380 3652 524386 3664
rect 571426 3652 571432 3664
rect 524380 3624 571432 3652
rect 524380 3612 524386 3624
rect 571426 3612 571432 3624
rect 571484 3612 571490 3664
rect 18322 3544 18328 3596
rect 18380 3584 18386 3596
rect 19242 3584 19248 3596
rect 18380 3556 19248 3584
rect 18380 3544 18386 3556
rect 19242 3544 19248 3556
rect 19300 3544 19306 3596
rect 19518 3544 19524 3596
rect 19576 3584 19582 3596
rect 24118 3584 24124 3596
rect 19576 3556 24124 3584
rect 19576 3544 19582 3556
rect 24118 3544 24124 3556
rect 24176 3544 24182 3596
rect 24302 3544 24308 3596
rect 24360 3584 24366 3596
rect 241514 3584 241520 3596
rect 24360 3556 241520 3584
rect 24360 3544 24366 3556
rect 241514 3544 241520 3556
rect 241572 3544 241578 3596
rect 275278 3544 275284 3596
rect 275336 3584 275342 3596
rect 276658 3584 276664 3596
rect 275336 3556 276664 3584
rect 275336 3544 275342 3556
rect 276658 3544 276664 3556
rect 276716 3544 276722 3596
rect 276753 3587 276811 3593
rect 276753 3553 276765 3587
rect 276799 3584 276811 3587
rect 276799 3556 287744 3584
rect 276799 3553 276811 3556
rect 276753 3547 276811 3553
rect 16022 3476 16028 3528
rect 16080 3516 16086 3528
rect 237558 3516 237564 3528
rect 16080 3488 237564 3516
rect 16080 3476 16086 3488
rect 237558 3476 237564 3488
rect 237616 3476 237622 3528
rect 238205 3519 238263 3525
rect 238205 3485 238217 3519
rect 238251 3516 238263 3519
rect 241790 3516 241796 3528
rect 238251 3488 241796 3516
rect 238251 3485 238263 3488
rect 238205 3479 238263 3485
rect 241790 3476 241796 3488
rect 241848 3476 241854 3528
rect 265802 3476 265808 3528
rect 265860 3516 265866 3528
rect 287606 3516 287612 3528
rect 265860 3488 287612 3516
rect 265860 3476 265866 3488
rect 287606 3476 287612 3488
rect 287664 3476 287670 3528
rect 287716 3516 287744 3556
rect 289538 3544 289544 3596
rect 289596 3584 289602 3596
rect 292577 3587 292635 3593
rect 292577 3584 292589 3587
rect 289596 3556 292589 3584
rect 289596 3544 289602 3556
rect 292577 3553 292589 3556
rect 292623 3553 292635 3587
rect 292577 3547 292635 3553
rect 296714 3544 296720 3596
rect 296772 3584 296778 3596
rect 381538 3584 381544 3596
rect 296772 3556 381544 3584
rect 296772 3544 296778 3556
rect 381538 3544 381544 3556
rect 381596 3544 381602 3596
rect 389450 3544 389456 3596
rect 389508 3584 389514 3596
rect 418157 3587 418215 3593
rect 418157 3584 418169 3587
rect 389508 3556 418169 3584
rect 389508 3544 389514 3556
rect 418157 3553 418169 3556
rect 418203 3553 418215 3587
rect 418157 3547 418215 3553
rect 439406 3544 439412 3596
rect 439464 3584 439470 3596
rect 455598 3584 455604 3596
rect 439464 3556 455604 3584
rect 439464 3544 439470 3556
rect 455598 3544 455604 3556
rect 455656 3544 455662 3596
rect 457254 3544 457260 3596
rect 457312 3584 457318 3596
rect 465074 3584 465080 3596
rect 457312 3556 465080 3584
rect 457312 3544 457318 3556
rect 465074 3544 465080 3556
rect 465132 3544 465138 3596
rect 484210 3544 484216 3596
rect 484268 3584 484274 3596
rect 494146 3584 494152 3596
rect 484268 3556 494152 3584
rect 484268 3544 484274 3556
rect 494146 3544 494152 3556
rect 494204 3544 494210 3596
rect 499390 3544 499396 3596
rect 499448 3584 499454 3596
rect 523862 3584 523868 3596
rect 499448 3556 523868 3584
rect 499448 3544 499454 3556
rect 523862 3544 523868 3556
rect 523920 3544 523926 3596
rect 525518 3544 525524 3596
rect 525576 3584 525582 3596
rect 525576 3556 570552 3584
rect 525576 3544 525582 3556
rect 289906 3516 289912 3528
rect 287716 3488 289912 3516
rect 289906 3476 289912 3488
rect 289964 3476 289970 3528
rect 302145 3519 302203 3525
rect 302145 3485 302157 3519
rect 302191 3516 302203 3519
rect 372801 3519 372859 3525
rect 372801 3516 372813 3519
rect 302191 3488 372813 3516
rect 302191 3485 302203 3488
rect 302145 3479 302203 3485
rect 372801 3485 372813 3488
rect 372847 3485 372859 3519
rect 372801 3479 372859 3485
rect 372893 3519 372951 3525
rect 372893 3485 372905 3519
rect 372939 3516 372951 3519
rect 376018 3516 376024 3528
rect 372939 3488 376024 3516
rect 372939 3485 372951 3488
rect 372893 3479 372951 3485
rect 376018 3476 376024 3488
rect 376076 3476 376082 3528
rect 382366 3476 382372 3528
rect 382424 3516 382430 3528
rect 423769 3519 423827 3525
rect 423769 3516 423781 3519
rect 382424 3488 423781 3516
rect 382424 3476 382430 3488
rect 423769 3485 423781 3488
rect 423815 3485 423827 3519
rect 423769 3479 423827 3485
rect 426342 3476 426348 3528
rect 426400 3516 426406 3528
rect 428458 3516 428464 3528
rect 426400 3488 428464 3516
rect 426400 3476 426406 3488
rect 428458 3476 428464 3488
rect 428516 3476 428522 3528
rect 452470 3476 452476 3528
rect 452528 3516 452534 3528
rect 460198 3516 460204 3528
rect 452528 3488 460204 3516
rect 452528 3476 452534 3488
rect 460198 3476 460204 3488
rect 460256 3476 460262 3528
rect 465626 3476 465632 3528
rect 465684 3516 465690 3528
rect 466362 3516 466368 3528
rect 465684 3488 466368 3516
rect 465684 3476 465690 3488
rect 466362 3476 466368 3488
rect 466420 3476 466426 3528
rect 487062 3476 487068 3528
rect 487120 3516 487126 3528
rect 498930 3516 498936 3528
rect 487120 3488 498936 3516
rect 487120 3476 487126 3488
rect 498930 3476 498936 3488
rect 498988 3476 498994 3528
rect 500770 3476 500776 3528
rect 500828 3516 500834 3528
rect 526254 3516 526260 3528
rect 500828 3488 526260 3516
rect 500828 3476 500834 3488
rect 526254 3476 526260 3488
rect 526312 3476 526318 3528
rect 528462 3476 528468 3528
rect 528520 3516 528526 3528
rect 569129 3519 569187 3525
rect 569129 3516 569141 3519
rect 528520 3488 569141 3516
rect 528520 3476 528526 3488
rect 569129 3485 569141 3488
rect 569175 3485 569187 3519
rect 569129 3479 569187 3485
rect 569218 3476 569224 3528
rect 569276 3516 569282 3528
rect 570230 3516 570236 3528
rect 569276 3488 570236 3516
rect 569276 3476 569282 3488
rect 570230 3476 570236 3488
rect 570288 3476 570294 3528
rect 570524 3516 570552 3556
rect 573358 3544 573364 3596
rect 573416 3584 573422 3596
rect 582190 3584 582196 3596
rect 573416 3556 582196 3584
rect 573416 3544 573422 3556
rect 582190 3544 582196 3556
rect 582248 3544 582254 3596
rect 573818 3516 573824 3528
rect 570524 3488 573824 3516
rect 573818 3476 573824 3488
rect 573876 3476 573882 3528
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 10318 3448 10324 3460
rect 5316 3420 10324 3448
rect 5316 3408 5322 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 14826 3408 14832 3460
rect 14884 3448 14890 3460
rect 236362 3448 236368 3460
rect 14884 3420 236368 3448
rect 14884 3408 14890 3420
rect 236362 3408 236368 3420
rect 236420 3408 236426 3460
rect 261018 3408 261024 3460
rect 261076 3448 261082 3460
rect 356054 3448 356060 3460
rect 261076 3420 356060 3448
rect 261076 3408 261082 3420
rect 356054 3408 356060 3420
rect 356112 3408 356118 3460
rect 371513 3451 371571 3457
rect 371513 3417 371525 3451
rect 371559 3448 371571 3451
rect 403805 3451 403863 3457
rect 371559 3420 403756 3448
rect 371559 3417 371571 3420
rect 371513 3411 371571 3417
rect 36170 3340 36176 3392
rect 36228 3380 36234 3392
rect 39298 3380 39304 3392
rect 36228 3352 39304 3380
rect 36228 3340 36234 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 50356 3352 58296 3380
rect 11238 3272 11244 3324
rect 11296 3312 11302 3324
rect 17218 3312 17224 3324
rect 11296 3284 17224 3312
rect 11296 3272 11302 3284
rect 17218 3272 17224 3284
rect 17276 3272 17282 3324
rect 20714 3272 20720 3324
rect 20772 3312 20778 3324
rect 28258 3312 28264 3324
rect 20772 3284 28264 3312
rect 20772 3272 20778 3284
rect 28258 3272 28264 3284
rect 28316 3272 28322 3324
rect 43346 3204 43352 3256
rect 43404 3244 43410 3256
rect 50356 3244 50384 3352
rect 54018 3272 54024 3324
rect 54076 3312 54082 3324
rect 57238 3312 57244 3324
rect 54076 3284 57244 3312
rect 54076 3272 54082 3284
rect 57238 3272 57244 3284
rect 57296 3272 57302 3324
rect 58268 3312 58296 3352
rect 59998 3340 60004 3392
rect 60056 3380 60062 3392
rect 60642 3380 60648 3392
rect 60056 3352 60648 3380
rect 60056 3340 60062 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 63586 3340 63592 3392
rect 63644 3380 63650 3392
rect 64782 3380 64788 3392
rect 63644 3352 64788 3380
rect 63644 3340 63650 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 70670 3340 70676 3392
rect 70728 3380 70734 3392
rect 71682 3380 71688 3392
rect 70728 3352 71688 3380
rect 70728 3340 70734 3352
rect 71682 3340 71688 3352
rect 71740 3340 71746 3392
rect 257338 3380 257344 3392
rect 71792 3352 257344 3380
rect 61378 3312 61384 3324
rect 58268 3284 61384 3312
rect 61378 3272 61384 3284
rect 61436 3272 61442 3324
rect 43404 3216 50384 3244
rect 43404 3204 43410 3216
rect 64782 3204 64788 3256
rect 64840 3244 64846 3256
rect 71792 3244 71820 3352
rect 257338 3340 257344 3352
rect 257396 3340 257402 3392
rect 268102 3340 268108 3392
rect 268160 3380 268166 3392
rect 276753 3383 276811 3389
rect 276753 3380 276765 3383
rect 268160 3352 276765 3380
rect 268160 3340 268166 3352
rect 276753 3349 276765 3352
rect 276799 3349 276811 3383
rect 276753 3343 276811 3349
rect 278866 3340 278872 3392
rect 278924 3380 278930 3392
rect 280062 3380 280068 3392
rect 278924 3352 280068 3380
rect 278924 3340 278930 3352
rect 280062 3340 280068 3352
rect 280120 3340 280126 3392
rect 282454 3340 282460 3392
rect 282512 3380 282518 3392
rect 294598 3380 294604 3392
rect 282512 3352 294604 3380
rect 282512 3340 282518 3352
rect 294598 3340 294604 3352
rect 294656 3340 294662 3392
rect 295518 3340 295524 3392
rect 295576 3380 295582 3392
rect 318794 3380 318800 3392
rect 295576 3352 318800 3380
rect 295576 3340 295582 3352
rect 318794 3340 318800 3352
rect 318852 3340 318858 3392
rect 324038 3340 324044 3392
rect 324096 3380 324102 3392
rect 346486 3380 346492 3392
rect 324096 3352 346492 3380
rect 324096 3340 324102 3352
rect 346486 3340 346492 3352
rect 346544 3340 346550 3392
rect 353754 3340 353760 3392
rect 353812 3380 353818 3392
rect 393869 3383 393927 3389
rect 393869 3380 393881 3383
rect 353812 3352 393881 3380
rect 353812 3340 353818 3352
rect 393869 3349 393881 3352
rect 393915 3349 393927 3383
rect 393869 3343 393927 3349
rect 396626 3340 396632 3392
rect 396684 3380 396690 3392
rect 403621 3383 403679 3389
rect 403621 3380 403633 3383
rect 396684 3352 403633 3380
rect 396684 3340 396690 3352
rect 403621 3349 403633 3352
rect 403667 3349 403679 3383
rect 403728 3380 403756 3420
rect 403805 3417 403817 3451
rect 403851 3448 403863 3451
rect 408402 3448 408408 3460
rect 403851 3420 408408 3448
rect 403851 3417 403863 3420
rect 403805 3411 403863 3417
rect 408402 3408 408408 3420
rect 408460 3408 408466 3460
rect 408494 3408 408500 3460
rect 408552 3448 408558 3460
rect 409782 3448 409788 3460
rect 408552 3420 409788 3448
rect 408552 3408 408558 3420
rect 409782 3408 409788 3420
rect 409840 3408 409846 3460
rect 409877 3451 409935 3457
rect 409877 3417 409889 3451
rect 409923 3448 409935 3451
rect 416225 3451 416283 3457
rect 416225 3448 416237 3451
rect 409923 3420 416237 3448
rect 409923 3417 409935 3420
rect 409877 3411 409935 3417
rect 416225 3417 416237 3420
rect 416271 3417 416283 3451
rect 444558 3448 444564 3460
rect 416225 3411 416283 3417
rect 422036 3420 444564 3448
rect 406289 3383 406347 3389
rect 406289 3380 406301 3383
rect 403728 3352 403848 3380
rect 403621 3343 403679 3349
rect 71866 3272 71872 3324
rect 71924 3312 71930 3324
rect 258718 3312 258724 3324
rect 71924 3284 258724 3312
rect 71924 3272 71930 3284
rect 258718 3272 258724 3284
rect 258776 3272 258782 3324
rect 292577 3315 292635 3321
rect 292577 3281 292589 3315
rect 292623 3312 292635 3315
rect 302145 3315 302203 3321
rect 302145 3312 302157 3315
rect 292623 3284 302157 3312
rect 292623 3281 292635 3284
rect 292577 3275 292635 3281
rect 302145 3281 302157 3284
rect 302191 3281 302203 3315
rect 302145 3275 302203 3281
rect 306190 3272 306196 3324
rect 306248 3312 306254 3324
rect 325602 3312 325608 3324
rect 306248 3284 325608 3312
rect 306248 3272 306254 3284
rect 325602 3272 325608 3284
rect 325660 3272 325666 3324
rect 335173 3315 335231 3321
rect 335173 3281 335185 3315
rect 335219 3312 335231 3315
rect 347958 3312 347964 3324
rect 335219 3284 347964 3312
rect 335219 3281 335231 3284
rect 335173 3275 335231 3281
rect 347958 3272 347964 3284
rect 348016 3272 348022 3324
rect 360930 3272 360936 3324
rect 360988 3312 360994 3324
rect 360988 3284 403756 3312
rect 360988 3272 360994 3284
rect 64840 3216 71820 3244
rect 64840 3204 64846 3216
rect 77846 3204 77852 3256
rect 77904 3244 77910 3256
rect 78582 3244 78588 3256
rect 77904 3216 78588 3244
rect 77904 3204 77910 3216
rect 78582 3204 78588 3216
rect 78640 3204 78646 3256
rect 81434 3204 81440 3256
rect 81492 3244 81498 3256
rect 82722 3244 82728 3256
rect 81492 3216 82728 3244
rect 81492 3204 81498 3216
rect 82722 3204 82728 3216
rect 82780 3204 82786 3256
rect 84838 3244 84844 3256
rect 82832 3216 84844 3244
rect 27890 3136 27896 3188
rect 27948 3176 27954 3188
rect 28902 3176 28908 3188
rect 27948 3148 28908 3176
rect 27948 3136 27954 3148
rect 28902 3136 28908 3148
rect 28960 3136 28966 3188
rect 29086 3136 29092 3188
rect 29144 3176 29150 3188
rect 32398 3176 32404 3188
rect 29144 3148 32404 3176
rect 29144 3136 29150 3148
rect 32398 3136 32404 3148
rect 32456 3136 32462 3188
rect 61194 3136 61200 3188
rect 61252 3176 61258 3188
rect 66898 3176 66904 3188
rect 61252 3148 66904 3176
rect 61252 3136 61258 3148
rect 66898 3136 66904 3148
rect 66956 3136 66962 3188
rect 82630 3136 82636 3188
rect 82688 3176 82694 3188
rect 82832 3176 82860 3216
rect 84838 3204 84844 3216
rect 84896 3204 84902 3256
rect 84930 3204 84936 3256
rect 84988 3244 84994 3256
rect 85482 3244 85488 3256
rect 84988 3216 85488 3244
rect 84988 3204 84994 3216
rect 85482 3204 85488 3216
rect 85540 3204 85546 3256
rect 88518 3204 88524 3256
rect 88576 3244 88582 3256
rect 89622 3244 89628 3256
rect 88576 3216 89628 3244
rect 88576 3204 88582 3216
rect 89622 3204 89628 3216
rect 89680 3204 89686 3256
rect 261478 3244 261484 3256
rect 89732 3216 261484 3244
rect 82688 3148 82860 3176
rect 82909 3179 82967 3185
rect 82688 3136 82694 3148
rect 82909 3145 82921 3179
rect 82955 3176 82967 3179
rect 89732 3176 89760 3216
rect 261478 3204 261484 3216
rect 261536 3204 261542 3256
rect 288342 3204 288348 3256
rect 288400 3244 288406 3256
rect 292942 3244 292948 3256
rect 288400 3216 292948 3244
rect 288400 3204 288406 3216
rect 292942 3204 292948 3216
rect 293000 3204 293006 3256
rect 302602 3204 302608 3256
rect 302660 3244 302666 3256
rect 320174 3244 320180 3256
rect 302660 3216 320180 3244
rect 302660 3204 302666 3216
rect 320174 3204 320180 3216
rect 320232 3204 320238 3256
rect 328822 3204 328828 3256
rect 328880 3244 328886 3256
rect 363598 3244 363604 3256
rect 328880 3216 363604 3244
rect 328880 3204 328886 3216
rect 363598 3204 363604 3216
rect 363656 3204 363662 3256
rect 370406 3204 370412 3256
rect 370464 3244 370470 3256
rect 403728 3253 403756 3284
rect 403621 3247 403679 3253
rect 403621 3244 403633 3247
rect 370464 3216 403633 3244
rect 370464 3204 370470 3216
rect 403621 3213 403633 3216
rect 403667 3213 403679 3247
rect 403621 3207 403679 3213
rect 403713 3247 403771 3253
rect 403713 3213 403725 3247
rect 403759 3213 403771 3247
rect 403820 3244 403848 3352
rect 404004 3352 406301 3380
rect 403897 3315 403955 3321
rect 403897 3281 403909 3315
rect 403943 3312 403955 3315
rect 404004 3312 404032 3352
rect 406289 3349 406301 3352
rect 406335 3349 406347 3383
rect 406289 3343 406347 3349
rect 407298 3340 407304 3392
rect 407356 3380 407362 3392
rect 409601 3383 409659 3389
rect 409601 3380 409613 3383
rect 407356 3352 409613 3380
rect 407356 3340 407362 3352
rect 409601 3349 409613 3352
rect 409647 3349 409659 3383
rect 409601 3343 409659 3349
rect 409690 3340 409696 3392
rect 409748 3380 409754 3392
rect 421929 3383 421987 3389
rect 421929 3380 421941 3383
rect 409748 3352 421941 3380
rect 409748 3340 409754 3352
rect 421929 3349 421941 3352
rect 421975 3349 421987 3383
rect 421929 3343 421987 3349
rect 403943 3284 404032 3312
rect 403943 3281 403955 3284
rect 403897 3275 403955 3281
rect 406102 3272 406108 3324
rect 406160 3312 406166 3324
rect 406160 3284 413324 3312
rect 406160 3272 406166 3284
rect 408497 3247 408555 3253
rect 408497 3244 408509 3247
rect 403820 3216 408509 3244
rect 403713 3207 403771 3213
rect 408497 3213 408509 3216
rect 408543 3213 408555 3247
rect 408497 3207 408555 3213
rect 408589 3247 408647 3253
rect 408589 3213 408601 3247
rect 408635 3244 408647 3247
rect 411898 3244 411904 3256
rect 408635 3216 411904 3244
rect 408635 3213 408647 3216
rect 408589 3207 408647 3213
rect 411898 3204 411904 3216
rect 411956 3204 411962 3256
rect 413296 3244 413324 3284
rect 416774 3272 416780 3324
rect 416832 3312 416838 3324
rect 417418 3312 417424 3324
rect 416832 3284 417424 3312
rect 416832 3272 416838 3284
rect 417418 3272 417424 3284
rect 417476 3272 417482 3324
rect 417970 3272 417976 3324
rect 418028 3312 418034 3324
rect 422036 3312 422064 3420
rect 444558 3408 444564 3420
rect 444616 3408 444622 3460
rect 446582 3408 446588 3460
rect 446640 3448 446646 3460
rect 459738 3448 459744 3460
rect 446640 3420 459744 3448
rect 446640 3408 446646 3420
rect 459738 3408 459744 3420
rect 459796 3408 459802 3460
rect 488350 3408 488356 3460
rect 488408 3448 488414 3460
rect 501230 3448 501236 3460
rect 488408 3420 501236 3448
rect 488408 3408 488414 3420
rect 501230 3408 501236 3420
rect 501288 3408 501294 3460
rect 502242 3408 502248 3460
rect 502300 3448 502306 3460
rect 528646 3448 528652 3460
rect 502300 3420 528652 3448
rect 502300 3408 502306 3420
rect 528646 3408 528652 3420
rect 528704 3408 528710 3460
rect 529842 3408 529848 3460
rect 529900 3448 529906 3460
rect 580994 3448 581000 3460
rect 529900 3420 581000 3448
rect 529900 3408 529906 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 424318 3380 424324 3392
rect 418028 3284 422064 3312
rect 422128 3352 424324 3380
rect 418028 3272 418034 3284
rect 421101 3247 421159 3253
rect 421101 3244 421113 3247
rect 413296 3216 421113 3244
rect 421101 3213 421113 3216
rect 421147 3213 421159 3247
rect 422128 3244 422156 3352
rect 424318 3340 424324 3352
rect 424376 3340 424382 3392
rect 425146 3340 425152 3392
rect 425204 3380 425210 3392
rect 425204 3352 432276 3380
rect 425204 3340 425210 3352
rect 422941 3315 422999 3321
rect 422941 3281 422953 3315
rect 422987 3312 422999 3315
rect 432248 3312 432276 3352
rect 432322 3340 432328 3392
rect 432380 3380 432386 3392
rect 447597 3383 447655 3389
rect 447597 3380 447609 3383
rect 432380 3352 447609 3380
rect 432380 3340 432386 3352
rect 447597 3349 447609 3352
rect 447643 3349 447655 3383
rect 449158 3380 449164 3392
rect 447597 3343 447655 3349
rect 447704 3352 449164 3380
rect 432693 3315 432751 3321
rect 432693 3312 432705 3315
rect 422987 3284 431632 3312
rect 432248 3284 432705 3312
rect 422987 3281 422999 3284
rect 422941 3275 422999 3281
rect 421101 3207 421159 3213
rect 421208 3216 422156 3244
rect 82955 3148 89760 3176
rect 82955 3145 82967 3148
rect 82909 3139 82967 3145
rect 89806 3136 89812 3188
rect 89864 3176 89870 3188
rect 262858 3176 262864 3188
rect 89864 3148 262864 3176
rect 89864 3136 89870 3148
rect 262858 3136 262864 3148
rect 262916 3136 262922 3188
rect 285950 3136 285956 3188
rect 286008 3176 286014 3188
rect 286962 3176 286968 3188
rect 286008 3148 286968 3176
rect 286008 3136 286014 3148
rect 286962 3136 286968 3148
rect 287020 3136 287026 3188
rect 293126 3136 293132 3188
rect 293184 3176 293190 3188
rect 293862 3176 293868 3188
rect 293184 3148 293868 3176
rect 293184 3136 293190 3148
rect 293862 3136 293868 3148
rect 293920 3136 293926 3188
rect 309778 3136 309784 3188
rect 309836 3176 309842 3188
rect 323578 3176 323584 3188
rect 309836 3148 323584 3176
rect 309836 3136 309842 3148
rect 323578 3136 323584 3148
rect 323636 3136 323642 3188
rect 327626 3136 327632 3188
rect 327684 3176 327690 3188
rect 335173 3179 335231 3185
rect 335173 3176 335185 3179
rect 327684 3148 335185 3176
rect 327684 3136 327690 3148
rect 335173 3145 335185 3148
rect 335219 3145 335231 3179
rect 335173 3139 335231 3145
rect 343082 3136 343088 3188
rect 343140 3176 343146 3188
rect 372893 3179 372951 3185
rect 372893 3176 372905 3179
rect 343140 3148 372905 3176
rect 343140 3136 343146 3148
rect 372893 3145 372905 3148
rect 372939 3145 372951 3179
rect 372893 3139 372951 3145
rect 381170 3136 381176 3188
rect 381228 3176 381234 3188
rect 421208 3176 421236 3216
rect 423950 3204 423956 3256
rect 424008 3244 424014 3256
rect 424962 3244 424968 3256
rect 424008 3216 424968 3244
rect 424008 3204 424014 3216
rect 424962 3204 424968 3216
rect 425020 3204 425026 3256
rect 381228 3148 421236 3176
rect 421929 3179 421987 3185
rect 381228 3136 381234 3148
rect 421929 3145 421941 3179
rect 421975 3176 421987 3179
rect 431218 3176 431224 3188
rect 421975 3148 431224 3176
rect 421975 3145 421987 3148
rect 421929 3139 421987 3145
rect 431218 3136 431224 3148
rect 431276 3136 431282 3188
rect 431604 3176 431632 3284
rect 432693 3281 432705 3284
rect 432739 3281 432751 3315
rect 432693 3275 432751 3281
rect 441798 3272 441804 3324
rect 441856 3312 441862 3324
rect 447704 3312 447732 3352
rect 449158 3340 449164 3352
rect 449216 3340 449222 3392
rect 482922 3340 482928 3392
rect 482980 3380 482986 3392
rect 489362 3380 489368 3392
rect 482980 3352 489368 3380
rect 482980 3340 482986 3352
rect 489362 3340 489368 3352
rect 489420 3340 489426 3392
rect 492490 3340 492496 3392
rect 492548 3380 492554 3392
rect 508406 3380 508412 3392
rect 492548 3352 508412 3380
rect 492548 3340 492554 3352
rect 508406 3340 508412 3352
rect 508464 3340 508470 3392
rect 514662 3340 514668 3392
rect 514720 3380 514726 3392
rect 552382 3380 552388 3392
rect 514720 3352 552388 3380
rect 514720 3340 514726 3352
rect 552382 3340 552388 3352
rect 552440 3340 552446 3392
rect 556798 3340 556804 3392
rect 556856 3380 556862 3392
rect 565538 3380 565544 3392
rect 556856 3352 565544 3380
rect 556856 3340 556862 3352
rect 565538 3340 565544 3352
rect 565596 3340 565602 3392
rect 569129 3383 569187 3389
rect 569129 3349 569141 3383
rect 569175 3380 569187 3383
rect 578602 3380 578608 3392
rect 569175 3352 578608 3380
rect 569175 3349 569187 3352
rect 569129 3343 569187 3349
rect 578602 3340 578608 3352
rect 578660 3340 578666 3392
rect 441856 3284 447732 3312
rect 441856 3272 441862 3284
rect 447778 3272 447784 3324
rect 447836 3312 447842 3324
rect 448422 3312 448428 3324
rect 447836 3284 448428 3312
rect 447836 3272 447842 3284
rect 448422 3272 448428 3284
rect 448480 3272 448486 3324
rect 464430 3272 464436 3324
rect 464488 3312 464494 3324
rect 464982 3312 464988 3324
rect 464488 3284 464988 3312
rect 464488 3272 464494 3284
rect 464982 3272 464988 3284
rect 465040 3272 465046 3324
rect 481542 3272 481548 3324
rect 481600 3312 481606 3324
rect 486970 3312 486976 3324
rect 481600 3284 486976 3312
rect 481600 3272 481606 3284
rect 486970 3272 486976 3284
rect 487028 3272 487034 3324
rect 488442 3272 488448 3324
rect 488500 3312 488506 3324
rect 502426 3312 502432 3324
rect 488500 3284 502432 3312
rect 488500 3272 488506 3284
rect 502426 3272 502432 3284
rect 502484 3272 502490 3324
rect 509789 3315 509847 3321
rect 509789 3281 509801 3315
rect 509835 3312 509847 3315
rect 516778 3312 516784 3324
rect 509835 3284 516784 3312
rect 509835 3281 509847 3284
rect 509789 3275 509847 3281
rect 516778 3272 516784 3284
rect 516836 3272 516842 3324
rect 540149 3315 540207 3321
rect 540149 3312 540161 3315
rect 516888 3284 540161 3312
rect 447597 3247 447655 3253
rect 447597 3213 447609 3247
rect 447643 3244 447655 3247
rect 451550 3244 451556 3256
rect 447643 3216 451556 3244
rect 447643 3213 447655 3216
rect 447597 3207 447655 3213
rect 451550 3204 451556 3216
rect 451608 3204 451614 3256
rect 485038 3204 485044 3256
rect 485096 3244 485102 3256
rect 488166 3244 488172 3256
rect 485096 3216 488172 3244
rect 485096 3204 485102 3216
rect 488166 3204 488172 3216
rect 488224 3204 488230 3256
rect 489822 3204 489828 3256
rect 489880 3244 489886 3256
rect 504818 3244 504824 3256
rect 489880 3216 504824 3244
rect 489880 3204 489886 3216
rect 504818 3204 504824 3216
rect 504876 3204 504882 3256
rect 511810 3204 511816 3256
rect 511868 3244 511874 3256
rect 516888 3244 516916 3284
rect 540149 3281 540161 3284
rect 540195 3281 540207 3315
rect 540149 3275 540207 3281
rect 540238 3272 540244 3324
rect 540296 3312 540302 3324
rect 542906 3312 542912 3324
rect 540296 3284 542912 3312
rect 540296 3272 540302 3284
rect 542906 3272 542912 3284
rect 542964 3272 542970 3324
rect 547230 3272 547236 3324
rect 547288 3312 547294 3324
rect 550082 3312 550088 3324
rect 547288 3284 550088 3312
rect 547288 3272 547294 3284
rect 550082 3272 550088 3284
rect 550140 3272 550146 3324
rect 558362 3312 558368 3324
rect 554884 3284 558368 3312
rect 511868 3216 516916 3244
rect 516965 3247 517023 3253
rect 511868 3204 511874 3216
rect 516965 3213 516977 3247
rect 517011 3244 517023 3247
rect 517011 3216 538996 3244
rect 517011 3213 517023 3216
rect 516965 3207 517023 3213
rect 435358 3176 435364 3188
rect 431604 3148 435364 3176
rect 435358 3136 435364 3148
rect 435416 3136 435422 3188
rect 493318 3136 493324 3188
rect 493376 3176 493382 3188
rect 496538 3176 496544 3188
rect 493376 3148 496544 3176
rect 493376 3136 493382 3148
rect 496538 3136 496544 3148
rect 496596 3136 496602 3188
rect 511902 3136 511908 3188
rect 511960 3176 511966 3188
rect 538968 3176 538996 3216
rect 540330 3204 540336 3256
rect 540388 3244 540394 3256
rect 544102 3244 544108 3256
rect 540388 3216 544108 3244
rect 540388 3204 540394 3216
rect 544102 3204 544108 3216
rect 544160 3204 544166 3256
rect 545758 3204 545764 3256
rect 545816 3244 545822 3256
rect 554774 3244 554780 3256
rect 545816 3216 554780 3244
rect 545816 3204 545822 3216
rect 554774 3204 554780 3216
rect 554832 3204 554838 3256
rect 545298 3176 545304 3188
rect 511960 3148 538904 3176
rect 538968 3148 545304 3176
rect 511960 3136 511966 3148
rect 95694 3068 95700 3120
rect 95752 3108 95758 3120
rect 96522 3108 96528 3120
rect 95752 3080 96528 3108
rect 95752 3068 95758 3080
rect 96522 3068 96528 3080
rect 96580 3068 96586 3120
rect 97258 3108 97264 3120
rect 96632 3080 97264 3108
rect 10042 3000 10048 3052
rect 10100 3040 10106 3052
rect 15838 3040 15844 3052
rect 10100 3012 15844 3040
rect 10100 3000 10106 3012
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 68278 3000 68284 3052
rect 68336 3040 68342 3052
rect 71038 3040 71044 3052
rect 68336 3012 71044 3040
rect 68336 3000 68342 3012
rect 71038 3000 71044 3012
rect 71096 3000 71102 3052
rect 93302 3000 93308 3052
rect 93360 3040 93366 3052
rect 96632 3040 96660 3080
rect 97258 3068 97264 3080
rect 97316 3068 97322 3120
rect 98086 3068 98092 3120
rect 98144 3108 98150 3120
rect 99190 3108 99196 3120
rect 98144 3080 99196 3108
rect 98144 3068 98150 3080
rect 99190 3068 99196 3080
rect 99248 3068 99254 3120
rect 102778 3068 102784 3120
rect 102836 3108 102842 3120
rect 103422 3108 103428 3120
rect 102836 3080 103428 3108
rect 102836 3068 102842 3080
rect 103422 3068 103428 3080
rect 103480 3068 103486 3120
rect 103974 3068 103980 3120
rect 104032 3108 104038 3120
rect 104802 3108 104808 3120
rect 104032 3080 104808 3108
rect 104032 3068 104038 3080
rect 104802 3068 104808 3080
rect 104860 3068 104866 3120
rect 106366 3068 106372 3120
rect 106424 3108 106430 3120
rect 107562 3108 107568 3120
rect 106424 3080 107568 3108
rect 106424 3068 106430 3080
rect 107562 3068 107568 3080
rect 107620 3068 107626 3120
rect 111150 3068 111156 3120
rect 111208 3108 111214 3120
rect 111702 3108 111708 3120
rect 111208 3080 111708 3108
rect 111208 3068 111214 3080
rect 111702 3068 111708 3080
rect 111760 3068 111766 3120
rect 264238 3108 264244 3120
rect 111812 3080 264244 3108
rect 93360 3012 96660 3040
rect 93360 3000 93366 3012
rect 96890 3000 96896 3052
rect 96948 3040 96954 3052
rect 111812 3040 111840 3080
rect 264238 3068 264244 3080
rect 264296 3068 264302 3120
rect 313366 3068 313372 3120
rect 313424 3108 313430 3120
rect 325510 3108 325516 3120
rect 313424 3080 325516 3108
rect 313424 3068 313430 3080
rect 325510 3068 325516 3080
rect 325568 3068 325574 3120
rect 335906 3068 335912 3120
rect 335964 3108 335970 3120
rect 366358 3108 366364 3120
rect 335964 3080 366364 3108
rect 335964 3068 335970 3080
rect 366358 3068 366364 3080
rect 366416 3068 366422 3120
rect 368014 3068 368020 3120
rect 368072 3108 368078 3120
rect 374641 3111 374699 3117
rect 374641 3108 374653 3111
rect 368072 3080 374653 3108
rect 368072 3068 368078 3080
rect 374641 3077 374653 3080
rect 374687 3077 374699 3111
rect 374641 3071 374699 3077
rect 375190 3068 375196 3120
rect 375248 3108 375254 3120
rect 403529 3111 403587 3117
rect 403529 3108 403541 3111
rect 375248 3080 403541 3108
rect 375248 3068 375254 3080
rect 403529 3077 403541 3080
rect 403575 3077 403587 3111
rect 403529 3071 403587 3077
rect 403621 3111 403679 3117
rect 403621 3077 403633 3111
rect 403667 3108 403679 3111
rect 408773 3111 408831 3117
rect 403667 3080 408724 3108
rect 403667 3077 403679 3080
rect 403621 3071 403679 3077
rect 264330 3040 264336 3052
rect 96948 3012 98776 3040
rect 96948 3000 96954 3012
rect 79042 2932 79048 2984
rect 79100 2972 79106 2984
rect 82909 2975 82967 2981
rect 82909 2972 82921 2975
rect 79100 2944 82921 2972
rect 79100 2932 79106 2944
rect 82909 2941 82921 2944
rect 82955 2941 82967 2975
rect 82909 2935 82967 2941
rect 86126 2932 86132 2984
rect 86184 2972 86190 2984
rect 98641 2975 98699 2981
rect 98641 2972 98653 2975
rect 86184 2944 98653 2972
rect 86184 2932 86190 2944
rect 98641 2941 98653 2944
rect 98687 2941 98699 2975
rect 98748 2972 98776 3012
rect 99392 3012 111840 3040
rect 111904 3012 264336 3040
rect 99392 2972 99420 3012
rect 106918 2972 106924 2984
rect 98748 2944 99420 2972
rect 100404 2944 106924 2972
rect 98641 2935 98699 2941
rect 75454 2864 75460 2916
rect 75512 2904 75518 2916
rect 100404 2904 100432 2944
rect 106918 2932 106924 2944
rect 106976 2932 106982 2984
rect 75512 2876 100432 2904
rect 75512 2864 75518 2876
rect 100478 2864 100484 2916
rect 100536 2904 100542 2916
rect 111904 2904 111932 3012
rect 264330 3000 264336 3012
rect 264388 3000 264394 3052
rect 320450 3000 320456 3052
rect 320508 3040 320514 3052
rect 328546 3040 328552 3052
rect 320508 3012 328552 3040
rect 320508 3000 320514 3012
rect 328546 3000 328552 3012
rect 328604 3000 328610 3052
rect 338298 3000 338304 3052
rect 338356 3040 338362 3052
rect 339402 3040 339408 3052
rect 338356 3012 339408 3040
rect 338356 3000 338362 3012
rect 339402 3000 339408 3012
rect 339460 3000 339466 3052
rect 350258 3000 350264 3052
rect 350316 3040 350322 3052
rect 374546 3040 374552 3052
rect 350316 3012 374552 3040
rect 350316 3000 350322 3012
rect 374546 3000 374552 3012
rect 374604 3000 374610 3052
rect 378778 3000 378784 3052
rect 378836 3040 378842 3052
rect 408586 3040 408592 3052
rect 378836 3012 408592 3040
rect 378836 3000 378842 3012
rect 408586 3000 408592 3012
rect 408644 3000 408650 3052
rect 408696 3040 408724 3080
rect 408773 3077 408785 3111
rect 408819 3108 408831 3111
rect 410610 3108 410616 3120
rect 408819 3080 410616 3108
rect 408819 3077 408831 3080
rect 408773 3071 408831 3077
rect 410610 3068 410616 3080
rect 410668 3068 410674 3120
rect 410705 3111 410763 3117
rect 410705 3077 410717 3111
rect 410751 3108 410763 3111
rect 416774 3108 416780 3120
rect 410751 3080 416780 3108
rect 410751 3077 410763 3080
rect 410705 3071 410763 3077
rect 416774 3068 416780 3080
rect 416832 3068 416838 3120
rect 416866 3068 416872 3120
rect 416924 3108 416930 3120
rect 438118 3108 438124 3120
rect 416924 3080 438124 3108
rect 416924 3068 416930 3080
rect 438118 3068 438124 3080
rect 438176 3068 438182 3120
rect 444190 3068 444196 3120
rect 444248 3108 444254 3120
rect 446490 3108 446496 3120
rect 444248 3080 446496 3108
rect 444248 3068 444254 3080
rect 446490 3068 446496 3080
rect 446548 3068 446554 3120
rect 501598 3068 501604 3120
rect 501656 3108 501662 3120
rect 506014 3108 506020 3120
rect 501656 3080 506020 3108
rect 501656 3068 501662 3080
rect 506014 3068 506020 3080
rect 506072 3068 506078 3120
rect 507762 3068 507768 3120
rect 507820 3108 507826 3120
rect 538122 3108 538128 3120
rect 507820 3080 538128 3108
rect 507820 3068 507826 3080
rect 538122 3068 538128 3080
rect 538180 3068 538186 3120
rect 538876 3108 538904 3148
rect 545298 3136 545304 3148
rect 545356 3136 545362 3188
rect 547138 3136 547144 3188
rect 547196 3176 547202 3188
rect 548886 3176 548892 3188
rect 547196 3148 548892 3176
rect 547196 3136 547202 3148
rect 548886 3136 548892 3148
rect 548944 3136 548950 3188
rect 549898 3136 549904 3188
rect 549956 3176 549962 3188
rect 554884 3176 554912 3284
rect 558362 3272 558368 3284
rect 558420 3272 558426 3324
rect 549956 3148 554912 3176
rect 549956 3136 549962 3148
rect 547690 3108 547696 3120
rect 538876 3080 547696 3108
rect 547690 3068 547696 3080
rect 547748 3068 547754 3120
rect 551186 3108 551192 3120
rect 547800 3080 551192 3108
rect 413278 3040 413284 3052
rect 408696 3012 413284 3040
rect 413278 3000 413284 3012
rect 413336 3000 413342 3052
rect 413370 3000 413376 3052
rect 413428 3040 413434 3052
rect 422941 3043 422999 3049
rect 422941 3040 422953 3043
rect 413428 3012 422953 3040
rect 413428 3000 413434 3012
rect 422941 3009 422953 3012
rect 422987 3009 422999 3043
rect 422941 3003 422999 3009
rect 506382 3000 506388 3052
rect 506440 3040 506446 3052
rect 535730 3040 535736 3052
rect 506440 3012 535736 3040
rect 506440 3000 506446 3012
rect 535730 3000 535736 3012
rect 535788 3000 535794 3052
rect 540149 3043 540207 3049
rect 540149 3009 540161 3043
rect 540195 3040 540207 3043
rect 546494 3040 546500 3052
rect 540195 3012 546500 3040
rect 540195 3009 540207 3012
rect 540149 3003 540207 3009
rect 546494 3000 546500 3012
rect 546552 3000 546558 3052
rect 112346 2932 112352 2984
rect 112404 2972 112410 2984
rect 113082 2972 113088 2984
rect 112404 2944 113088 2972
rect 112404 2932 112410 2944
rect 113082 2932 113088 2944
rect 113140 2932 113146 2984
rect 113542 2932 113548 2984
rect 113600 2972 113606 2984
rect 114462 2972 114468 2984
rect 113600 2944 114468 2972
rect 113600 2932 113606 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 115934 2932 115940 2984
rect 115992 2972 115998 2984
rect 116946 2972 116952 2984
rect 115992 2944 116952 2972
rect 115992 2932 115998 2944
rect 116946 2932 116952 2944
rect 117004 2932 117010 2984
rect 119430 2932 119436 2984
rect 119488 2972 119494 2984
rect 119982 2972 119988 2984
rect 119488 2944 119988 2972
rect 119488 2932 119494 2944
rect 119982 2932 119988 2944
rect 120040 2932 120046 2984
rect 120626 2932 120632 2984
rect 120684 2972 120690 2984
rect 121362 2972 121368 2984
rect 120684 2944 121368 2972
rect 120684 2932 120690 2944
rect 121362 2932 121368 2944
rect 121420 2932 121426 2984
rect 266906 2972 266912 2984
rect 121564 2944 266912 2972
rect 100536 2876 111932 2904
rect 100536 2864 100542 2876
rect 114738 2864 114744 2916
rect 114796 2904 114802 2916
rect 121457 2907 121515 2913
rect 121457 2904 121469 2907
rect 114796 2876 121469 2904
rect 114796 2864 114802 2876
rect 121457 2873 121469 2876
rect 121503 2873 121515 2907
rect 121457 2867 121515 2873
rect 98641 2839 98699 2845
rect 98641 2805 98653 2839
rect 98687 2836 98699 2839
rect 105538 2836 105544 2848
rect 98687 2808 105544 2836
rect 98687 2805 98699 2808
rect 98641 2799 98699 2805
rect 105538 2796 105544 2808
rect 105596 2796 105602 2848
rect 107562 2796 107568 2848
rect 107620 2836 107626 2848
rect 121564 2836 121592 2944
rect 266906 2932 266912 2944
rect 266964 2932 266970 2984
rect 341886 2932 341892 2984
rect 341944 2972 341950 2984
rect 351822 2972 351828 2984
rect 341944 2944 351828 2972
rect 341944 2932 341950 2944
rect 351822 2932 351828 2944
rect 351880 2932 351886 2984
rect 363322 2932 363328 2984
rect 363380 2972 363386 2984
rect 371513 2975 371571 2981
rect 371513 2972 371525 2975
rect 363380 2944 371525 2972
rect 363380 2932 363386 2944
rect 371513 2941 371525 2944
rect 371559 2941 371571 2975
rect 371513 2935 371571 2941
rect 371602 2932 371608 2984
rect 371660 2972 371666 2984
rect 372522 2972 372528 2984
rect 371660 2944 372528 2972
rect 371660 2932 371666 2944
rect 372522 2932 372528 2944
rect 372580 2932 372586 2984
rect 377582 2932 377588 2984
rect 377640 2972 377646 2984
rect 413462 2972 413468 2984
rect 377640 2944 413468 2972
rect 377640 2932 377646 2944
rect 413462 2932 413468 2944
rect 413520 2932 413526 2984
rect 421101 2975 421159 2981
rect 421101 2941 421113 2975
rect 421147 2972 421159 2975
rect 427078 2972 427084 2984
rect 421147 2944 427084 2972
rect 421147 2941 421159 2944
rect 421101 2935 421159 2941
rect 427078 2932 427084 2944
rect 427136 2932 427142 2984
rect 505002 2932 505008 2984
rect 505060 2972 505066 2984
rect 533430 2972 533436 2984
rect 505060 2944 533436 2972
rect 505060 2932 505066 2944
rect 533430 2932 533436 2944
rect 533488 2932 533494 2984
rect 121641 2907 121699 2913
rect 121641 2873 121653 2907
rect 121687 2904 121699 2907
rect 268378 2904 268384 2916
rect 121687 2876 268384 2904
rect 121687 2873 121699 2876
rect 121641 2867 121699 2873
rect 268378 2864 268384 2876
rect 268436 2864 268442 2916
rect 384666 2864 384672 2916
rect 384724 2904 384730 2916
rect 408497 2907 408555 2913
rect 408497 2904 408509 2907
rect 384724 2876 408509 2904
rect 384724 2864 384730 2876
rect 408497 2873 408509 2876
rect 408543 2873 408555 2907
rect 408497 2867 408555 2873
rect 408586 2864 408592 2916
rect 408644 2904 408650 2916
rect 416038 2904 416044 2916
rect 408644 2876 416044 2904
rect 408644 2864 408650 2876
rect 416038 2864 416044 2876
rect 416096 2864 416102 2916
rect 418157 2907 418215 2913
rect 418157 2873 418169 2907
rect 418203 2904 418215 2907
rect 426713 2907 426771 2913
rect 426713 2904 426725 2907
rect 418203 2876 426725 2904
rect 418203 2873 418215 2876
rect 418157 2867 418215 2873
rect 426713 2873 426725 2876
rect 426759 2873 426771 2907
rect 426713 2867 426771 2873
rect 462038 2864 462044 2916
rect 462096 2904 462102 2916
rect 466730 2904 466736 2916
rect 462096 2876 466736 2904
rect 462096 2864 462102 2876
rect 466730 2864 466736 2876
rect 466788 2864 466794 2916
rect 503714 2864 503720 2916
rect 503772 2904 503778 2916
rect 531038 2904 531044 2916
rect 503772 2876 531044 2904
rect 503772 2864 503778 2876
rect 531038 2864 531044 2876
rect 531096 2864 531102 2916
rect 542998 2864 543004 2916
rect 543056 2904 543062 2916
rect 547800 2904 547828 3080
rect 551186 3068 551192 3080
rect 551244 3068 551250 3120
rect 571978 3000 571984 3052
rect 572036 3040 572042 3052
rect 577406 3040 577412 3052
rect 572036 3012 577412 3040
rect 572036 3000 572042 3012
rect 577406 3000 577412 3012
rect 577464 3000 577470 3052
rect 543056 2876 547828 2904
rect 543056 2864 543062 2876
rect 107620 2808 121592 2836
rect 107620 2796 107626 2808
rect 121822 2796 121828 2848
rect 121880 2836 121886 2848
rect 269758 2836 269764 2848
rect 121880 2808 269764 2836
rect 121880 2796 121886 2808
rect 269758 2796 269764 2808
rect 269816 2796 269822 2848
rect 310974 2796 310980 2848
rect 311032 2836 311038 2848
rect 385678 2836 385684 2848
rect 311032 2808 385684 2836
rect 311032 2796 311038 2808
rect 385678 2796 385684 2808
rect 385736 2796 385742 2848
rect 395430 2796 395436 2848
rect 395488 2836 395494 2848
rect 420178 2836 420184 2848
rect 395488 2808 420184 2836
rect 395488 2796 395494 2808
rect 420178 2796 420184 2808
rect 420236 2796 420242 2848
rect 471514 2796 471520 2848
rect 471572 2836 471578 2848
rect 471882 2836 471888 2848
rect 471572 2808 471888 2836
rect 471572 2796 471578 2808
rect 471882 2796 471888 2808
rect 471940 2796 471946 2848
rect 516686 2796 516692 2848
rect 516744 2836 516750 2848
rect 527450 2836 527456 2848
rect 516744 2808 527456 2836
rect 516744 2796 516750 2808
rect 527450 2796 527456 2808
rect 527508 2796 527514 2848
rect 529198 2796 529204 2848
rect 529256 2836 529262 2848
rect 541710 2836 541716 2848
rect 529256 2808 541716 2836
rect 529256 2796 529262 2808
rect 541710 2796 541716 2808
rect 541768 2796 541774 2848
rect 373994 1912 374000 1964
rect 374052 1952 374058 1964
rect 375282 1952 375288 1964
rect 374052 1924 375288 1952
rect 374052 1912 374058 1924
rect 375282 1912 375288 1924
rect 375340 1912 375346 1964
rect 480346 960 480352 1012
rect 480404 1000 480410 1012
rect 481082 1000 481088 1012
rect 480404 972 481088 1000
rect 480404 960 480410 972
rect 481082 960 481088 972
rect 481140 960 481146 1012
rect 345474 688 345480 740
rect 345532 728 345538 740
rect 346302 728 346308 740
rect 345532 700 346308 728
rect 345532 688 345538 700
rect 346302 688 346308 700
rect 346360 688 346366 740
rect 139670 552 139676 604
rect 139728 592 139734 604
rect 140682 592 140688 604
rect 139728 564 140688 592
rect 139728 552 139734 564
rect 140682 552 140688 564
rect 140740 552 140746 604
rect 172974 552 172980 604
rect 173032 592 173038 604
rect 173802 592 173808 604
rect 173032 564 173808 592
rect 173032 552 173038 564
rect 173802 552 173808 564
rect 173860 552 173866 604
rect 180150 552 180156 604
rect 180208 592 180214 604
rect 180702 592 180708 604
rect 180208 564 180708 592
rect 180208 552 180214 564
rect 180702 552 180708 564
rect 180760 552 180766 604
rect 205082 552 205088 604
rect 205140 592 205146 604
rect 205542 592 205548 604
rect 205140 564 205548 592
rect 205140 552 205146 564
rect 205542 552 205548 564
rect 205600 552 205606 604
rect 206278 552 206284 604
rect 206336 592 206342 604
rect 206922 592 206928 604
rect 206336 564 206928 592
rect 206336 552 206342 564
rect 206922 552 206928 564
rect 206980 552 206986 604
rect 220538 552 220544 604
rect 220596 592 220602 604
rect 220722 592 220728 604
rect 220596 564 220728 592
rect 220596 552 220602 564
rect 220722 552 220728 564
rect 220780 552 220786 604
rect 393038 592 393044 604
rect 392999 564 393044 592
rect 393038 552 393044 564
rect 393096 552 393102 604
rect 435818 552 435824 604
rect 435876 592 435882 604
rect 436002 592 436008 604
rect 435876 564 436008 592
rect 435876 552 435882 564
rect 436002 552 436008 564
rect 436060 552 436066 604
rect 453666 552 453672 604
rect 453724 592 453730 604
rect 453942 592 453948 604
rect 453724 564 453948 592
rect 453724 552 453730 564
rect 453942 552 453948 564
rect 454000 552 454006 604
rect 499758 552 499764 604
rect 499816 592 499822 604
rect 500126 592 500132 604
rect 499816 564 500132 592
rect 499816 552 499822 564
rect 500126 552 500132 564
rect 500184 552 500190 604
rect 506658 552 506664 604
rect 506716 592 506722 604
rect 507210 592 507216 604
rect 506716 564 507216 592
rect 506716 552 506722 564
rect 507210 552 507216 564
rect 507268 552 507274 604
rect 513558 552 513564 604
rect 513616 592 513622 604
rect 514386 592 514392 604
rect 513616 564 514392 592
rect 513616 552 513622 564
rect 514386 552 514392 564
rect 514444 552 514450 604
rect 520366 552 520372 604
rect 520424 592 520430 604
rect 521470 592 521476 604
rect 520424 564 521476 592
rect 520424 552 520430 564
rect 521470 552 521476 564
rect 521528 552 521534 604
<< via1 >>
rect 218980 700952 219032 701004
rect 393320 700952 393372 701004
rect 355968 700884 356020 700936
rect 543464 700884 543516 700936
rect 202788 700816 202840 700868
rect 390560 700816 390612 700868
rect 170312 700748 170364 700800
rect 396080 700748 396132 700800
rect 154120 700680 154172 700732
rect 401600 700680 401652 700732
rect 137836 700612 137888 700664
rect 398840 700612 398892 700664
rect 105452 700544 105504 700596
rect 404360 700544 404412 700596
rect 89168 700476 89220 700528
rect 409880 700476 409932 700528
rect 72976 700408 73028 700460
rect 407120 700408 407172 700460
rect 40500 700340 40552 700392
rect 411260 700340 411312 700392
rect 24308 700272 24360 700324
rect 416780 700272 416832 700324
rect 353208 700204 353260 700256
rect 527180 700204 527232 700256
rect 267648 700136 267700 700188
rect 383660 700136 383712 700188
rect 362868 700068 362920 700120
rect 478512 700068 478564 700120
rect 360108 700000 360160 700052
rect 462320 700000 462372 700052
rect 283840 699932 283892 699984
rect 385040 699932 385092 699984
rect 332508 699864 332560 699916
rect 375380 699864 375432 699916
rect 371148 699796 371200 699848
rect 413652 699796 413704 699848
rect 348792 699728 348844 699780
rect 378140 699728 378192 699780
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 364984 699660 365036 699712
rect 365628 699660 365680 699712
rect 368388 699660 368440 699712
rect 397460 699660 397512 699712
rect 344928 696940 344980 696992
rect 580172 696940 580224 696992
rect 429384 688576 429436 688628
rect 429844 688576 429896 688628
rect 559104 688576 559156 688628
rect 559656 688576 559708 688628
rect 347688 685856 347740 685908
rect 580172 685856 580224 685908
rect 429292 684428 429344 684480
rect 559012 684428 559064 684480
rect 3516 681708 3568 681760
rect 419540 681708 419592 681760
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 342168 673480 342220 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 425060 667904 425112 667956
rect 429660 666544 429712 666596
rect 494152 666544 494204 666596
rect 559380 666544 559432 666596
rect 429476 656863 429528 656872
rect 429476 656829 429485 656863
rect 429485 656829 429519 656863
rect 429519 656829 429528 656863
rect 429476 656820 429528 656829
rect 559196 656863 559248 656872
rect 559196 656829 559205 656863
rect 559205 656829 559239 656863
rect 559239 656829 559248 656863
rect 559196 656820 559248 656829
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 422300 652740 422352 652792
rect 336648 650020 336700 650072
rect 580172 650020 580224 650072
rect 429568 647232 429620 647284
rect 559288 647232 559340 647284
rect 365168 643968 365220 644020
rect 429568 643968 429620 644020
rect 300768 643900 300820 643952
rect 380992 643900 381044 643952
rect 357348 643832 357400 643884
rect 494244 643832 494296 643884
rect 235908 643764 235960 643816
rect 388904 643764 388956 643816
rect 349436 643696 349488 643748
rect 559288 643696 559340 643748
rect 365628 643084 365680 643136
rect 373080 643084 373132 643136
rect 331036 643016 331088 643068
rect 530400 643016 530452 643068
rect 323124 642948 323176 643000
rect 531228 642948 531280 643000
rect 315212 642880 315264 642932
rect 531044 642880 531096 642932
rect 296812 642812 296864 642864
rect 530768 642812 530820 642864
rect 309968 642744 310020 642796
rect 580172 642744 580224 642796
rect 270500 642676 270552 642728
rect 580448 642676 580500 642728
rect 5448 642608 5500 642660
rect 433616 642608 433668 642660
rect 5356 642540 5408 642592
rect 441528 642540 441580 642592
rect 3240 642472 3292 642524
rect 438860 642472 438912 642524
rect 8024 642404 8076 642456
rect 446772 642404 446824 642456
rect 5172 642336 5224 642388
rect 449440 642336 449492 642388
rect 7932 642268 7984 642320
rect 454684 642268 454736 642320
rect 3332 642200 3384 642252
rect 459928 642200 459980 642252
rect 6368 642132 6420 642184
rect 465172 642132 465224 642184
rect 4988 642064 5040 642116
rect 470508 642064 470560 642116
rect 6276 641996 6328 642048
rect 480996 641996 481048 642048
rect 4068 641928 4120 641980
rect 486240 641928 486292 641980
rect 3976 641860 4028 641912
rect 496820 641860 496872 641912
rect 3884 641792 3936 641844
rect 502064 641792 502116 641844
rect 3792 641724 3844 641776
rect 512552 641724 512604 641776
rect 320456 641112 320508 641164
rect 530492 641112 530544 641164
rect 312544 641044 312596 641096
rect 531136 641044 531188 641096
rect 302056 640976 302108 641028
rect 530860 640976 530912 641028
rect 294144 640908 294196 640960
rect 529572 640908 529624 640960
rect 286232 640840 286284 640892
rect 529480 640840 529532 640892
rect 278320 640772 278372 640824
rect 530584 640772 530636 640824
rect 265164 640704 265216 640756
rect 580356 640704 580408 640756
rect 7840 640636 7892 640688
rect 467840 640636 467892 640688
rect 7748 640568 7800 640620
rect 475752 640568 475804 640620
rect 4804 640500 4856 640552
rect 499396 640500 499448 640552
rect 6184 640432 6236 640484
rect 507308 640432 507360 640484
rect 7656 640364 7708 640416
rect 515220 640364 515272 640416
rect 7564 640296 7616 640348
rect 523132 640296 523184 640348
rect 428096 639931 428148 639940
rect 428096 639897 428105 639931
rect 428105 639897 428139 639931
rect 428139 639897 428148 639931
rect 428096 639888 428148 639897
rect 436100 639931 436152 639940
rect 436100 639897 436109 639931
rect 436109 639897 436143 639931
rect 436143 639897 436152 639931
rect 436100 639888 436152 639897
rect 443828 639931 443880 639940
rect 443828 639897 443837 639931
rect 443837 639897 443871 639931
rect 443871 639897 443880 639931
rect 443828 639888 443880 639897
rect 451740 639931 451792 639940
rect 451740 639897 451749 639931
rect 451749 639897 451783 639931
rect 451783 639897 451792 639931
rect 451740 639888 451792 639897
rect 520280 639931 520332 639940
rect 520280 639897 520289 639931
rect 520289 639897 520323 639931
rect 520323 639897 520332 639931
rect 520280 639888 520332 639897
rect 333888 639820 333940 639872
rect 529756 639820 529808 639872
rect 325976 639752 326028 639804
rect 529664 639752 529716 639804
rect 328460 639684 328512 639736
rect 338028 639684 338080 639736
rect 339224 639684 339276 639736
rect 579804 639684 579856 639736
rect 307576 639616 307628 639668
rect 580908 639616 580960 639668
rect 299480 639548 299532 639600
rect 580816 639548 580868 639600
rect 291752 639480 291804 639532
rect 580724 639480 580776 639532
rect 284024 639412 284076 639464
rect 580632 639412 580684 639464
rect 275928 639344 275980 639396
rect 580540 639344 580592 639396
rect 268200 639276 268252 639328
rect 580264 639276 580316 639328
rect 6736 639208 6788 639260
rect 6644 639140 6696 639192
rect 6552 639072 6604 639124
rect 6460 639004 6512 639056
rect 3608 638936 3660 638988
rect 529756 627852 529808 627904
rect 580080 627852 580132 627904
rect 3148 624928 3200 624980
rect 6736 624928 6788 624980
rect 2780 610512 2832 610564
rect 5448 610512 5500 610564
rect 530308 604392 530360 604444
rect 580080 604392 580132 604444
rect 3148 596028 3200 596080
rect 8116 596028 8168 596080
rect 530400 593308 530452 593360
rect 580080 593308 580132 593360
rect 529664 580932 529716 580984
rect 580080 580932 580132 580984
rect 3148 567536 3200 567588
rect 6644 567536 6696 567588
rect 530492 557472 530544 557524
rect 580080 557472 580132 557524
rect 2780 553052 2832 553104
rect 5356 553052 5408 553104
rect 531228 546388 531280 546440
rect 580080 546388 580132 546440
rect 531136 510552 531188 510604
rect 580080 510552 580132 510604
rect 3240 510348 3292 510400
rect 6552 510348 6604 510400
rect 531044 499468 531096 499520
rect 580080 499468 580132 499520
rect 2780 496408 2832 496460
rect 5172 496408 5224 496460
rect 3240 481244 3292 481296
rect 8024 481244 8076 481296
rect 530952 463632 531004 463684
rect 579804 463632 579856 463684
rect 3148 452412 3200 452464
rect 6460 452412 6512 452464
rect 530860 440172 530912 440224
rect 580172 440172 580224 440224
rect 2780 437996 2832 438048
rect 5264 437996 5316 438048
rect 3240 424260 3292 424312
rect 7932 424260 7984 424312
rect 530768 416712 530820 416764
rect 580172 416712 580224 416764
rect 529572 393252 529624 393304
rect 579620 393252 579672 393304
rect 3240 380604 3292 380656
rect 6368 380604 6420 380656
rect 2780 366732 2832 366784
rect 5080 366732 5132 366784
rect 529664 346332 529716 346384
rect 580172 346332 580224 346384
rect 356704 338376 356756 338428
rect 357348 338376 357400 338428
rect 71044 338036 71096 338088
rect 264888 338036 264940 338088
rect 332508 338036 332560 338088
rect 400220 338036 400272 338088
rect 412088 338036 412140 338088
rect 419172 338036 419224 338088
rect 420276 338036 420328 338088
rect 445484 338036 445536 338088
rect 512276 338036 512328 338088
rect 547144 338036 547196 338088
rect 66904 337968 66956 338020
rect 261208 337968 261260 338020
rect 322756 337968 322808 338020
rect 395252 337968 395304 338020
rect 402612 337968 402664 338020
rect 416688 337968 416740 338020
rect 443644 337968 443696 338020
rect 451924 337968 451976 338020
rect 459008 337968 459060 338020
rect 490840 337968 490892 338020
rect 512828 337968 512880 338020
rect 547236 337968 547288 338020
rect 57244 337900 57296 337952
rect 257528 337900 257580 337952
rect 309784 337900 309836 337952
rect 50344 337832 50396 337884
rect 251364 337832 251416 337884
rect 268384 337832 268436 337884
rect 288716 337832 288768 337884
rect 311900 337832 311952 337884
rect 312268 337832 312320 337884
rect 313464 337832 313516 337884
rect 314108 337832 314160 337884
rect 314660 337832 314712 337884
rect 315396 337832 315448 337884
rect 316040 337900 316092 337952
rect 316684 337900 316736 337952
rect 317604 337900 317656 337952
rect 318340 337900 318392 337952
rect 320180 337900 320232 337952
rect 320916 337900 320968 337952
rect 385684 337900 385736 337952
rect 389732 337900 389784 337952
rect 387984 337832 388036 337884
rect 407764 337900 407816 337952
rect 415492 337900 415544 337952
rect 391204 337832 391256 337884
rect 397092 337832 397144 337884
rect 405004 337832 405056 337884
rect 411812 337832 411864 337884
rect 413284 337832 413336 337884
rect 420368 337900 420420 337952
rect 439964 337900 440016 337952
rect 442264 337900 442316 337952
rect 449808 337900 449860 337952
rect 453396 337900 453448 337952
rect 462044 337900 462096 337952
rect 490196 337900 490248 337952
rect 501604 337900 501656 337952
rect 503444 337900 503496 337952
rect 503628 337900 503680 337952
rect 520832 337900 520884 337952
rect 556804 337900 556856 337952
rect 416136 337832 416188 337884
rect 443000 337832 443052 337884
rect 449256 337832 449308 337884
rect 457168 337832 457220 337884
rect 497556 337832 497608 337884
rect 509884 337832 509936 337884
rect 514668 337832 514720 337884
rect 553400 337832 553452 337884
rect 46204 337764 46256 337816
rect 247684 337764 247736 337816
rect 269764 337764 269816 337816
rect 292396 337764 292448 337816
rect 294604 337764 294656 337816
rect 375104 337764 375156 337816
rect 376024 337764 376076 337816
rect 406292 337764 406344 337816
rect 409788 337764 409840 337816
rect 436928 337764 436980 337816
rect 437480 337764 437532 337816
rect 438768 337764 438820 337816
rect 445024 337764 445076 337816
rect 456524 337764 456576 337816
rect 463608 337764 463660 337816
rect 468116 337764 468168 337816
rect 489000 337764 489052 337816
rect 502616 337764 502668 337816
rect 504272 337764 504324 337816
rect 505008 337764 505060 337816
rect 39304 337696 39356 337748
rect 240416 337696 240468 337748
rect 258724 337696 258776 337748
rect 266728 337696 266780 337748
rect 287704 337696 287756 337748
rect 369584 337696 369636 337748
rect 374644 337696 374696 337748
rect 409972 337696 410024 337748
rect 412548 337696 412600 337748
rect 441804 337696 441856 337748
rect 442356 337696 442408 337748
rect 454684 337696 454736 337748
rect 487160 337696 487212 337748
rect 499764 337696 499816 337748
rect 499948 337696 500000 337748
rect 500868 337696 500920 337748
rect 501236 337696 501288 337748
rect 505468 337696 505520 337748
rect 506388 337696 506440 337748
rect 507952 337764 508004 337816
rect 509148 337764 509200 337816
rect 515864 337764 515916 337816
rect 554872 337764 554924 337816
rect 32404 337628 32456 337680
rect 253388 337628 253440 337680
rect 255688 337628 255740 337680
rect 264336 337628 264388 337680
rect 281448 337628 281500 337680
rect 283564 337628 283616 337680
rect 365904 337628 365956 337680
rect 366916 337628 366968 337680
rect 418528 337628 418580 337680
rect 420828 337628 420880 337680
rect 446128 337628 446180 337680
rect 456064 337628 456116 337680
rect 463884 337628 463936 337680
rect 466368 337628 466420 337680
rect 469404 337628 469456 337680
rect 475476 337628 475528 337680
rect 477684 337628 477736 337680
rect 485872 337628 485924 337680
rect 489184 337628 489236 337680
rect 491392 337628 491444 337680
rect 492496 337628 492548 337680
rect 495072 337628 495124 337680
rect 496084 337628 496136 337680
rect 496912 337628 496964 337680
rect 498844 337628 498896 337680
rect 28264 337560 28316 337612
rect 3332 337492 3384 337544
rect 7840 337492 7892 337544
rect 17224 337492 17276 337544
rect 228180 337492 228232 337544
rect 234896 337492 234948 337544
rect 248328 337560 248380 337612
rect 244648 337492 244700 337544
rect 246304 337492 246356 337544
rect 290004 337560 290056 337612
rect 293868 337560 293920 337612
rect 380624 337560 380676 337612
rect 391572 337560 391624 337612
rect 393228 337560 393280 337612
rect 432052 337560 432104 337612
rect 441252 337560 441304 337612
rect 452844 337560 452896 337612
rect 453948 337560 454000 337612
rect 463240 337560 463292 337612
rect 492680 337560 492732 337612
rect 510804 337628 510856 337680
rect 518348 337696 518400 337748
rect 560300 337696 560352 337748
rect 516784 337628 516836 337680
rect 502432 337560 502484 337612
rect 503536 337560 503588 337612
rect 508596 337560 508648 337612
rect 526904 337628 526956 337680
rect 262864 337492 262916 337544
rect 285036 337492 285088 337544
rect 286968 337492 287020 337544
rect 376944 337492 376996 337544
rect 384028 337492 384080 337544
rect 389088 337492 389140 337544
rect 24124 337424 24176 337476
rect 15844 337356 15896 337408
rect 228180 337356 228232 337408
rect 235448 337356 235500 337408
rect 261484 337424 261536 337476
rect 239772 337356 239824 337408
rect 257344 337356 257396 337408
rect 263048 337356 263100 337408
rect 61384 337288 61436 337340
rect 251732 337288 251784 337340
rect 251824 337288 251876 337340
rect 253204 337288 253256 337340
rect 255964 337288 256016 337340
rect 259368 337288 259420 337340
rect 264244 337424 264296 337476
rect 279608 337424 279660 337476
rect 280068 337424 280120 337476
rect 373264 337424 373316 337476
rect 375288 337424 375340 337476
rect 422208 337424 422260 337476
rect 275928 337356 275980 337408
rect 276664 337356 276716 337408
rect 371424 337356 371476 337408
rect 372528 337356 372580 337408
rect 421012 337356 421064 337408
rect 432604 337492 432656 337544
rect 435732 337492 435784 337544
rect 451004 337492 451056 337544
rect 451188 337492 451240 337544
rect 461400 337492 461452 337544
rect 479800 337492 479852 337544
rect 485964 337492 486016 337544
rect 494520 337492 494572 337544
rect 513564 337492 513616 337544
rect 528928 337492 528980 337544
rect 563152 337628 563204 337680
rect 529388 337560 529440 337612
rect 573364 337560 573416 337612
rect 446404 337424 446456 337476
rect 446496 337424 446548 337476
rect 458364 337424 458416 337476
rect 485320 337424 485372 337476
rect 493324 337424 493376 337476
rect 496268 337424 496320 337476
rect 429568 337356 429620 337408
rect 447324 337356 447376 337408
rect 453304 337356 453356 337408
rect 460756 337356 460808 337408
rect 460848 337356 460900 337408
rect 466920 337356 466972 337408
rect 482836 337356 482888 337408
rect 491484 337356 491536 337408
rect 510988 337424 511040 337476
rect 511816 337424 511868 337476
rect 515312 337424 515364 337476
rect 517612 337356 517664 337408
rect 519544 337424 519596 337476
rect 567200 337492 567252 337544
rect 529480 337424 529532 337476
rect 569224 337424 569276 337476
rect 531320 337356 531372 337408
rect 571984 337356 572036 337408
rect 270408 337288 270460 337340
rect 284944 337288 284996 337340
rect 338948 337288 339000 337340
rect 403900 337288 403952 337340
rect 411168 337288 411220 337340
rect 84844 337220 84896 337272
rect 272248 337220 272300 337272
rect 283656 337220 283708 337272
rect 337108 337220 337160 337272
rect 339408 337220 339460 337272
rect 97264 337152 97316 337204
rect 277768 337152 277820 337204
rect 316684 337152 316736 337204
rect 346308 337220 346360 337272
rect 407488 337220 407540 337272
rect 409144 337220 409196 337272
rect 428372 337288 428424 337340
rect 428556 337288 428608 337340
rect 450360 337288 450412 337340
rect 506664 337288 506716 337340
rect 413468 337220 413520 337272
rect 104808 337084 104860 337136
rect 283196 337084 283248 337136
rect 353208 337084 353260 337136
rect 417608 337152 417660 337204
rect 422208 337220 422260 337272
rect 424968 337220 425020 337272
rect 447968 337220 448020 337272
rect 448428 337220 448480 337272
rect 460204 337220 460256 337272
rect 495716 337220 495768 337272
rect 496728 337220 496780 337272
rect 506756 337220 506808 337272
rect 507768 337220 507820 337272
rect 424048 337152 424100 337204
rect 433248 337152 433300 337204
rect 449164 337152 449216 337204
rect 498108 337152 498160 337204
rect 520372 337288 520424 337340
rect 517152 337220 517204 337272
rect 549904 337288 549956 337340
rect 522028 337220 522080 337272
rect 558184 337220 558236 337272
rect 509056 337152 509108 337204
rect 540244 337152 540296 337204
rect 357348 337084 357400 337136
rect 413652 337084 413704 337136
rect 414664 337084 414716 337136
rect 422852 337084 422904 337136
rect 423588 337084 423640 337136
rect 111708 337016 111760 337068
rect 286876 337016 286928 337068
rect 360108 337016 360160 337068
rect 414848 337016 414900 337068
rect 420184 337016 420236 337068
rect 431868 337016 431920 337068
rect 451648 337084 451700 337136
rect 507308 337084 507360 337136
rect 538220 337084 538272 337136
rect 118608 336948 118660 337000
rect 290556 336948 290608 337000
rect 366456 336948 366508 337000
rect 417332 336948 417384 337000
rect 424416 336948 424468 337000
rect 431224 336948 431276 337000
rect 125508 336880 125560 336932
rect 294236 336880 294288 336932
rect 366364 336880 366416 336932
rect 395436 336880 395488 336932
rect 400772 336880 400824 336932
rect 413376 336880 413428 336932
rect 427084 336880 427136 336932
rect 436008 337016 436060 337068
rect 454040 337016 454092 337068
rect 482192 337016 482244 337068
rect 482836 337016 482888 337068
rect 509792 337016 509844 337068
rect 540336 337016 540388 337068
rect 434628 336948 434680 337000
rect 464344 336948 464396 337000
rect 466276 336948 466328 337000
rect 479156 336948 479208 337000
rect 484584 336948 484636 337000
rect 516508 336948 516560 337000
rect 517428 336948 517480 337000
rect 517704 336948 517756 337000
rect 518808 336948 518860 337000
rect 518992 336948 519044 337000
rect 520096 336948 520148 337000
rect 545764 336948 545816 337000
rect 440608 336880 440660 336932
rect 105544 336812 105596 336864
rect 274088 336812 274140 336864
rect 363604 336812 363656 336864
rect 398932 336812 398984 336864
rect 106924 336744 106976 336796
rect 268568 336744 268620 336796
rect 347964 336744 348016 336796
rect 348792 336744 348844 336796
rect 363696 336744 363748 336796
rect 356520 336676 356572 336728
rect 356704 336676 356756 336728
rect 381544 336744 381596 336796
rect 382464 336744 382516 336796
rect 382924 336744 382976 336796
rect 386144 336744 386196 336796
rect 389916 336744 389968 336796
rect 393412 336744 393464 336796
rect 396724 336744 396776 336796
rect 404452 336812 404504 336864
rect 410616 336812 410668 336864
rect 416412 336812 416464 336864
rect 427728 336812 427780 336864
rect 429108 336812 429160 336864
rect 435364 336812 435416 336864
rect 442448 336812 442500 336864
rect 401048 336744 401100 336796
rect 408132 336744 408184 336796
rect 410524 336744 410576 336796
rect 413008 336744 413060 336796
rect 416044 336744 416096 336796
rect 424232 336744 424284 336796
rect 424324 336744 424376 336796
rect 425888 336744 425940 336796
rect 430488 336744 430540 336796
rect 437480 336744 437532 336796
rect 438124 336744 438176 336796
rect 444288 336744 444340 336796
rect 446404 336744 446456 336796
rect 453488 336880 453540 336932
rect 462964 336880 463016 336932
rect 464436 336880 464488 336932
rect 464988 336812 465040 336864
rect 468760 336880 468812 336932
rect 476764 336880 476816 336932
rect 477408 336880 477460 336932
rect 478512 336880 478564 336932
rect 483204 336880 483256 336932
rect 498752 336880 498804 336932
rect 499488 336880 499540 336932
rect 504916 336880 504968 336932
rect 534080 336880 534132 336932
rect 467748 336812 467800 336864
rect 469956 336812 470008 336864
rect 480996 336812 481048 336864
rect 485044 336812 485096 336864
rect 513472 336812 513524 336864
rect 543004 336812 543056 336864
rect 447784 336744 447836 336796
rect 455328 336744 455380 336796
rect 460204 336744 460256 336796
rect 462596 336744 462648 336796
rect 464436 336744 464488 336796
rect 465724 336744 465776 336796
rect 469864 336744 469916 336796
rect 471244 336744 471296 336796
rect 474924 336744 474976 336796
rect 476028 336744 476080 336796
rect 476120 336744 476172 336796
rect 477592 336744 477644 336796
rect 477960 336744 478012 336796
rect 478788 336744 478840 336796
rect 480352 336744 480404 336796
rect 481548 336744 481600 336796
rect 481640 336744 481692 336796
rect 482928 336744 482980 336796
rect 483480 336744 483532 336796
rect 484308 336744 484360 336796
rect 484676 336744 484728 336796
rect 485688 336744 485740 336796
rect 503444 336744 503496 336796
rect 524512 336744 524564 336796
rect 525616 336744 525668 336796
rect 526352 336744 526404 336796
rect 382648 336676 382700 336728
rect 527548 336744 527600 336796
rect 528468 336744 528520 336796
rect 528744 336744 528796 336796
rect 529848 336744 529900 336796
rect 382464 336608 382516 336660
rect 230664 335588 230716 335640
rect 231492 335588 231544 335640
rect 237472 335588 237524 335640
rect 238300 335588 238352 335640
rect 241520 335588 241572 335640
rect 241980 335588 242032 335640
rect 243084 335588 243136 335640
rect 243820 335588 243872 335640
rect 245660 335588 245712 335640
rect 246212 335588 246264 335640
rect 248420 335588 248472 335640
rect 249156 335588 249208 335640
rect 302332 335588 302384 335640
rect 303068 335588 303120 335640
rect 303620 335588 303672 335640
rect 304356 335588 304408 335640
rect 307852 335588 307904 335640
rect 308036 335588 308088 335640
rect 310704 335588 310756 335640
rect 311164 335588 311216 335640
rect 323124 335588 323176 335640
rect 323860 335588 323912 335640
rect 325700 335588 325752 335640
rect 326436 335588 326488 335640
rect 328644 335588 328696 335640
rect 329380 335588 329432 335640
rect 335360 335588 335412 335640
rect 336188 335588 336240 335640
rect 340880 335588 340932 335640
rect 341708 335588 341760 335640
rect 345020 335588 345072 335640
rect 345940 335588 345992 335640
rect 349160 335588 349212 335640
rect 349620 335588 349672 335640
rect 350540 335588 350592 335640
rect 351460 335588 351512 335640
rect 354680 335588 354732 335640
rect 355140 335588 355192 335640
rect 357624 335588 357676 335640
rect 358268 335588 358320 335640
rect 360200 335588 360252 335640
rect 360660 335588 360712 335640
rect 361672 335588 361724 335640
rect 362500 335588 362552 335640
rect 362960 335588 363012 335640
rect 363788 335588 363840 335640
rect 377036 335631 377088 335640
rect 377036 335597 377045 335631
rect 377045 335597 377079 335631
rect 377079 335597 377088 335631
rect 377036 335588 377088 335597
rect 378232 335588 378284 335640
rect 379060 335588 379112 335640
rect 405924 335588 405976 335640
rect 406660 335588 406712 335640
rect 422300 335588 422352 335640
rect 423220 335588 423272 335640
rect 430580 335588 430632 335640
rect 431132 335588 431184 335640
rect 334072 335384 334124 335436
rect 318984 335316 319036 335368
rect 319628 335316 319680 335368
rect 294512 335248 294564 335300
rect 356520 335291 356572 335300
rect 356520 335257 356529 335291
rect 356529 335257 356563 335291
rect 356563 335257 356572 335291
rect 356520 335248 356572 335257
rect 334164 335180 334216 335232
rect 252744 334568 252796 334620
rect 253296 334568 253348 334620
rect 296812 334432 296864 334484
rect 297548 334432 297600 334484
rect 428004 334296 428056 334348
rect 428464 334296 428516 334348
rect 299480 333888 299532 333940
rect 300124 333888 300176 333940
rect 259644 333276 259696 333328
rect 260288 333276 260340 333328
rect 352012 333276 352064 333328
rect 352656 333276 352708 333328
rect 466552 333276 466604 333328
rect 467104 333276 467156 333328
rect 339500 333208 339552 333260
rect 340420 333208 340472 333260
rect 343640 332188 343692 332240
rect 344100 332188 344152 332240
rect 306380 331916 306432 331968
rect 306748 331916 306800 331968
rect 324412 331848 324464 331900
rect 325056 331848 325108 331900
rect 327264 331848 327316 331900
rect 327448 331848 327500 331900
rect 333980 331576 334032 331628
rect 334256 331576 334308 331628
rect 295800 331236 295852 331288
rect 295616 331168 295668 331220
rect 305184 331168 305236 331220
rect 416780 331168 416832 331220
rect 416964 331168 417016 331220
rect 422300 331168 422352 331220
rect 422484 331168 422536 331220
rect 305276 331100 305328 331152
rect 381176 331143 381228 331152
rect 381176 331109 381185 331143
rect 381185 331109 381219 331143
rect 381219 331109 381228 331143
rect 381176 331100 381228 331109
rect 254216 330420 254268 330472
rect 254768 330420 254820 330472
rect 371516 328516 371568 328568
rect 236276 328448 236328 328500
rect 236920 328448 236972 328500
rect 241796 328448 241848 328500
rect 242348 328448 242400 328500
rect 265256 328448 265308 328500
rect 265624 328448 265676 328500
rect 267096 328448 267148 328500
rect 270776 328448 270828 328500
rect 271144 328448 271196 328500
rect 309416 328448 309468 328500
rect 309692 328448 309744 328500
rect 330024 328448 330076 328500
rect 330576 328448 330628 328500
rect 331496 328448 331548 328500
rect 331680 328448 331732 328500
rect 334440 328448 334492 328500
rect 334808 328448 334860 328500
rect 336924 328448 336976 328500
rect 337200 328448 337252 328500
rect 342628 328448 342680 328500
rect 342996 328448 343048 328500
rect 353576 328448 353628 328500
rect 353944 328448 353996 328500
rect 359096 328448 359148 328500
rect 359464 328448 359516 328500
rect 364616 328448 364668 328500
rect 364800 328448 364852 328500
rect 367284 328448 367336 328500
rect 367836 328448 367888 328500
rect 370136 328448 370188 328500
rect 370320 328448 370372 328500
rect 371332 328448 371384 328500
rect 381084 328448 381136 328500
rect 386696 328448 386748 328500
rect 386880 328448 386932 328500
rect 232228 328380 232280 328432
rect 232320 328380 232372 328432
rect 392308 328423 392360 328432
rect 392308 328389 392317 328423
rect 392317 328389 392351 328423
rect 392351 328389 392360 328423
rect 392308 328380 392360 328389
rect 393228 328423 393280 328432
rect 393228 328389 393237 328423
rect 393237 328389 393271 328423
rect 393271 328389 393280 328423
rect 393228 328380 393280 328389
rect 397828 328423 397880 328432
rect 397828 328389 397837 328423
rect 397837 328389 397871 328423
rect 397871 328389 397880 328423
rect 397828 328380 397880 328389
rect 400312 328380 400364 328432
rect 400588 328380 400640 328432
rect 416964 328380 417016 328432
rect 422484 328380 422536 328432
rect 428004 328380 428056 328432
rect 433708 328423 433760 328432
rect 433708 328389 433717 328423
rect 433717 328389 433751 328423
rect 433751 328389 433760 328423
rect 433708 328380 433760 328389
rect 472164 328380 472216 328432
rect 377036 327131 377088 327140
rect 377036 327097 377045 327131
rect 377045 327097 377079 327131
rect 377079 327097 377088 327131
rect 377036 327088 377088 327097
rect 477316 327088 477368 327140
rect 480352 327088 480404 327140
rect 281632 327020 281684 327072
rect 282000 327020 282052 327072
rect 292764 327063 292816 327072
rect 292764 327029 292773 327063
rect 292773 327029 292807 327063
rect 292807 327029 292816 327063
rect 292764 327020 292816 327029
rect 357624 327020 357676 327072
rect 382464 327063 382516 327072
rect 382464 327029 382473 327063
rect 382473 327029 382507 327063
rect 382507 327029 382516 327063
rect 382464 327020 382516 327029
rect 400312 327063 400364 327072
rect 400312 327029 400321 327063
rect 400321 327029 400355 327063
rect 400355 327029 400364 327063
rect 400312 327020 400364 327029
rect 294052 325703 294104 325712
rect 294052 325669 294061 325703
rect 294061 325669 294095 325703
rect 294095 325669 294104 325703
rect 294052 325660 294104 325669
rect 321652 325660 321704 325712
rect 322112 325660 322164 325712
rect 451372 325660 451424 325712
rect 451556 325660 451608 325712
rect 348056 324300 348108 324352
rect 348240 324300 348292 324352
rect 232320 324275 232372 324284
rect 232320 324241 232329 324275
rect 232329 324241 232363 324275
rect 232363 324241 232372 324275
rect 232320 324232 232372 324241
rect 277308 323552 277360 323604
rect 277584 323552 277636 323604
rect 530676 322872 530728 322924
rect 579620 322872 579672 322924
rect 249984 321691 250036 321700
rect 249984 321657 249993 321691
rect 249993 321657 250027 321691
rect 250027 321657 250036 321691
rect 249984 321648 250036 321657
rect 261024 321648 261076 321700
rect 259644 321623 259696 321632
rect 259644 321589 259653 321623
rect 259653 321589 259687 321623
rect 259687 321589 259696 321623
rect 259644 321580 259696 321589
rect 327264 321580 327316 321632
rect 261024 321512 261076 321564
rect 348056 321580 348108 321632
rect 359096 321580 359148 321632
rect 387984 321580 388036 321632
rect 408684 321580 408736 321632
rect 466552 321623 466604 321632
rect 466552 321589 466561 321623
rect 466561 321589 466595 321623
rect 466595 321589 466604 321623
rect 466552 321580 466604 321589
rect 347964 321512 348016 321564
rect 359004 321512 359056 321564
rect 327264 321444 327316 321496
rect 408776 321444 408828 321496
rect 388076 321376 388128 321428
rect 252744 318860 252796 318912
rect 233424 318792 233476 318844
rect 233516 318792 233568 318844
rect 236276 318792 236328 318844
rect 236368 318792 236420 318844
rect 252560 318792 252612 318844
rect 259644 318835 259696 318844
rect 259644 318801 259653 318835
rect 259653 318801 259687 318835
rect 259687 318801 259696 318835
rect 259644 318792 259696 318801
rect 375564 318792 375616 318844
rect 375748 318792 375800 318844
rect 376944 318792 376996 318844
rect 377036 318792 377088 318844
rect 392400 318792 392452 318844
rect 393228 318835 393280 318844
rect 393228 318801 393237 318835
rect 393237 318801 393271 318835
rect 393271 318801 393280 318835
rect 393228 318792 393280 318801
rect 397920 318792 397972 318844
rect 400496 318792 400548 318844
rect 416872 318835 416924 318844
rect 416872 318801 416881 318835
rect 416881 318801 416915 318835
rect 416915 318801 416924 318835
rect 416872 318792 416924 318801
rect 422392 318835 422444 318844
rect 422392 318801 422401 318835
rect 422401 318801 422435 318835
rect 422435 318801 422444 318835
rect 422392 318792 422444 318801
rect 427912 318835 427964 318844
rect 427912 318801 427921 318835
rect 427921 318801 427955 318835
rect 427955 318801 427964 318835
rect 427912 318792 427964 318801
rect 433800 318792 433852 318844
rect 466552 318835 466604 318844
rect 466552 318801 466561 318835
rect 466561 318801 466595 318835
rect 466595 318801 466604 318835
rect 466552 318792 466604 318801
rect 472072 318835 472124 318844
rect 472072 318801 472081 318835
rect 472081 318801 472115 318835
rect 472115 318801 472124 318835
rect 472072 318792 472124 318801
rect 283012 318724 283064 318776
rect 283104 318724 283156 318776
rect 288624 318767 288676 318776
rect 288624 318733 288633 318767
rect 288633 318733 288667 318767
rect 288667 318733 288676 318767
rect 288624 318724 288676 318733
rect 365812 318724 365864 318776
rect 365904 318724 365956 318776
rect 371332 318724 371384 318776
rect 371424 318724 371476 318776
rect 386696 318767 386748 318776
rect 386696 318733 386705 318767
rect 386705 318733 386739 318767
rect 386739 318733 386748 318767
rect 386696 318724 386748 318733
rect 382464 317543 382516 317552
rect 382464 317509 382473 317543
rect 382473 317509 382507 317543
rect 382507 317509 382516 317543
rect 382464 317500 382516 317509
rect 249984 317475 250036 317484
rect 249984 317441 249993 317475
rect 249993 317441 250027 317475
rect 250027 317441 250036 317475
rect 249984 317432 250036 317441
rect 292764 317475 292816 317484
rect 292764 317441 292773 317475
rect 292773 317441 292807 317475
rect 292807 317441 292816 317475
rect 292764 317432 292816 317441
rect 334440 317432 334492 317484
rect 334532 317432 334584 317484
rect 356520 317475 356572 317484
rect 356520 317441 356529 317475
rect 356529 317441 356563 317475
rect 356563 317441 356572 317475
rect 356520 317432 356572 317441
rect 357532 317475 357584 317484
rect 357532 317441 357541 317475
rect 357541 317441 357575 317475
rect 357575 317441 357584 317475
rect 357532 317432 357584 317441
rect 255412 317364 255464 317416
rect 281632 317407 281684 317416
rect 281632 317373 281641 317407
rect 281641 317373 281675 317407
rect 281675 317373 281684 317407
rect 281632 317364 281684 317373
rect 283012 317407 283064 317416
rect 283012 317373 283021 317407
rect 283021 317373 283055 317407
rect 283055 317373 283064 317407
rect 283012 317364 283064 317373
rect 327264 317364 327316 317416
rect 332692 317364 332744 317416
rect 332876 317364 332928 317416
rect 365812 317364 365864 317416
rect 365904 317364 365956 317416
rect 371332 317407 371384 317416
rect 371332 317373 371341 317407
rect 371341 317373 371375 317407
rect 371375 317373 371384 317407
rect 371332 317364 371384 317373
rect 376944 317407 376996 317416
rect 376944 317373 376953 317407
rect 376953 317373 376987 317407
rect 376987 317373 376996 317407
rect 376944 317364 376996 317373
rect 381084 317364 381136 317416
rect 381360 317364 381412 317416
rect 382464 317407 382516 317416
rect 382464 317373 382473 317407
rect 382473 317373 382507 317407
rect 382507 317373 382516 317407
rect 382464 317364 382516 317373
rect 480352 317407 480404 317416
rect 480352 317373 480361 317407
rect 480361 317373 480395 317407
rect 480395 317373 480404 317407
rect 480352 317364 480404 317373
rect 255688 317296 255740 317348
rect 327264 317228 327316 317280
rect 451556 316072 451608 316124
rect 451740 316072 451792 316124
rect 294144 316004 294196 316056
rect 294328 316004 294380 316056
rect 321468 316004 321520 316056
rect 321744 316004 321796 316056
rect 352104 316004 352156 316056
rect 352288 316004 352340 316056
rect 255688 315936 255740 315988
rect 400496 315979 400548 315988
rect 400496 315945 400505 315979
rect 400505 315945 400539 315979
rect 400539 315945 400548 315979
rect 400496 315936 400548 315945
rect 408776 315979 408828 315988
rect 408776 315945 408785 315979
rect 408785 315945 408819 315979
rect 408819 315945 408828 315979
rect 408776 315936 408828 315945
rect 451556 315979 451608 315988
rect 451556 315945 451565 315979
rect 451565 315945 451599 315979
rect 451599 315945 451608 315979
rect 451556 315936 451608 315945
rect 232412 314644 232464 314696
rect 232320 313259 232372 313268
rect 232320 313225 232329 313259
rect 232329 313225 232363 313259
rect 232363 313225 232372 313259
rect 232320 313216 232372 313225
rect 249892 312536 249944 312588
rect 250076 312536 250128 312588
rect 277584 311967 277636 311976
rect 277584 311933 277593 311967
rect 277593 311933 277627 311967
rect 277627 311933 277636 311967
rect 277584 311924 277636 311933
rect 294144 311924 294196 311976
rect 397552 311856 397604 311908
rect 397920 311856 397972 311908
rect 433432 311856 433484 311908
rect 433800 311856 433852 311908
rect 294144 311788 294196 311840
rect 318892 311788 318944 311840
rect 319076 311788 319128 311840
rect 346584 311831 346636 311840
rect 346584 311797 346593 311831
rect 346593 311797 346627 311831
rect 346627 311797 346636 311831
rect 346584 311788 346636 311797
rect 416780 311788 416832 311840
rect 416964 311788 417016 311840
rect 422300 311788 422352 311840
rect 422484 311788 422536 311840
rect 427820 311788 427872 311840
rect 428004 311788 428056 311840
rect 466460 311788 466512 311840
rect 466644 311788 466696 311840
rect 471980 311788 472032 311840
rect 472164 311788 472216 311840
rect 321468 311176 321520 311228
rect 321744 311176 321796 311228
rect 392032 310904 392084 310956
rect 392492 310904 392544 310956
rect 342628 309204 342680 309256
rect 252560 309136 252612 309188
rect 252744 309136 252796 309188
rect 267096 309179 267148 309188
rect 267096 309145 267105 309179
rect 267105 309145 267139 309179
rect 267139 309145 267148 309179
rect 267096 309136 267148 309145
rect 288624 309179 288676 309188
rect 288624 309145 288633 309179
rect 288633 309145 288667 309179
rect 288667 309145 288676 309179
rect 288624 309136 288676 309145
rect 305184 309136 305236 309188
rect 305276 309136 305328 309188
rect 336832 309136 336884 309188
rect 336924 309136 336976 309188
rect 342444 309136 342496 309188
rect 346584 309179 346636 309188
rect 346584 309145 346593 309179
rect 346593 309145 346627 309179
rect 346627 309145 346636 309179
rect 346584 309136 346636 309145
rect 353484 309136 353536 309188
rect 353576 309136 353628 309188
rect 364524 309136 364576 309188
rect 364616 309136 364668 309188
rect 367376 309136 367428 309188
rect 367468 309136 367520 309188
rect 386696 309179 386748 309188
rect 386696 309145 386705 309179
rect 386705 309145 386739 309179
rect 386739 309145 386748 309179
rect 386696 309136 386748 309145
rect 270684 309111 270736 309120
rect 270684 309077 270693 309111
rect 270693 309077 270727 309111
rect 270727 309077 270736 309111
rect 270684 309068 270736 309077
rect 309324 309111 309376 309120
rect 309324 309077 309333 309111
rect 309333 309077 309367 309111
rect 309367 309077 309376 309111
rect 309324 309068 309376 309077
rect 319076 309068 319128 309120
rect 371332 309111 371384 309120
rect 371332 309077 371341 309111
rect 371341 309077 371375 309111
rect 371375 309077 371384 309111
rect 371332 309068 371384 309077
rect 416964 309068 417016 309120
rect 422484 309111 422536 309120
rect 422484 309077 422493 309111
rect 422493 309077 422527 309111
rect 422527 309077 422536 309111
rect 422484 309068 422536 309077
rect 428004 309111 428056 309120
rect 428004 309077 428013 309111
rect 428013 309077 428047 309111
rect 428047 309077 428056 309111
rect 428004 309068 428056 309077
rect 433432 309111 433484 309120
rect 433432 309077 433441 309111
rect 433441 309077 433475 309111
rect 433475 309077 433484 309111
rect 433432 309068 433484 309077
rect 466644 309068 466696 309120
rect 472164 309068 472216 309120
rect 277492 309000 277544 309052
rect 342444 309043 342496 309052
rect 342444 309009 342453 309043
rect 342453 309009 342487 309043
rect 342487 309009 342496 309043
rect 342444 309000 342496 309009
rect 2780 308796 2832 308848
rect 4988 308796 5040 308848
rect 287152 307844 287204 307896
rect 287336 307844 287388 307896
rect 261024 307776 261076 307828
rect 261116 307776 261168 307828
rect 267096 307819 267148 307828
rect 267096 307785 267105 307819
rect 267105 307785 267139 307819
rect 267139 307785 267148 307819
rect 267096 307776 267148 307785
rect 281632 307819 281684 307828
rect 281632 307785 281641 307819
rect 281641 307785 281675 307819
rect 281675 307785 281684 307819
rect 281632 307776 281684 307785
rect 283012 307819 283064 307828
rect 283012 307785 283021 307819
rect 283021 307785 283055 307819
rect 283055 307785 283064 307819
rect 283012 307776 283064 307785
rect 376944 307819 376996 307828
rect 376944 307785 376953 307819
rect 376953 307785 376987 307819
rect 376987 307785 376996 307819
rect 376944 307776 376996 307785
rect 382464 307819 382516 307828
rect 382464 307785 382473 307819
rect 382473 307785 382507 307819
rect 382507 307785 382516 307819
rect 382464 307776 382516 307785
rect 480352 307819 480404 307828
rect 480352 307785 480361 307819
rect 480361 307785 480395 307819
rect 480395 307785 480404 307819
rect 480352 307776 480404 307785
rect 243084 307708 243136 307760
rect 277584 307751 277636 307760
rect 277584 307717 277593 307751
rect 277593 307717 277627 307751
rect 277627 307717 277636 307751
rect 277584 307708 277636 307717
rect 287336 307708 287388 307760
rect 295524 307751 295576 307760
rect 295524 307717 295533 307751
rect 295533 307717 295567 307751
rect 295567 307717 295576 307751
rect 295524 307708 295576 307717
rect 364524 307751 364576 307760
rect 364524 307717 364533 307751
rect 364533 307717 364567 307751
rect 364567 307717 364576 307751
rect 364524 307708 364576 307717
rect 332692 306416 332744 306468
rect 332876 306416 332928 306468
rect 352104 306348 352156 306400
rect 352288 306348 352340 306400
rect 357532 306348 357584 306400
rect 357716 306348 357768 306400
rect 236368 304920 236420 304972
rect 236552 304920 236604 304972
rect 281632 302268 281684 302320
rect 283012 302268 283064 302320
rect 298284 302268 298336 302320
rect 233332 302200 233384 302252
rect 233516 302200 233568 302252
rect 281816 302064 281868 302116
rect 283104 302064 283156 302116
rect 298376 302064 298428 302116
rect 408776 302107 408828 302116
rect 408776 302073 408785 302107
rect 408785 302073 408819 302107
rect 408819 302073 408828 302107
rect 408776 302064 408828 302073
rect 451556 302107 451608 302116
rect 451556 302073 451565 302107
rect 451565 302073 451599 302107
rect 451599 302073 451608 302107
rect 451556 302064 451608 302073
rect 422484 299931 422536 299940
rect 422484 299897 422493 299931
rect 422493 299897 422527 299931
rect 422527 299897 422536 299931
rect 422484 299888 422536 299897
rect 342536 299548 342588 299600
rect 347964 299548 348016 299600
rect 353484 299548 353536 299600
rect 265164 299480 265216 299532
rect 265256 299480 265308 299532
rect 270776 299480 270828 299532
rect 309416 299480 309468 299532
rect 318984 299523 319036 299532
rect 318984 299489 318993 299523
rect 318993 299489 319027 299523
rect 319027 299489 319036 299523
rect 318984 299480 319036 299489
rect 241796 299455 241848 299464
rect 241796 299421 241805 299455
rect 241805 299421 241839 299455
rect 241839 299421 241848 299455
rect 241796 299412 241848 299421
rect 249984 299455 250036 299464
rect 249984 299421 249993 299455
rect 249993 299421 250027 299455
rect 250027 299421 250036 299455
rect 249984 299412 250036 299421
rect 281816 299412 281868 299464
rect 283104 299455 283156 299464
rect 283104 299421 283113 299455
rect 283113 299421 283147 299455
rect 283147 299421 283156 299455
rect 283104 299412 283156 299421
rect 288624 299455 288676 299464
rect 288624 299421 288633 299455
rect 288633 299421 288667 299455
rect 288667 299421 288676 299455
rect 288624 299412 288676 299421
rect 305184 299455 305236 299464
rect 305184 299421 305193 299455
rect 305193 299421 305227 299455
rect 305227 299421 305236 299455
rect 305184 299412 305236 299421
rect 310704 299455 310756 299464
rect 310704 299421 310713 299455
rect 310713 299421 310747 299455
rect 310747 299421 310756 299455
rect 310704 299412 310756 299421
rect 331404 299412 331456 299464
rect 331496 299412 331548 299464
rect 346584 299455 346636 299464
rect 346584 299421 346593 299455
rect 346593 299421 346627 299455
rect 346627 299421 346636 299455
rect 346584 299412 346636 299421
rect 416872 299523 416924 299532
rect 416872 299489 416881 299523
rect 416881 299489 416915 299523
rect 416915 299489 416924 299523
rect 416872 299480 416924 299489
rect 428004 299523 428056 299532
rect 428004 299489 428013 299523
rect 428013 299489 428047 299523
rect 428047 299489 428056 299523
rect 428004 299480 428056 299489
rect 433708 299480 433760 299532
rect 466552 299523 466604 299532
rect 466552 299489 466561 299523
rect 466561 299489 466595 299523
rect 466595 299489 466604 299523
rect 466552 299480 466604 299489
rect 472072 299523 472124 299532
rect 472072 299489 472081 299523
rect 472081 299489 472115 299523
rect 472115 299489 472124 299523
rect 472072 299480 472124 299489
rect 370044 299412 370096 299464
rect 370136 299412 370188 299464
rect 376944 299455 376996 299464
rect 376944 299421 376953 299455
rect 376953 299421 376987 299455
rect 376987 299421 376996 299455
rect 376944 299412 376996 299421
rect 400496 299455 400548 299464
rect 400496 299421 400505 299455
rect 400505 299421 400539 299455
rect 400539 299421 400548 299455
rect 400496 299412 400548 299421
rect 530584 299412 530636 299464
rect 579712 299412 579764 299464
rect 347964 299344 348016 299396
rect 353484 299344 353536 299396
rect 242992 298231 243044 298240
rect 242992 298197 243001 298231
rect 243001 298197 243035 298231
rect 243035 298197 243044 298231
rect 242992 298188 243044 298197
rect 277584 298231 277636 298240
rect 277584 298197 277593 298231
rect 277593 298197 277627 298231
rect 277627 298197 277636 298231
rect 277584 298188 277636 298197
rect 255504 298163 255556 298172
rect 255504 298129 255513 298163
rect 255513 298129 255547 298163
rect 255547 298129 255556 298163
rect 255504 298120 255556 298129
rect 261024 298120 261076 298172
rect 261208 298120 261260 298172
rect 287244 298163 287296 298172
rect 287244 298129 287253 298163
rect 287253 298129 287287 298163
rect 287287 298129 287296 298163
rect 287244 298120 287296 298129
rect 242992 298095 243044 298104
rect 242992 298061 243001 298095
rect 243001 298061 243035 298095
rect 243035 298061 243044 298095
rect 242992 298052 243044 298061
rect 265256 298052 265308 298104
rect 267096 298052 267148 298104
rect 270776 298052 270828 298104
rect 270868 298052 270920 298104
rect 277584 298095 277636 298104
rect 277584 298061 277593 298095
rect 277593 298061 277627 298095
rect 277627 298061 277636 298095
rect 277584 298052 277636 298061
rect 292764 298052 292816 298104
rect 334256 298163 334308 298172
rect 334256 298129 334265 298163
rect 334265 298129 334299 298163
rect 334299 298129 334308 298163
rect 334256 298120 334308 298129
rect 364616 298120 364668 298172
rect 347964 298095 348016 298104
rect 347964 298061 347973 298095
rect 347973 298061 348007 298095
rect 348007 298061 348016 298095
rect 347964 298052 348016 298061
rect 352104 298095 352156 298104
rect 352104 298061 352113 298095
rect 352113 298061 352147 298095
rect 352147 298061 352156 298095
rect 352104 298052 352156 298061
rect 353484 298052 353536 298104
rect 353576 298052 353628 298104
rect 370044 298095 370096 298104
rect 370044 298061 370053 298095
rect 370053 298061 370087 298095
rect 370087 298061 370096 298095
rect 370044 298052 370096 298061
rect 375472 298095 375524 298104
rect 375472 298061 375481 298095
rect 375481 298061 375515 298095
rect 375515 298061 375524 298095
rect 375472 298052 375524 298061
rect 397736 298095 397788 298104
rect 397736 298061 397745 298095
rect 397745 298061 397779 298095
rect 397779 298061 397788 298095
rect 397736 298052 397788 298061
rect 480352 298095 480404 298104
rect 480352 298061 480361 298095
rect 480361 298061 480395 298095
rect 480395 298061 480404 298095
rect 480352 298052 480404 298061
rect 382464 297984 382516 298036
rect 382556 297984 382608 298036
rect 332784 296692 332836 296744
rect 332968 296692 333020 296744
rect 334256 296735 334308 296744
rect 334256 296701 334265 296735
rect 334265 296701 334299 296735
rect 334299 296701 334308 296735
rect 334256 296692 334308 296701
rect 298376 296667 298428 296676
rect 298376 296633 298385 296667
rect 298385 296633 298419 296667
rect 298419 296633 298428 296667
rect 298376 296624 298428 296633
rect 236276 295264 236328 295316
rect 236460 295264 236512 295316
rect 3332 294924 3384 294976
rect 7748 294924 7800 294976
rect 232320 294899 232372 294908
rect 232320 294865 232329 294899
rect 232329 294865 232363 294899
rect 232363 294865 232372 294899
rect 232320 294856 232372 294865
rect 232320 293904 232372 293956
rect 232412 293904 232464 293956
rect 295708 293224 295760 293276
rect 255504 292612 255556 292664
rect 321744 292612 321796 292664
rect 327264 292612 327316 292664
rect 330024 292612 330076 292664
rect 367376 292612 367428 292664
rect 392216 292544 392268 292596
rect 408776 292612 408828 292664
rect 451556 292612 451608 292664
rect 232412 292519 232464 292528
rect 232412 292485 232421 292519
rect 232421 292485 232455 292519
rect 232455 292485 232464 292519
rect 232412 292476 232464 292485
rect 236460 292519 236512 292528
rect 236460 292485 236469 292519
rect 236469 292485 236503 292519
rect 236503 292485 236512 292519
rect 236460 292476 236512 292485
rect 244464 292476 244516 292528
rect 255504 292476 255556 292528
rect 321744 292476 321796 292528
rect 327264 292476 327316 292528
rect 330024 292476 330076 292528
rect 367376 292476 367428 292528
rect 392124 292476 392176 292528
rect 408684 292476 408736 292528
rect 451464 292476 451516 292528
rect 466460 292476 466512 292528
rect 466644 292476 466696 292528
rect 471980 292476 472032 292528
rect 472164 292476 472216 292528
rect 244464 292340 244516 292392
rect 364524 291363 364576 291372
rect 364524 291329 364533 291363
rect 364533 291329 364567 291363
rect 364567 291329 364576 291363
rect 364524 291320 364576 291329
rect 241796 289867 241848 289876
rect 241796 289833 241805 289867
rect 241805 289833 241839 289867
rect 241839 289833 241848 289867
rect 241796 289824 241848 289833
rect 249984 289867 250036 289876
rect 249984 289833 249993 289867
rect 249993 289833 250027 289867
rect 250027 289833 250036 289867
rect 249984 289824 250036 289833
rect 281632 289867 281684 289876
rect 281632 289833 281641 289867
rect 281641 289833 281675 289867
rect 281675 289833 281684 289867
rect 281632 289824 281684 289833
rect 283104 289867 283156 289876
rect 283104 289833 283113 289867
rect 283113 289833 283147 289867
rect 283147 289833 283156 289867
rect 283104 289824 283156 289833
rect 288624 289867 288676 289876
rect 288624 289833 288633 289867
rect 288633 289833 288667 289867
rect 288667 289833 288676 289867
rect 288624 289824 288676 289833
rect 305184 289867 305236 289876
rect 305184 289833 305193 289867
rect 305193 289833 305227 289867
rect 305227 289833 305236 289867
rect 305184 289824 305236 289833
rect 309324 289824 309376 289876
rect 309600 289824 309652 289876
rect 310704 289867 310756 289876
rect 310704 289833 310713 289867
rect 310713 289833 310747 289867
rect 310747 289833 310756 289867
rect 310704 289824 310756 289833
rect 324504 289824 324556 289876
rect 324688 289824 324740 289876
rect 346584 289867 346636 289876
rect 346584 289833 346593 289867
rect 346593 289833 346627 289867
rect 346627 289833 346636 289867
rect 346584 289824 346636 289833
rect 376944 289867 376996 289876
rect 376944 289833 376953 289867
rect 376953 289833 376987 289867
rect 376987 289833 376996 289867
rect 376944 289824 376996 289833
rect 381084 289824 381136 289876
rect 381360 289824 381412 289876
rect 252744 289799 252796 289808
rect 252744 289765 252753 289799
rect 252753 289765 252787 289799
rect 252787 289765 252796 289799
rect 252744 289756 252796 289765
rect 254124 289799 254176 289808
rect 254124 289765 254133 289799
rect 254133 289765 254167 289799
rect 254167 289765 254176 289799
rect 254124 289756 254176 289765
rect 259644 289799 259696 289808
rect 259644 289765 259653 289799
rect 259653 289765 259687 289799
rect 259687 289765 259696 289799
rect 259644 289756 259696 289765
rect 334256 289799 334308 289808
rect 334256 289765 334265 289799
rect 334265 289765 334299 289799
rect 334299 289765 334308 289799
rect 334256 289756 334308 289765
rect 356428 289756 356480 289808
rect 375472 289799 375524 289808
rect 375472 289765 375481 289799
rect 375481 289765 375515 289799
rect 375515 289765 375524 289799
rect 375472 289756 375524 289765
rect 309324 289731 309376 289740
rect 309324 289697 309333 289731
rect 309333 289697 309367 289731
rect 309367 289697 309376 289731
rect 309324 289688 309376 289697
rect 356520 289688 356572 289740
rect 265164 288439 265216 288448
rect 265164 288405 265173 288439
rect 265173 288405 265207 288439
rect 265207 288405 265216 288439
rect 265164 288396 265216 288405
rect 292672 288439 292724 288448
rect 292672 288405 292681 288439
rect 292681 288405 292715 288439
rect 292715 288405 292724 288439
rect 292672 288396 292724 288405
rect 348056 288396 348108 288448
rect 370044 288439 370096 288448
rect 370044 288405 370053 288439
rect 370053 288405 370087 288439
rect 370087 288405 370096 288439
rect 370044 288396 370096 288405
rect 397736 288439 397788 288448
rect 397736 288405 397745 288439
rect 397745 288405 397779 288439
rect 397779 288405 397788 288439
rect 397736 288396 397788 288405
rect 480352 288439 480404 288448
rect 480352 288405 480361 288439
rect 480361 288405 480395 288439
rect 480395 288405 480404 288439
rect 480352 288396 480404 288405
rect 408684 288371 408736 288380
rect 408684 288337 408693 288371
rect 408693 288337 408727 288371
rect 408727 288337 408736 288371
rect 408684 288328 408736 288337
rect 352104 287963 352156 287972
rect 352104 287929 352113 287963
rect 352113 287929 352147 287963
rect 352147 287929 352156 287963
rect 352104 287920 352156 287929
rect 298468 287036 298520 287088
rect 386604 287079 386656 287088
rect 386604 287045 386613 287079
rect 386613 287045 386647 287079
rect 386647 287045 386656 287079
rect 386604 287036 386656 287045
rect 364616 284928 364668 284980
rect 236460 284359 236512 284368
rect 236460 284325 236469 284359
rect 236469 284325 236503 284359
rect 236503 284325 236512 284359
rect 236460 284316 236512 284325
rect 232412 282931 232464 282940
rect 232412 282897 232421 282931
rect 232421 282897 232455 282931
rect 232455 282897 232464 282931
rect 232412 282888 232464 282897
rect 233332 282888 233384 282940
rect 233516 282888 233568 282940
rect 342536 282931 342588 282940
rect 342536 282897 342545 282931
rect 342545 282897 342579 282931
rect 342579 282897 342588 282931
rect 342536 282888 342588 282897
rect 370044 282888 370096 282940
rect 381084 282888 381136 282940
rect 422300 282888 422352 282940
rect 422484 282888 422536 282940
rect 427820 282888 427872 282940
rect 428004 282888 428056 282940
rect 334440 282752 334492 282804
rect 375472 282820 375524 282872
rect 370136 282752 370188 282804
rect 375656 282752 375708 282804
rect 400496 282820 400548 282872
rect 381176 282752 381228 282804
rect 400496 282684 400548 282736
rect 342536 280279 342588 280288
rect 342536 280245 342545 280279
rect 342545 280245 342579 280279
rect 342579 280245 342588 280279
rect 342536 280236 342588 280245
rect 243176 280168 243228 280220
rect 252744 280211 252796 280220
rect 252744 280177 252753 280211
rect 252753 280177 252787 280211
rect 252787 280177 252796 280211
rect 252744 280168 252796 280177
rect 265072 280168 265124 280220
rect 265256 280168 265308 280220
rect 267004 280211 267056 280220
rect 267004 280177 267013 280211
rect 267013 280177 267047 280211
rect 267047 280177 267056 280211
rect 267004 280168 267056 280177
rect 277676 280168 277728 280220
rect 281724 280168 281776 280220
rect 281908 280168 281960 280220
rect 292672 280168 292724 280220
rect 292764 280168 292816 280220
rect 309416 280168 309468 280220
rect 324412 280168 324464 280220
rect 324688 280168 324740 280220
rect 397460 280168 397512 280220
rect 3148 280100 3200 280152
rect 6276 280100 6328 280152
rect 241796 280143 241848 280152
rect 241796 280109 241805 280143
rect 241805 280109 241839 280143
rect 241839 280109 241848 280143
rect 241796 280100 241848 280109
rect 270592 280100 270644 280152
rect 270868 280100 270920 280152
rect 288624 280143 288676 280152
rect 288624 280109 288633 280143
rect 288633 280109 288667 280143
rect 288667 280109 288676 280143
rect 288624 280100 288676 280109
rect 295432 280100 295484 280152
rect 295708 280100 295760 280152
rect 298468 280100 298520 280152
rect 305184 280143 305236 280152
rect 305184 280109 305193 280143
rect 305193 280109 305227 280143
rect 305227 280109 305236 280143
rect 305184 280100 305236 280109
rect 310704 280143 310756 280152
rect 310704 280109 310713 280143
rect 310713 280109 310747 280143
rect 310747 280109 310756 280143
rect 310704 280100 310756 280109
rect 318984 280100 319036 280152
rect 319076 280100 319128 280152
rect 321744 280143 321796 280152
rect 321744 280109 321753 280143
rect 321753 280109 321787 280143
rect 321787 280109 321796 280143
rect 321744 280100 321796 280109
rect 327264 280143 327316 280152
rect 327264 280109 327273 280143
rect 327273 280109 327307 280143
rect 327307 280109 327316 280143
rect 327264 280100 327316 280109
rect 331404 280100 331456 280152
rect 331496 280100 331548 280152
rect 334440 280100 334492 280152
rect 346584 280143 346636 280152
rect 346584 280109 346593 280143
rect 346593 280109 346627 280143
rect 346627 280109 346636 280143
rect 346584 280100 346636 280109
rect 348056 280100 348108 280152
rect 348148 280100 348200 280152
rect 352104 280100 352156 280152
rect 352288 280100 352340 280152
rect 353484 280100 353536 280152
rect 353576 280100 353628 280152
rect 359004 280100 359056 280152
rect 359096 280100 359148 280152
rect 364524 280100 364576 280152
rect 364616 280100 364668 280152
rect 365904 280100 365956 280152
rect 365996 280100 366048 280152
rect 369768 280100 369820 280152
rect 370136 280100 370188 280152
rect 371424 280100 371476 280152
rect 371516 280100 371568 280152
rect 375196 280100 375248 280152
rect 375656 280100 375708 280152
rect 382464 280143 382516 280152
rect 382464 280109 382473 280143
rect 382473 280109 382507 280143
rect 382507 280109 382516 280143
rect 382464 280100 382516 280109
rect 416872 280143 416924 280152
rect 416872 280109 416881 280143
rect 416881 280109 416915 280143
rect 416915 280109 416924 280143
rect 416872 280100 416924 280109
rect 433616 280143 433668 280152
rect 433616 280109 433625 280143
rect 433625 280109 433659 280143
rect 433659 280109 433668 280143
rect 433616 280100 433668 280109
rect 466552 280143 466604 280152
rect 466552 280109 466561 280143
rect 466561 280109 466595 280143
rect 466595 280109 466604 280143
rect 466552 280100 466604 280109
rect 472072 280143 472124 280152
rect 472072 280109 472081 280143
rect 472081 280109 472115 280143
rect 472115 280109 472124 280143
rect 472072 280100 472124 280109
rect 298284 280032 298336 280084
rect 381176 280032 381228 280084
rect 397460 280032 397512 280084
rect 357624 278740 357676 278792
rect 357808 278740 357860 278792
rect 386696 278740 386748 278792
rect 397644 278740 397696 278792
rect 397736 278740 397788 278792
rect 408776 278740 408828 278792
rect 451280 278740 451332 278792
rect 451556 278740 451608 278792
rect 270592 278715 270644 278724
rect 270592 278681 270601 278715
rect 270601 278681 270635 278715
rect 270635 278681 270644 278715
rect 270592 278672 270644 278681
rect 397644 278579 397696 278588
rect 397644 278545 397653 278579
rect 397653 278545 397687 278579
rect 397687 278545 397696 278579
rect 397644 278536 397696 278545
rect 254216 277380 254268 277432
rect 259736 277380 259788 277432
rect 356428 277380 356480 277432
rect 356704 277380 356756 277432
rect 545672 274932 545724 274984
rect 550548 274932 550600 274984
rect 369768 274796 369820 274848
rect 370136 274796 370188 274848
rect 295432 273955 295484 273964
rect 295432 273921 295441 273955
rect 295441 273921 295475 273955
rect 295475 273921 295484 273955
rect 295432 273912 295484 273921
rect 451556 273751 451608 273760
rect 451556 273717 451565 273751
rect 451565 273717 451599 273751
rect 451599 273717 451608 273751
rect 451556 273708 451608 273717
rect 232136 273300 232188 273352
rect 232412 273300 232464 273352
rect 330024 273300 330076 273352
rect 356428 273343 356480 273352
rect 356428 273309 356437 273343
rect 356437 273309 356471 273343
rect 356471 273309 356480 273343
rect 356428 273300 356480 273309
rect 357624 273300 357676 273352
rect 367376 273300 367428 273352
rect 236276 273232 236328 273284
rect 386604 273275 386656 273284
rect 386604 273241 386613 273275
rect 386613 273241 386647 273275
rect 386647 273241 386656 273275
rect 386604 273232 386656 273241
rect 408776 273300 408828 273352
rect 244464 273164 244516 273216
rect 272064 273164 272116 273216
rect 283104 273164 283156 273216
rect 294144 273164 294196 273216
rect 330024 273164 330076 273216
rect 334348 273207 334400 273216
rect 334348 273173 334357 273207
rect 334357 273173 334391 273207
rect 334391 273173 334400 273207
rect 334348 273164 334400 273173
rect 357624 273164 357676 273216
rect 367376 273164 367428 273216
rect 376944 273164 376996 273216
rect 400404 273164 400456 273216
rect 400588 273164 400640 273216
rect 408684 273164 408736 273216
rect 244464 273028 244516 273080
rect 249984 273028 250036 273080
rect 272064 273028 272116 273080
rect 283104 273028 283156 273080
rect 294144 273028 294196 273080
rect 376944 273028 376996 273080
rect 249984 272892 250036 272944
rect 321744 272187 321796 272196
rect 321744 272153 321753 272187
rect 321753 272153 321787 272187
rect 321787 272153 321796 272187
rect 321744 272144 321796 272153
rect 327264 272187 327316 272196
rect 327264 272153 327273 272187
rect 327273 272153 327307 272187
rect 327307 272153 327316 272187
rect 327264 272144 327316 272153
rect 232136 271847 232188 271856
rect 232136 271813 232145 271847
rect 232145 271813 232179 271847
rect 232179 271813 232188 271847
rect 232136 271804 232188 271813
rect 241796 270555 241848 270564
rect 241796 270521 241805 270555
rect 241805 270521 241839 270555
rect 241839 270521 241848 270555
rect 241796 270512 241848 270521
rect 288624 270555 288676 270564
rect 288624 270521 288633 270555
rect 288633 270521 288667 270555
rect 288667 270521 288676 270555
rect 288624 270512 288676 270521
rect 305184 270555 305236 270564
rect 305184 270521 305193 270555
rect 305193 270521 305227 270555
rect 305227 270521 305236 270555
rect 305184 270512 305236 270521
rect 309324 270512 309376 270564
rect 309600 270512 309652 270564
rect 310704 270555 310756 270564
rect 310704 270521 310713 270555
rect 310713 270521 310747 270555
rect 310747 270521 310756 270555
rect 310704 270512 310756 270521
rect 346584 270555 346636 270564
rect 346584 270521 346593 270555
rect 346593 270521 346627 270555
rect 346627 270521 346636 270555
rect 346584 270512 346636 270521
rect 381084 270555 381136 270564
rect 381084 270521 381093 270555
rect 381093 270521 381127 270555
rect 381127 270521 381136 270555
rect 381084 270512 381136 270521
rect 382464 270555 382516 270564
rect 382464 270521 382473 270555
rect 382473 270521 382507 270555
rect 382507 270521 382516 270555
rect 382464 270512 382516 270521
rect 416964 270512 417016 270564
rect 433708 270512 433760 270564
rect 466644 270512 466696 270564
rect 472164 270512 472216 270564
rect 243084 270487 243136 270496
rect 243084 270453 243093 270487
rect 243093 270453 243127 270487
rect 243127 270453 243136 270487
rect 243084 270444 243136 270453
rect 252744 270487 252796 270496
rect 252744 270453 252753 270487
rect 252753 270453 252787 270487
rect 252787 270453 252796 270487
rect 252744 270444 252796 270453
rect 267096 270487 267148 270496
rect 267096 270453 267105 270487
rect 267105 270453 267139 270487
rect 267139 270453 267148 270487
rect 267096 270444 267148 270453
rect 356428 270487 356480 270496
rect 356428 270453 356437 270487
rect 356437 270453 356471 270487
rect 356471 270453 356480 270487
rect 356428 270444 356480 270453
rect 400588 270444 400640 270496
rect 309324 270419 309376 270428
rect 309324 270385 309333 270419
rect 309333 270385 309367 270419
rect 309367 270385 309376 270419
rect 309324 270376 309376 270385
rect 381084 270419 381136 270428
rect 381084 270385 381093 270419
rect 381093 270385 381127 270419
rect 381127 270385 381136 270419
rect 381084 270376 381136 270385
rect 386604 269195 386656 269204
rect 386604 269161 386613 269195
rect 386613 269161 386647 269195
rect 386647 269161 386656 269195
rect 386604 269152 386656 269161
rect 287244 269084 287296 269136
rect 287428 269084 287480 269136
rect 393228 269084 393280 269136
rect 393412 269084 393464 269136
rect 397920 269084 397972 269136
rect 480168 269084 480220 269136
rect 480352 269084 480404 269136
rect 281816 269059 281868 269068
rect 281816 269025 281825 269059
rect 281825 269025 281859 269059
rect 281859 269025 281868 269059
rect 281816 269016 281868 269025
rect 292672 269059 292724 269068
rect 292672 269025 292681 269059
rect 292681 269025 292715 269059
rect 292715 269025 292724 269059
rect 292672 269016 292724 269025
rect 375196 269016 375248 269068
rect 375656 269016 375708 269068
rect 347872 267724 347924 267776
rect 348240 267724 348292 267776
rect 386604 264256 386656 264308
rect 392216 264256 392268 264308
rect 233332 263576 233384 263628
rect 233516 263576 233568 263628
rect 236000 263508 236052 263560
rect 356428 263644 356480 263696
rect 324412 263619 324464 263628
rect 324412 263585 324421 263619
rect 324421 263585 324455 263619
rect 324455 263585 324464 263619
rect 324412 263576 324464 263585
rect 334348 263576 334400 263628
rect 342536 263619 342588 263628
rect 342536 263585 342545 263619
rect 342545 263585 342579 263619
rect 342579 263585 342588 263619
rect 342536 263576 342588 263585
rect 353484 263576 353536 263628
rect 331312 263508 331364 263560
rect 295616 263440 295668 263492
rect 331496 263440 331548 263492
rect 334440 263440 334492 263492
rect 408684 263576 408736 263628
rect 422300 263576 422352 263628
rect 422484 263576 422536 263628
rect 427820 263576 427872 263628
rect 428004 263576 428056 263628
rect 356520 263508 356572 263560
rect 353576 263440 353628 263492
rect 408776 263440 408828 263492
rect 451556 263483 451608 263492
rect 451556 263449 451565 263483
rect 451565 263449 451599 263483
rect 451599 263449 451608 263483
rect 451556 263440 451608 263449
rect 232320 262216 232372 262268
rect 243176 260856 243228 260908
rect 252744 260899 252796 260908
rect 252744 260865 252753 260899
rect 252753 260865 252787 260899
rect 252787 260865 252796 260899
rect 252744 260856 252796 260865
rect 267096 260899 267148 260908
rect 267096 260865 267105 260899
rect 267105 260865 267139 260899
rect 267139 260865 267148 260899
rect 267096 260856 267148 260865
rect 270776 260856 270828 260908
rect 309416 260856 309468 260908
rect 324412 260899 324464 260908
rect 324412 260865 324421 260899
rect 324421 260865 324455 260899
rect 324455 260865 324464 260899
rect 324412 260856 324464 260865
rect 342536 260899 342588 260908
rect 342536 260865 342545 260899
rect 342545 260865 342579 260899
rect 342579 260865 342588 260899
rect 342536 260856 342588 260865
rect 359096 260856 359148 260908
rect 359188 260856 359240 260908
rect 381176 260856 381228 260908
rect 397644 260856 397696 260908
rect 397920 260856 397972 260908
rect 400496 260899 400548 260908
rect 400496 260865 400505 260899
rect 400505 260865 400539 260899
rect 400539 260865 400548 260899
rect 400496 260856 400548 260865
rect 241796 260831 241848 260840
rect 241796 260797 241805 260831
rect 241805 260797 241839 260831
rect 241839 260797 241848 260831
rect 241796 260788 241848 260797
rect 265256 260831 265308 260840
rect 265256 260797 265265 260831
rect 265265 260797 265299 260831
rect 265299 260797 265308 260831
rect 265256 260788 265308 260797
rect 272064 260831 272116 260840
rect 272064 260797 272073 260831
rect 272073 260797 272107 260831
rect 272107 260797 272116 260831
rect 272064 260788 272116 260797
rect 277584 260788 277636 260840
rect 277676 260788 277728 260840
rect 288624 260831 288676 260840
rect 288624 260797 288633 260831
rect 288633 260797 288667 260831
rect 288667 260797 288676 260831
rect 288624 260788 288676 260797
rect 294144 260831 294196 260840
rect 294144 260797 294153 260831
rect 294153 260797 294187 260831
rect 294187 260797 294196 260831
rect 294144 260788 294196 260797
rect 295616 260788 295668 260840
rect 305184 260831 305236 260840
rect 305184 260797 305193 260831
rect 305193 260797 305227 260831
rect 305227 260797 305236 260831
rect 305184 260788 305236 260797
rect 310704 260831 310756 260840
rect 310704 260797 310713 260831
rect 310713 260797 310747 260831
rect 310747 260797 310756 260831
rect 310704 260788 310756 260797
rect 318984 260788 319036 260840
rect 319076 260788 319128 260840
rect 321744 260831 321796 260840
rect 321744 260797 321753 260831
rect 321753 260797 321787 260831
rect 321787 260797 321796 260831
rect 321744 260788 321796 260797
rect 327264 260831 327316 260840
rect 327264 260797 327273 260831
rect 327273 260797 327307 260831
rect 327307 260797 327316 260831
rect 327264 260788 327316 260797
rect 331128 260788 331180 260840
rect 331496 260788 331548 260840
rect 334440 260788 334492 260840
rect 346584 260831 346636 260840
rect 346584 260797 346593 260831
rect 346593 260797 346627 260831
rect 346627 260797 346636 260831
rect 346584 260788 346636 260797
rect 382464 260831 382516 260840
rect 382464 260797 382473 260831
rect 382473 260797 382507 260831
rect 382507 260797 382516 260831
rect 382464 260788 382516 260797
rect 416872 260831 416924 260840
rect 416872 260797 416881 260831
rect 416881 260797 416915 260831
rect 416915 260797 416924 260831
rect 416872 260788 416924 260797
rect 433616 260831 433668 260840
rect 433616 260797 433625 260831
rect 433625 260797 433659 260831
rect 433659 260797 433668 260831
rect 433616 260788 433668 260797
rect 466552 260831 466604 260840
rect 466552 260797 466561 260831
rect 466561 260797 466595 260831
rect 466595 260797 466604 260831
rect 466552 260788 466604 260797
rect 472072 260831 472124 260840
rect 472072 260797 472081 260831
rect 472081 260797 472115 260831
rect 472115 260797 472124 260831
rect 472072 260788 472124 260797
rect 292764 260720 292816 260772
rect 309416 260720 309468 260772
rect 342536 260720 342588 260772
rect 282000 259428 282052 259480
rect 351828 259428 351880 259480
rect 352012 259428 352064 259480
rect 386512 259471 386564 259480
rect 386512 259437 386521 259471
rect 386521 259437 386555 259471
rect 386555 259437 386564 259471
rect 386512 259428 386564 259437
rect 392032 259471 392084 259480
rect 392032 259437 392041 259471
rect 392041 259437 392075 259471
rect 392075 259437 392084 259471
rect 392032 259428 392084 259437
rect 393228 259428 393280 259480
rect 393412 259428 393464 259480
rect 451556 259403 451608 259412
rect 451556 259369 451565 259403
rect 451565 259369 451599 259403
rect 451599 259369 451608 259403
rect 451556 259360 451608 259369
rect 356428 258000 356480 258052
rect 356612 258000 356664 258052
rect 408776 258000 408828 258052
rect 408960 258000 409012 258052
rect 254216 253988 254268 254040
rect 259736 253988 259788 254040
rect 261024 253988 261076 254040
rect 330024 253988 330076 254040
rect 370136 253988 370188 254040
rect 375656 253988 375708 254040
rect 232136 253920 232188 253972
rect 232320 253920 232372 253972
rect 397736 253920 397788 253972
rect 236276 253895 236328 253904
rect 236276 253861 236285 253895
rect 236285 253861 236319 253895
rect 236319 253861 236328 253895
rect 236276 253852 236328 253861
rect 244464 253852 244516 253904
rect 261024 253852 261076 253904
rect 283104 253852 283156 253904
rect 330024 253852 330076 253904
rect 376944 253852 376996 253904
rect 387984 253852 388036 253904
rect 400404 253852 400456 253904
rect 400588 253852 400640 253904
rect 244464 253716 244516 253768
rect 249984 253716 250036 253768
rect 267096 253716 267148 253768
rect 283104 253716 283156 253768
rect 376944 253716 376996 253768
rect 387984 253716 388036 253768
rect 267188 253648 267240 253700
rect 249984 253580 250036 253632
rect 334348 251311 334400 251320
rect 334348 251277 334357 251311
rect 334357 251277 334391 251311
rect 334391 251277 334400 251311
rect 334348 251268 334400 251277
rect 381268 251268 381320 251320
rect 241796 251243 241848 251252
rect 241796 251209 241805 251243
rect 241805 251209 241839 251243
rect 241839 251209 241848 251243
rect 241796 251200 241848 251209
rect 265256 251243 265308 251252
rect 265256 251209 265265 251243
rect 265265 251209 265299 251243
rect 265299 251209 265308 251243
rect 265256 251200 265308 251209
rect 270684 251200 270736 251252
rect 270960 251200 271012 251252
rect 272064 251243 272116 251252
rect 272064 251209 272073 251243
rect 272073 251209 272107 251243
rect 272107 251209 272116 251243
rect 272064 251200 272116 251209
rect 288624 251243 288676 251252
rect 288624 251209 288633 251243
rect 288633 251209 288667 251243
rect 288667 251209 288676 251243
rect 288624 251200 288676 251209
rect 294144 251243 294196 251252
rect 294144 251209 294153 251243
rect 294153 251209 294187 251243
rect 294187 251209 294196 251243
rect 294144 251200 294196 251209
rect 295524 251243 295576 251252
rect 295524 251209 295533 251243
rect 295533 251209 295567 251243
rect 295567 251209 295576 251243
rect 295524 251200 295576 251209
rect 305184 251243 305236 251252
rect 305184 251209 305193 251243
rect 305193 251209 305227 251243
rect 305227 251209 305236 251243
rect 305184 251200 305236 251209
rect 309324 251243 309376 251252
rect 309324 251209 309333 251243
rect 309333 251209 309367 251243
rect 309367 251209 309376 251243
rect 309324 251200 309376 251209
rect 310704 251243 310756 251252
rect 310704 251209 310713 251243
rect 310713 251209 310747 251243
rect 310747 251209 310756 251243
rect 310704 251200 310756 251209
rect 321744 251243 321796 251252
rect 321744 251209 321753 251243
rect 321753 251209 321787 251243
rect 321787 251209 321796 251243
rect 321744 251200 321796 251209
rect 327264 251243 327316 251252
rect 327264 251209 327273 251243
rect 327273 251209 327307 251243
rect 327307 251209 327316 251243
rect 327264 251200 327316 251209
rect 342444 251243 342496 251252
rect 342444 251209 342453 251243
rect 342453 251209 342487 251243
rect 342487 251209 342496 251243
rect 342444 251200 342496 251209
rect 346584 251243 346636 251252
rect 346584 251209 346593 251243
rect 346593 251209 346627 251243
rect 346627 251209 346636 251243
rect 346584 251200 346636 251209
rect 352012 251200 352064 251252
rect 352104 251200 352156 251252
rect 381084 251200 381136 251252
rect 382464 251243 382516 251252
rect 382464 251209 382473 251243
rect 382473 251209 382507 251243
rect 382507 251209 382516 251243
rect 382464 251200 382516 251209
rect 292764 251175 292816 251184
rect 292764 251141 292773 251175
rect 292773 251141 292807 251175
rect 292807 251141 292816 251175
rect 292764 251132 292816 251141
rect 298284 251132 298336 251184
rect 298560 251132 298612 251184
rect 334348 251175 334400 251184
rect 334348 251141 334357 251175
rect 334357 251141 334391 251175
rect 334391 251141 334400 251175
rect 334348 251132 334400 251141
rect 353576 251175 353628 251184
rect 353576 251141 353585 251175
rect 353585 251141 353619 251175
rect 353619 251141 353628 251175
rect 353576 251132 353628 251141
rect 386512 251132 386564 251184
rect 386880 251132 386932 251184
rect 393228 251268 393280 251320
rect 416964 251200 417016 251252
rect 433708 251200 433760 251252
rect 466644 251200 466696 251252
rect 472164 251200 472216 251252
rect 400588 251132 400640 251184
rect 407672 251132 407724 251184
rect 407764 251132 407816 251184
rect 393136 251064 393188 251116
rect 348056 250087 348108 250096
rect 348056 250053 348065 250087
rect 348065 250053 348099 250087
rect 348099 250053 348108 250087
rect 348056 250044 348108 250053
rect 359096 249908 359148 249960
rect 287152 249840 287204 249892
rect 287336 249840 287388 249892
rect 359004 249840 359056 249892
rect 364524 249840 364576 249892
rect 364616 249840 364668 249892
rect 397552 249815 397604 249824
rect 397552 249781 397561 249815
rect 397561 249781 397595 249815
rect 397595 249781 397604 249815
rect 397552 249772 397604 249781
rect 480168 249772 480220 249824
rect 480352 249772 480404 249824
rect 254124 248523 254176 248532
rect 254124 248489 254133 248523
rect 254133 248489 254167 248523
rect 254167 248489 254176 248523
rect 254124 248480 254176 248489
rect 259644 248523 259696 248532
rect 259644 248489 259653 248523
rect 259653 248489 259687 248523
rect 259687 248489 259696 248523
rect 259644 248480 259696 248489
rect 370044 248523 370096 248532
rect 370044 248489 370053 248523
rect 370053 248489 370087 248523
rect 370087 248489 370096 248523
rect 370044 248480 370096 248489
rect 375564 248523 375616 248532
rect 375564 248489 375573 248523
rect 375573 248489 375607 248523
rect 375607 248489 375616 248523
rect 375564 248480 375616 248489
rect 254124 248387 254176 248396
rect 254124 248353 254133 248387
rect 254133 248353 254167 248387
rect 254167 248353 254176 248387
rect 254124 248344 254176 248353
rect 259368 248344 259420 248396
rect 259644 248344 259696 248396
rect 282000 248344 282052 248396
rect 282184 248344 282236 248396
rect 356336 248344 356388 248396
rect 356428 248344 356480 248396
rect 370044 248344 370096 248396
rect 370320 248344 370372 248396
rect 375564 248387 375616 248396
rect 375564 248353 375573 248387
rect 375573 248353 375607 248387
rect 375607 248353 375616 248387
rect 375564 248344 375616 248353
rect 397552 244987 397604 244996
rect 397552 244953 397561 244987
rect 397561 244953 397595 244987
rect 397595 244953 397604 244987
rect 397552 244944 397604 244953
rect 233332 244264 233384 244316
rect 233516 244264 233568 244316
rect 231952 244196 232004 244248
rect 232136 244196 232188 244248
rect 265164 244332 265216 244384
rect 243084 244264 243136 244316
rect 254124 244239 254176 244248
rect 254124 244205 254133 244239
rect 254133 244205 254167 244239
rect 254167 244205 254176 244239
rect 254124 244196 254176 244205
rect 270684 244264 270736 244316
rect 324412 244307 324464 244316
rect 324412 244273 324421 244307
rect 324421 244273 324455 244307
rect 324455 244273 324464 244307
rect 324412 244264 324464 244273
rect 364524 244264 364576 244316
rect 381084 244264 381136 244316
rect 422300 244264 422352 244316
rect 422484 244264 422536 244316
rect 427820 244264 427872 244316
rect 428004 244264 428056 244316
rect 243176 244128 243228 244180
rect 265164 244128 265216 244180
rect 270776 244128 270828 244180
rect 334348 244171 334400 244180
rect 334348 244137 334357 244171
rect 334357 244137 334391 244171
rect 334391 244137 334400 244171
rect 334348 244128 334400 244137
rect 364616 244128 364668 244180
rect 381176 244128 381228 244180
rect 451556 244171 451608 244180
rect 451556 244137 451565 244171
rect 451565 244137 451599 244171
rect 451599 244137 451608 244171
rect 451556 244128 451608 244137
rect 375564 242811 375616 242820
rect 375564 242777 375573 242811
rect 375573 242777 375607 242811
rect 375607 242777 375616 242811
rect 375564 242768 375616 242777
rect 324412 241587 324464 241596
rect 324412 241553 324421 241587
rect 324421 241553 324455 241587
rect 324455 241553 324464 241587
rect 324412 241544 324464 241553
rect 266820 241476 266872 241528
rect 266912 241476 266964 241528
rect 295708 241476 295760 241528
rect 295800 241476 295852 241528
rect 309508 241476 309560 241528
rect 309600 241476 309652 241528
rect 331128 241476 331180 241528
rect 331496 241476 331548 241528
rect 348056 241519 348108 241528
rect 348056 241485 348065 241519
rect 348065 241485 348099 241519
rect 348099 241485 348108 241519
rect 348056 241476 348108 241485
rect 353576 241519 353628 241528
rect 353576 241485 353585 241519
rect 353585 241485 353619 241519
rect 353619 241485 353628 241519
rect 353576 241476 353628 241485
rect 392032 241476 392084 241528
rect 392124 241476 392176 241528
rect 400496 241519 400548 241528
rect 400496 241485 400505 241519
rect 400505 241485 400539 241519
rect 400539 241485 400548 241519
rect 400496 241476 400548 241485
rect 324412 241408 324464 241460
rect 324504 241408 324556 241460
rect 466552 241408 466604 241460
rect 466644 241408 466696 241460
rect 287244 240116 287296 240168
rect 287428 240116 287480 240168
rect 292764 240159 292816 240168
rect 292764 240125 292773 240159
rect 292773 240125 292807 240159
rect 292807 240125 292816 240159
rect 292764 240116 292816 240125
rect 359096 240116 359148 240168
rect 359280 240116 359332 240168
rect 392952 240116 393004 240168
rect 393228 240116 393280 240168
rect 397644 240116 397696 240168
rect 407488 240116 407540 240168
rect 407764 240116 407816 240168
rect 292764 240023 292816 240032
rect 292764 239989 292773 240023
rect 292773 239989 292807 240023
rect 292807 239989 292816 240023
rect 292764 239980 292816 239989
rect 356520 238620 356572 238672
rect 356612 238620 356664 238672
rect 2780 237124 2832 237176
rect 4896 237124 4948 237176
rect 236276 234651 236328 234660
rect 236276 234617 236285 234651
rect 236285 234617 236319 234651
rect 236319 234617 236328 234651
rect 236276 234608 236328 234617
rect 255596 234608 255648 234660
rect 261116 234608 261168 234660
rect 281908 234676 281960 234728
rect 397644 234676 397696 234728
rect 321836 234608 321888 234660
rect 330116 234608 330168 234660
rect 357716 234608 357768 234660
rect 367468 234608 367520 234660
rect 381176 234608 381228 234660
rect 451556 234676 451608 234728
rect 255504 234540 255556 234592
rect 261024 234540 261076 234592
rect 281816 234540 281868 234592
rect 309324 234540 309376 234592
rect 309600 234540 309652 234592
rect 321744 234540 321796 234592
rect 330024 234540 330076 234592
rect 357624 234540 357676 234592
rect 367376 234540 367428 234592
rect 376944 234540 376996 234592
rect 381084 234540 381136 234592
rect 387984 234540 388036 234592
rect 397644 234540 397696 234592
rect 400404 234540 400456 234592
rect 400588 234540 400640 234592
rect 451464 234540 451516 234592
rect 351828 234472 351880 234524
rect 352104 234472 352156 234524
rect 376944 234404 376996 234456
rect 387984 234404 388036 234456
rect 359096 233860 359148 233912
rect 359280 233860 359332 233912
rect 369768 233860 369820 233912
rect 370320 233860 370372 233912
rect 265164 231956 265216 232008
rect 334348 231956 334400 232008
rect 265256 231820 265308 231872
rect 271880 231820 271932 231872
rect 272064 231820 272116 231872
rect 277584 231820 277636 231872
rect 277676 231820 277728 231872
rect 293960 231820 294012 231872
rect 294144 231820 294196 231872
rect 295524 231820 295576 231872
rect 295800 231820 295852 231872
rect 298284 231820 298336 231872
rect 298560 231820 298612 231872
rect 305184 231820 305236 231872
rect 305368 231820 305420 231872
rect 310704 231820 310756 231872
rect 310888 231820 310940 231872
rect 318984 231820 319036 231872
rect 319076 231820 319128 231872
rect 331496 231820 331548 231872
rect 334440 231820 334492 231872
rect 346584 231820 346636 231872
rect 346768 231820 346820 231872
rect 364616 231820 364668 231872
rect 382280 231820 382332 231872
rect 382464 231820 382516 231872
rect 386604 231820 386656 231872
rect 386880 231820 386932 231872
rect 416964 231820 417016 231872
rect 417148 231820 417200 231872
rect 433432 231820 433484 231872
rect 433708 231820 433760 231872
rect 472164 231820 472216 231872
rect 472348 231820 472400 231872
rect 259644 231795 259696 231804
rect 259644 231761 259653 231795
rect 259653 231761 259687 231795
rect 259687 231761 259696 231795
rect 259644 231752 259696 231761
rect 309324 231795 309376 231804
rect 309324 231761 309333 231795
rect 309333 231761 309367 231795
rect 309367 231761 309376 231795
rect 309324 231752 309376 231761
rect 364524 231752 364576 231804
rect 347964 230528 348016 230580
rect 348056 230528 348108 230580
rect 353484 230528 353536 230580
rect 353576 230528 353628 230580
rect 242716 230460 242768 230512
rect 242808 230460 242860 230512
rect 270592 230460 270644 230512
rect 270684 230460 270736 230512
rect 292764 230503 292816 230512
rect 292764 230469 292773 230503
rect 292773 230469 292807 230503
rect 292807 230469 292816 230503
rect 292764 230460 292816 230469
rect 480168 230460 480220 230512
rect 480352 230460 480404 230512
rect 281816 229032 281868 229084
rect 332876 229032 332928 229084
rect 333060 229032 333112 229084
rect 331312 227783 331364 227792
rect 331312 227749 331321 227783
rect 331321 227749 331355 227783
rect 331355 227749 331364 227783
rect 331312 227740 331364 227749
rect 236276 225088 236328 225140
rect 233332 224952 233384 225004
rect 233516 224952 233568 225004
rect 236276 224952 236328 225004
rect 270776 224952 270828 225004
rect 347964 224952 348016 225004
rect 353484 224952 353536 225004
rect 381084 224952 381136 225004
rect 422300 224952 422352 225004
rect 422484 224952 422536 225004
rect 427820 224952 427872 225004
rect 428004 224952 428056 225004
rect 451372 224952 451424 225004
rect 270684 224884 270736 224936
rect 236276 224859 236328 224868
rect 236276 224825 236285 224859
rect 236285 224825 236319 224859
rect 236319 224825 236328 224859
rect 236276 224816 236328 224825
rect 348056 224816 348108 224868
rect 353576 224816 353628 224868
rect 408684 224884 408736 224936
rect 408868 224884 408920 224936
rect 381176 224816 381228 224868
rect 242808 222164 242860 222216
rect 243176 222164 243228 222216
rect 252744 222164 252796 222216
rect 252928 222164 252980 222216
rect 259736 222164 259788 222216
rect 295524 222164 295576 222216
rect 295800 222164 295852 222216
rect 298284 222164 298336 222216
rect 298560 222164 298612 222216
rect 309508 222164 309560 222216
rect 392124 222164 392176 222216
rect 392308 222164 392360 222216
rect 400404 222164 400456 222216
rect 400496 222164 400548 222216
rect 451280 222207 451332 222216
rect 451280 222173 451289 222207
rect 451289 222173 451323 222207
rect 451323 222173 451332 222207
rect 451280 222164 451332 222173
rect 466552 222096 466604 222148
rect 466644 222096 466696 222148
rect 243084 222071 243136 222080
rect 243084 222037 243093 222071
rect 243093 222037 243127 222071
rect 243127 222037 243136 222071
rect 243084 222028 243136 222037
rect 292764 220872 292816 220924
rect 266728 220804 266780 220856
rect 266912 220804 266964 220856
rect 292672 220804 292724 220856
rect 327264 220804 327316 220856
rect 327448 220804 327500 220856
rect 351828 220804 351880 220856
rect 352012 220804 352064 220856
rect 358912 220804 358964 220856
rect 359096 220804 359148 220856
rect 364432 220804 364484 220856
rect 364708 220804 364760 220856
rect 369768 220804 369820 220856
rect 369952 220804 370004 220856
rect 375472 220804 375524 220856
rect 375564 220804 375616 220856
rect 287244 220668 287296 220720
rect 287336 220668 287388 220720
rect 375472 220668 375524 220720
rect 375840 220668 375892 220720
rect 334348 219419 334400 219428
rect 334348 219385 334357 219419
rect 334357 219385 334391 219419
rect 334391 219385 334400 219419
rect 334348 219376 334400 219385
rect 358912 217948 358964 218000
rect 359004 217948 359056 218000
rect 259736 217404 259788 217456
rect 259644 217336 259696 217388
rect 231860 216588 231912 216640
rect 232044 216588 232096 216640
rect 321744 215976 321796 216028
rect 321928 215976 321980 216028
rect 324504 215976 324556 216028
rect 324688 215976 324740 216028
rect 270684 215407 270736 215416
rect 270684 215373 270693 215407
rect 270693 215373 270727 215407
rect 270727 215373 270736 215407
rect 270684 215364 270736 215373
rect 236276 215339 236328 215348
rect 236276 215305 236285 215339
rect 236285 215305 236319 215339
rect 236319 215305 236328 215339
rect 236276 215296 236328 215305
rect 255596 215296 255648 215348
rect 261116 215296 261168 215348
rect 330116 215296 330168 215348
rect 357716 215296 357768 215348
rect 367468 215296 367520 215348
rect 408776 215339 408828 215348
rect 408776 215305 408785 215339
rect 408785 215305 408819 215339
rect 408819 215305 408828 215339
rect 408776 215296 408828 215305
rect 255504 215228 255556 215280
rect 261024 215228 261076 215280
rect 283104 215228 283156 215280
rect 330024 215228 330076 215280
rect 357624 215228 357676 215280
rect 367376 215228 367428 215280
rect 376944 215228 376996 215280
rect 387984 215228 388036 215280
rect 283104 215092 283156 215144
rect 376944 215092 376996 215144
rect 387984 215092 388036 215144
rect 364340 212823 364392 212832
rect 364340 212789 364349 212823
rect 364349 212789 364383 212823
rect 364383 212789 364392 212823
rect 364340 212780 364392 212789
rect 265164 212644 265216 212696
rect 254216 212576 254268 212628
rect 356520 212576 356572 212628
rect 243176 212508 243228 212560
rect 252744 212508 252796 212560
rect 252836 212508 252888 212560
rect 254124 212508 254176 212560
rect 265256 212508 265308 212560
rect 271880 212508 271932 212560
rect 272064 212508 272116 212560
rect 277584 212508 277636 212560
rect 277676 212508 277728 212560
rect 288440 212508 288492 212560
rect 288624 212508 288676 212560
rect 298284 212508 298336 212560
rect 298560 212508 298612 212560
rect 305184 212508 305236 212560
rect 305368 212508 305420 212560
rect 308128 212508 308180 212560
rect 308312 212508 308364 212560
rect 310704 212508 310756 212560
rect 310888 212508 310940 212560
rect 318984 212508 319036 212560
rect 319076 212508 319128 212560
rect 346584 212508 346636 212560
rect 346768 212508 346820 212560
rect 347964 212508 348016 212560
rect 348148 212508 348200 212560
rect 352012 212508 352064 212560
rect 352104 212508 352156 212560
rect 353484 212508 353536 212560
rect 353668 212508 353720 212560
rect 356428 212508 356480 212560
rect 364432 212508 364484 212560
rect 382280 212508 382332 212560
rect 382464 212508 382516 212560
rect 386604 212508 386656 212560
rect 386880 212508 386932 212560
rect 400312 212508 400364 212560
rect 400588 212508 400640 212560
rect 408776 212551 408828 212560
rect 408776 212517 408785 212551
rect 408785 212517 408819 212551
rect 408819 212517 408828 212551
rect 408776 212508 408828 212517
rect 416964 212508 417016 212560
rect 417148 212508 417200 212560
rect 433432 212508 433484 212560
rect 433708 212508 433760 212560
rect 472164 212508 472216 212560
rect 472348 212508 472400 212560
rect 259644 212483 259696 212492
rect 259644 212449 259653 212483
rect 259653 212449 259687 212483
rect 259687 212449 259696 212483
rect 259644 212440 259696 212449
rect 270684 212483 270736 212492
rect 270684 212449 270693 212483
rect 270693 212449 270727 212483
rect 270727 212449 270736 212483
rect 270684 212440 270736 212449
rect 281816 212440 281868 212492
rect 334440 212440 334492 212492
rect 369952 212483 370004 212492
rect 369952 212449 369961 212483
rect 369961 212449 369995 212483
rect 369995 212449 370004 212483
rect 369952 212440 370004 212449
rect 364340 212415 364392 212424
rect 364340 212381 364349 212415
rect 364349 212381 364383 212415
rect 364383 212381 364392 212415
rect 364340 212372 364392 212381
rect 292672 211148 292724 211200
rect 292764 211148 292816 211200
rect 255320 211080 255372 211132
rect 255504 211080 255556 211132
rect 270684 211123 270736 211132
rect 270684 211089 270693 211123
rect 270693 211089 270727 211123
rect 270727 211089 270736 211123
rect 270684 211080 270736 211089
rect 351828 211080 351880 211132
rect 352012 211080 352064 211132
rect 295524 209763 295576 209772
rect 295524 209729 295533 209763
rect 295533 209729 295567 209763
rect 295567 209729 295576 209763
rect 295524 209720 295576 209729
rect 331128 209720 331180 209772
rect 331312 209720 331364 209772
rect 332692 209720 332744 209772
rect 332876 209720 332928 209772
rect 386604 209720 386656 209772
rect 386788 209720 386840 209772
rect 364156 208403 364208 208412
rect 364156 208369 364165 208403
rect 364165 208369 364199 208403
rect 364199 208369 364208 208403
rect 364156 208360 364208 208369
rect 236368 207000 236420 207052
rect 236644 206864 236696 206916
rect 233332 205640 233384 205692
rect 233516 205640 233568 205692
rect 243176 205683 243228 205692
rect 243176 205649 243185 205683
rect 243185 205649 243219 205683
rect 243219 205649 243228 205683
rect 243176 205640 243228 205649
rect 265256 205683 265308 205692
rect 265256 205649 265265 205683
rect 265265 205649 265299 205683
rect 265299 205649 265308 205683
rect 265256 205640 265308 205649
rect 292764 205640 292816 205692
rect 298284 205640 298336 205692
rect 336832 205683 336884 205692
rect 336832 205649 336841 205683
rect 336841 205649 336875 205683
rect 336875 205649 336884 205683
rect 336832 205640 336884 205649
rect 347964 205640 348016 205692
rect 422300 205640 422352 205692
rect 422484 205640 422536 205692
rect 427820 205640 427872 205692
rect 428004 205640 428056 205692
rect 270684 205615 270736 205624
rect 270684 205581 270693 205615
rect 270693 205581 270727 205615
rect 270727 205581 270736 205615
rect 270684 205572 270736 205581
rect 298376 205572 298428 205624
rect 348056 205572 348108 205624
rect 292856 205504 292908 205556
rect 336740 204348 336792 204400
rect 338120 204348 338172 204400
rect 375196 204348 375248 204400
rect 384948 204348 385000 204400
rect 425060 204348 425112 204400
rect 434536 204348 434588 204400
rect 521660 204348 521712 204400
rect 526444 204348 526496 204400
rect 309324 202920 309376 202972
rect 309416 202920 309468 202972
rect 480352 202920 480404 202972
rect 243176 202895 243228 202904
rect 243176 202861 243185 202895
rect 243185 202861 243219 202895
rect 243219 202861 243228 202895
rect 243176 202852 243228 202861
rect 259736 202852 259788 202904
rect 265256 202895 265308 202904
rect 265256 202861 265265 202895
rect 265265 202861 265299 202895
rect 265299 202861 265308 202895
rect 265256 202852 265308 202861
rect 281724 202852 281776 202904
rect 281908 202852 281960 202904
rect 327264 202852 327316 202904
rect 327356 202852 327408 202904
rect 336832 202895 336884 202904
rect 336832 202861 336841 202895
rect 336841 202861 336875 202895
rect 336875 202861 336884 202895
rect 336832 202852 336884 202861
rect 364156 202852 364208 202904
rect 364616 202852 364668 202904
rect 369952 202895 370004 202904
rect 369952 202861 369961 202895
rect 369961 202861 369995 202895
rect 369995 202861 370004 202895
rect 369952 202852 370004 202861
rect 295524 202827 295576 202836
rect 295524 202793 295533 202827
rect 295533 202793 295567 202827
rect 295567 202793 295576 202827
rect 295524 202784 295576 202793
rect 318984 202784 319036 202836
rect 319076 202784 319128 202836
rect 400496 202784 400548 202836
rect 400588 202784 400640 202836
rect 243084 202759 243136 202768
rect 243084 202725 243093 202759
rect 243093 202725 243127 202759
rect 243127 202725 243136 202759
rect 243084 202716 243136 202725
rect 480260 201535 480312 201544
rect 480260 201501 480269 201535
rect 480269 201501 480303 201535
rect 480303 201501 480312 201535
rect 480260 201492 480312 201501
rect 255504 201424 255556 201476
rect 255596 201424 255648 201476
rect 281908 201467 281960 201476
rect 281908 201433 281917 201467
rect 281917 201433 281951 201467
rect 281951 201433 281960 201467
rect 281908 201424 281960 201433
rect 287336 201424 287388 201476
rect 309416 201424 309468 201476
rect 321744 201424 321796 201476
rect 321928 201424 321980 201476
rect 324504 201424 324556 201476
rect 324688 201424 324740 201476
rect 352104 201467 352156 201476
rect 352104 201433 352113 201467
rect 352113 201433 352147 201467
rect 352147 201433 352156 201467
rect 352104 201424 352156 201433
rect 369952 201467 370004 201476
rect 369952 201433 369961 201467
rect 369961 201433 369995 201467
rect 369995 201433 370004 201467
rect 369952 201424 370004 201433
rect 287428 201356 287480 201408
rect 255504 200107 255556 200116
rect 255504 200073 255513 200107
rect 255513 200073 255547 200107
rect 255547 200073 255556 200107
rect 255504 200064 255556 200073
rect 294144 200064 294196 200116
rect 294236 200064 294288 200116
rect 295524 200064 295576 200116
rect 386604 200064 386656 200116
rect 386880 200064 386932 200116
rect 332784 198679 332836 198688
rect 332784 198645 332793 198679
rect 332793 198645 332827 198679
rect 332827 198645 332836 198679
rect 332784 198636 332836 198645
rect 386604 198679 386656 198688
rect 386604 198645 386613 198679
rect 386613 198645 386647 198679
rect 386647 198645 386656 198679
rect 386604 198636 386656 198645
rect 236460 198568 236512 198620
rect 236644 198568 236696 198620
rect 259736 198092 259788 198144
rect 259644 198024 259696 198076
rect 359096 197276 359148 197328
rect 342720 196596 342772 196648
rect 342904 196596 342956 196648
rect 365720 196596 365772 196648
rect 365904 196596 365956 196648
rect 270776 196052 270828 196104
rect 364616 196052 364668 196104
rect 364800 196052 364852 196104
rect 375656 196052 375708 196104
rect 433708 196095 433760 196104
rect 433708 196061 433717 196095
rect 433717 196061 433751 196095
rect 433751 196061 433760 196095
rect 433708 196052 433760 196061
rect 367468 195984 367520 196036
rect 480260 195984 480312 196036
rect 277492 195916 277544 195968
rect 277676 195916 277728 195968
rect 367376 195916 367428 195968
rect 376944 195916 376996 195968
rect 387984 195916 388036 195968
rect 480352 195848 480404 195900
rect 376944 195780 376996 195832
rect 387984 195780 388036 195832
rect 265256 193264 265308 193316
rect 356520 193264 356572 193316
rect 243176 193196 243228 193248
rect 252836 193196 252888 193248
rect 253020 193196 253072 193248
rect 265164 193196 265216 193248
rect 267004 193196 267056 193248
rect 267096 193196 267148 193248
rect 288440 193196 288492 193248
rect 288624 193196 288676 193248
rect 292764 193196 292816 193248
rect 292948 193196 293000 193248
rect 298284 193196 298336 193248
rect 298468 193196 298520 193248
rect 305184 193196 305236 193248
rect 305368 193196 305420 193248
rect 308128 193196 308180 193248
rect 308312 193196 308364 193248
rect 327264 193196 327316 193248
rect 327356 193196 327408 193248
rect 330024 193196 330076 193248
rect 334348 193196 334400 193248
rect 334440 193196 334492 193248
rect 336740 193196 336792 193248
rect 336832 193196 336884 193248
rect 346584 193196 346636 193248
rect 346768 193196 346820 193248
rect 347964 193196 348016 193248
rect 348148 193196 348200 193248
rect 353484 193196 353536 193248
rect 353668 193196 353720 193248
rect 356428 193196 356480 193248
rect 375564 193239 375616 193248
rect 375564 193205 375573 193239
rect 375573 193205 375607 193239
rect 375607 193205 375616 193239
rect 375564 193196 375616 193205
rect 382280 193196 382332 193248
rect 382464 193196 382516 193248
rect 392124 193196 392176 193248
rect 392216 193196 392268 193248
rect 397736 193196 397788 193248
rect 397920 193196 397972 193248
rect 408776 193196 408828 193248
rect 408960 193196 409012 193248
rect 416964 193196 417016 193248
rect 417148 193196 417200 193248
rect 433708 193239 433760 193248
rect 433708 193205 433717 193239
rect 433717 193205 433751 193239
rect 433751 193205 433760 193239
rect 433708 193196 433760 193205
rect 472164 193196 472216 193248
rect 472348 193196 472400 193248
rect 270592 193171 270644 193180
rect 270592 193137 270601 193171
rect 270601 193137 270635 193171
rect 270635 193137 270644 193171
rect 270592 193128 270644 193137
rect 281908 193171 281960 193180
rect 281908 193137 281917 193171
rect 281917 193137 281951 193171
rect 281951 193137 281960 193171
rect 281908 193128 281960 193137
rect 330116 193128 330168 193180
rect 352104 193171 352156 193180
rect 352104 193137 352113 193171
rect 352113 193137 352147 193171
rect 352147 193137 352156 193171
rect 352104 193128 352156 193137
rect 369952 193171 370004 193180
rect 369952 193137 369961 193171
rect 369961 193137 369995 193171
rect 369995 193137 370004 193171
rect 369952 193128 370004 193137
rect 231952 191768 232004 191820
rect 232044 191768 232096 191820
rect 270592 191811 270644 191820
rect 270592 191777 270601 191811
rect 270601 191777 270635 191811
rect 270635 191777 270644 191811
rect 270592 191768 270644 191777
rect 255504 190519 255556 190528
rect 255504 190485 255513 190519
rect 255513 190485 255547 190519
rect 255547 190485 255556 190519
rect 255504 190476 255556 190485
rect 364524 190451 364576 190460
rect 364524 190417 364533 190451
rect 364533 190417 364567 190451
rect 364567 190417 364576 190451
rect 364524 190408 364576 190417
rect 332784 189091 332836 189100
rect 332784 189057 332793 189091
rect 332793 189057 332827 189091
rect 332827 189057 332836 189091
rect 332784 189048 332836 189057
rect 236276 187688 236328 187740
rect 236460 187688 236512 187740
rect 359096 187688 359148 187740
rect 236276 187595 236328 187604
rect 236276 187561 236285 187595
rect 236285 187561 236319 187595
rect 236319 187561 236328 187595
rect 236276 187552 236328 187561
rect 451648 186464 451700 186516
rect 272064 186396 272116 186448
rect 277676 186396 277728 186448
rect 298284 186439 298336 186448
rect 298284 186405 298293 186439
rect 298293 186405 298327 186439
rect 298327 186405 298336 186439
rect 298284 186396 298336 186405
rect 321744 186396 321796 186448
rect 324504 186396 324556 186448
rect 233332 186328 233384 186380
rect 233516 186328 233568 186380
rect 243176 186328 243228 186380
rect 243084 186260 243136 186312
rect 327264 186396 327316 186448
rect 357624 186439 357676 186448
rect 357624 186405 357633 186439
rect 357633 186405 357667 186439
rect 357667 186405 357676 186439
rect 357624 186396 357676 186405
rect 422300 186328 422352 186380
rect 422484 186328 422536 186380
rect 427820 186328 427872 186380
rect 428004 186328 428056 186380
rect 451648 186328 451700 186380
rect 327172 186260 327224 186312
rect 364524 186303 364576 186312
rect 364524 186269 364533 186303
rect 364533 186269 364567 186303
rect 364567 186269 364576 186303
rect 364524 186260 364576 186269
rect 386604 186303 386656 186312
rect 386604 186269 386613 186303
rect 386613 186269 386647 186303
rect 386647 186269 386656 186303
rect 386604 186260 386656 186269
rect 277676 186192 277728 186244
rect 382464 183608 382516 183660
rect 252836 183540 252888 183592
rect 253020 183540 253072 183592
rect 271972 183583 272024 183592
rect 271972 183549 271981 183583
rect 271981 183549 272015 183583
rect 272015 183549 272024 183583
rect 271972 183540 272024 183549
rect 287244 183540 287296 183592
rect 287428 183540 287480 183592
rect 298284 183583 298336 183592
rect 298284 183549 298293 183583
rect 298293 183549 298327 183583
rect 298327 183549 298336 183583
rect 298284 183540 298336 183549
rect 309508 183540 309560 183592
rect 321652 183583 321704 183592
rect 321652 183549 321661 183583
rect 321661 183549 321695 183583
rect 321695 183549 321704 183583
rect 321652 183540 321704 183549
rect 324412 183583 324464 183592
rect 324412 183549 324421 183583
rect 324421 183549 324455 183583
rect 324455 183549 324464 183583
rect 324412 183540 324464 183549
rect 329932 183540 329984 183592
rect 330116 183540 330168 183592
rect 331404 183540 331456 183592
rect 331496 183540 331548 183592
rect 334348 183540 334400 183592
rect 334440 183540 334492 183592
rect 336740 183540 336792 183592
rect 336832 183540 336884 183592
rect 347964 183540 348016 183592
rect 348056 183540 348108 183592
rect 352012 183540 352064 183592
rect 352196 183540 352248 183592
rect 353484 183540 353536 183592
rect 353576 183540 353628 183592
rect 356428 183540 356480 183592
rect 356520 183540 356572 183592
rect 270684 183472 270736 183524
rect 295708 183515 295760 183524
rect 295708 183481 295717 183515
rect 295717 183481 295751 183515
rect 295751 183481 295760 183515
rect 295708 183472 295760 183481
rect 382464 183472 382516 183524
rect 416872 183472 416924 183524
rect 416964 183472 417016 183524
rect 332784 182180 332836 182232
rect 231952 182112 232004 182164
rect 232136 182112 232188 182164
rect 265164 182112 265216 182164
rect 265256 182112 265308 182164
rect 267188 182155 267240 182164
rect 267188 182121 267197 182155
rect 267197 182121 267231 182155
rect 267231 182121 267240 182155
rect 267188 182112 267240 182121
rect 287244 182112 287296 182164
rect 287428 182112 287480 182164
rect 292856 182112 292908 182164
rect 292948 182112 293000 182164
rect 298284 182112 298336 182164
rect 298468 182112 298520 182164
rect 331496 182112 331548 182164
rect 331588 182112 331640 182164
rect 332692 182112 332744 182164
rect 334440 182112 334492 182164
rect 334532 182112 334584 182164
rect 336832 182155 336884 182164
rect 336832 182121 336841 182155
rect 336841 182121 336875 182155
rect 336875 182121 336884 182155
rect 336832 182112 336884 182121
rect 365720 182112 365772 182164
rect 365904 182112 365956 182164
rect 372620 181160 372672 181212
rect 382188 181160 382240 181212
rect 364340 181024 364392 181076
rect 553308 180956 553360 181008
rect 554964 180956 555016 181008
rect 475936 180888 475988 180940
rect 476120 180888 476172 180940
rect 364340 180820 364392 180872
rect 425060 180820 425112 180872
rect 434536 180820 434588 180872
rect 521660 180820 521712 180872
rect 526444 180820 526496 180872
rect 255504 180795 255556 180804
rect 255504 180761 255513 180795
rect 255513 180761 255547 180795
rect 255547 180761 255556 180795
rect 255504 180752 255556 180761
rect 348056 180752 348108 180804
rect 352012 180752 352064 180804
rect 353576 180752 353628 180804
rect 357624 179435 357676 179444
rect 357624 179401 357633 179435
rect 357633 179401 357667 179435
rect 357667 179401 357676 179435
rect 357624 179392 357676 179401
rect 359096 179256 359148 179308
rect 359188 179256 359240 179308
rect 252836 178780 252888 178832
rect 480352 178780 480404 178832
rect 480352 178644 480404 178696
rect 236460 178032 236512 178084
rect 364616 176740 364668 176792
rect 386696 176740 386748 176792
rect 329932 176672 329984 176724
rect 244464 176604 244516 176656
rect 346584 176604 346636 176656
rect 364616 176604 364668 176656
rect 386696 176604 386748 176656
rect 397736 176647 397788 176656
rect 397736 176613 397745 176647
rect 397745 176613 397779 176647
rect 397779 176613 397788 176647
rect 397736 176604 397788 176613
rect 330024 176536 330076 176588
rect 336832 176579 336884 176588
rect 336832 176545 336841 176579
rect 336841 176545 336875 176579
rect 336875 176545 336884 176579
rect 336832 176536 336884 176545
rect 244464 176468 244516 176520
rect 249984 176468 250036 176520
rect 346584 176468 346636 176520
rect 249984 176332 250036 176384
rect 309508 174020 309560 174072
rect 241796 173884 241848 173936
rect 241980 173884 242032 173936
rect 243176 173884 243228 173936
rect 243268 173884 243320 173936
rect 252744 173927 252796 173936
rect 252744 173893 252753 173927
rect 252753 173893 252787 173927
rect 252787 173893 252796 173927
rect 252744 173884 252796 173893
rect 254124 173884 254176 173936
rect 254308 173884 254360 173936
rect 259736 173884 259788 173936
rect 259828 173884 259880 173936
rect 266452 173884 266504 173936
rect 266544 173884 266596 173936
rect 270684 173884 270736 173936
rect 270868 173884 270920 173936
rect 271972 173884 272024 173936
rect 272064 173884 272116 173936
rect 288440 173884 288492 173936
rect 288624 173884 288676 173936
rect 294236 173952 294288 174004
rect 308128 173884 308180 173936
rect 308220 173884 308272 173936
rect 310704 173884 310756 173936
rect 310888 173884 310940 173936
rect 321652 173884 321704 173936
rect 321744 173884 321796 173936
rect 324412 173884 324464 173936
rect 324504 173884 324556 173936
rect 327172 173884 327224 173936
rect 327264 173884 327316 173936
rect 370044 173884 370096 173936
rect 370136 173884 370188 173936
rect 397736 173927 397788 173936
rect 397736 173893 397745 173927
rect 397745 173893 397779 173927
rect 397779 173893 397788 173927
rect 397736 173884 397788 173893
rect 408776 173884 408828 173936
rect 408960 173884 409012 173936
rect 422484 173884 422536 173936
rect 422668 173884 422720 173936
rect 433616 173884 433668 173936
rect 433708 173884 433760 173936
rect 472164 173884 472216 173936
rect 472348 173884 472400 173936
rect 294144 173816 294196 173868
rect 309508 173816 309560 173868
rect 267188 173315 267240 173324
rect 267188 173281 267197 173315
rect 267197 173281 267231 173315
rect 267231 173281 267240 173315
rect 267188 173272 267240 173281
rect 295616 172524 295668 172576
rect 295708 172524 295760 172576
rect 254124 172499 254176 172508
rect 254124 172465 254133 172499
rect 254133 172465 254167 172499
rect 254167 172465 254176 172499
rect 254124 172456 254176 172465
rect 259736 172456 259788 172508
rect 272064 172456 272116 172508
rect 292764 172499 292816 172508
rect 292764 172465 292773 172499
rect 292773 172465 292807 172499
rect 292807 172465 292816 172499
rect 292764 172456 292816 172465
rect 332692 172456 332744 172508
rect 332784 172456 332836 172508
rect 342536 172456 342588 172508
rect 451740 172456 451792 172508
rect 452016 172456 452068 172508
rect 288348 170076 288400 170128
rect 296628 170076 296680 170128
rect 328368 170008 328420 170060
rect 336648 170008 336700 170060
rect 365720 169940 365772 169992
rect 368296 169940 368348 169992
rect 454040 169940 454092 169992
rect 458180 169940 458232 169992
rect 514576 169940 514628 169992
rect 516876 169940 516928 169992
rect 475936 169872 475988 169924
rect 476120 169872 476172 169924
rect 309048 169804 309100 169856
rect 317328 169804 317380 169856
rect 425060 169804 425112 169856
rect 434536 169804 434588 169856
rect 524236 169804 524288 169856
rect 526444 169804 526496 169856
rect 299388 169668 299440 169720
rect 302976 169668 303028 169720
rect 376944 169056 376996 169108
rect 377128 169056 377180 169108
rect 480352 169056 480404 169108
rect 480536 169056 480588 169108
rect 321468 168580 321520 168632
rect 321744 168580 321796 168632
rect 382280 167628 382332 167680
rect 243176 167084 243228 167136
rect 233332 167016 233384 167068
rect 233516 167016 233568 167068
rect 270684 167016 270736 167068
rect 318892 167016 318944 167068
rect 319076 167016 319128 167068
rect 254124 166991 254176 167000
rect 254124 166957 254133 166991
rect 254133 166957 254167 166991
rect 254167 166957 254176 166991
rect 254124 166948 254176 166957
rect 255504 166991 255556 167000
rect 255504 166957 255513 166991
rect 255513 166957 255547 166991
rect 255547 166957 255556 166991
rect 255504 166948 255556 166957
rect 356520 167084 356572 167136
rect 400404 167016 400456 167068
rect 400588 167016 400640 167068
rect 422300 167016 422352 167068
rect 422484 167016 422536 167068
rect 466460 167016 466512 167068
rect 466644 167016 466696 167068
rect 270776 166880 270828 166932
rect 356428 166880 356480 166932
rect 2780 165112 2832 165164
rect 4804 165112 4856 165164
rect 231952 164228 232004 164280
rect 232044 164228 232096 164280
rect 298192 164228 298244 164280
rect 298284 164228 298336 164280
rect 393228 164228 393280 164280
rect 265256 164160 265308 164212
rect 266912 164160 266964 164212
rect 267004 164160 267056 164212
rect 292764 164203 292816 164212
rect 292764 164169 292773 164203
rect 292773 164169 292807 164203
rect 292807 164169 292816 164203
rect 292764 164160 292816 164169
rect 308036 164160 308088 164212
rect 308220 164160 308272 164212
rect 310704 164160 310756 164212
rect 310888 164160 310940 164212
rect 327172 164160 327224 164212
rect 329932 164160 329984 164212
rect 330116 164160 330168 164212
rect 370136 164160 370188 164212
rect 376944 164203 376996 164212
rect 376944 164169 376953 164203
rect 376953 164169 376987 164203
rect 376987 164169 376996 164203
rect 376944 164160 376996 164169
rect 386696 164160 386748 164212
rect 386788 164160 386840 164212
rect 397736 164203 397788 164212
rect 397736 164169 397745 164203
rect 397745 164169 397779 164203
rect 397779 164169 397788 164203
rect 397736 164160 397788 164169
rect 400496 164203 400548 164212
rect 400496 164169 400505 164203
rect 400505 164169 400539 164203
rect 400539 164169 400548 164203
rect 400496 164160 400548 164169
rect 408408 164160 408460 164212
rect 408592 164160 408644 164212
rect 416872 164160 416924 164212
rect 416964 164160 417016 164212
rect 422392 164203 422444 164212
rect 422392 164169 422401 164203
rect 422401 164169 422435 164203
rect 422435 164169 422444 164203
rect 422392 164160 422444 164169
rect 466552 164203 466604 164212
rect 466552 164169 466561 164203
rect 466561 164169 466595 164203
rect 466595 164169 466604 164203
rect 466552 164160 466604 164169
rect 472072 164160 472124 164212
rect 472348 164160 472400 164212
rect 480352 164160 480404 164212
rect 327264 164092 327316 164144
rect 393228 164092 393280 164144
rect 242992 162911 243044 162920
rect 242992 162877 243001 162911
rect 243001 162877 243035 162911
rect 243035 162877 243044 162911
rect 242992 162868 243044 162877
rect 259644 162911 259696 162920
rect 259644 162877 259653 162911
rect 259653 162877 259687 162911
rect 259687 162877 259696 162911
rect 259644 162868 259696 162877
rect 271972 162911 272024 162920
rect 271972 162877 271981 162911
rect 271981 162877 272015 162911
rect 272015 162877 272024 162911
rect 271972 162868 272024 162877
rect 342352 162911 342404 162920
rect 342352 162877 342361 162911
rect 342361 162877 342395 162911
rect 342395 162877 342404 162911
rect 342352 162868 342404 162877
rect 347964 162911 348016 162920
rect 347964 162877 347973 162911
rect 347973 162877 348007 162911
rect 348007 162877 348016 162911
rect 347964 162868 348016 162877
rect 352104 162911 352156 162920
rect 352104 162877 352113 162911
rect 352113 162877 352147 162911
rect 352147 162877 352156 162911
rect 352104 162868 352156 162877
rect 353484 162911 353536 162920
rect 353484 162877 353493 162911
rect 353493 162877 353527 162911
rect 353527 162877 353536 162911
rect 353484 162868 353536 162877
rect 298284 162843 298336 162852
rect 298284 162809 298293 162843
rect 298293 162809 298327 162843
rect 298327 162809 298336 162843
rect 298284 162800 298336 162809
rect 308220 162800 308272 162852
rect 308404 162800 308456 162852
rect 327264 162800 327316 162852
rect 327448 162800 327500 162852
rect 393228 162843 393280 162852
rect 393228 162809 393237 162843
rect 393237 162809 393271 162843
rect 393271 162809 393280 162843
rect 393228 162800 393280 162809
rect 451740 162800 451792 162852
rect 334532 161415 334584 161424
rect 334532 161381 334541 161415
rect 334541 161381 334575 161415
rect 334575 161381 334584 161415
rect 334532 161372 334584 161381
rect 356428 161347 356480 161356
rect 356428 161313 356437 161347
rect 356437 161313 356471 161347
rect 356471 161313 356480 161347
rect 356428 161304 356480 161313
rect 321468 159332 321520 159384
rect 321744 159332 321796 159384
rect 252560 157972 252612 158024
rect 252744 157972 252796 158024
rect 271972 158015 272024 158024
rect 271972 157981 271981 158015
rect 271981 157981 272015 158015
rect 272015 157981 272024 158015
rect 271972 157972 272024 157981
rect 405740 157700 405792 157752
rect 415308 157700 415360 157752
rect 387984 157428 388036 157480
rect 521660 157428 521712 157480
rect 526444 157428 526496 157480
rect 232044 157360 232096 157412
rect 232136 157292 232188 157344
rect 298284 157335 298336 157344
rect 298284 157301 298293 157335
rect 298293 157301 298327 157335
rect 298327 157301 298336 157335
rect 298284 157292 298336 157301
rect 324504 157360 324556 157412
rect 346584 157292 346636 157344
rect 387984 157292 388036 157344
rect 400496 157335 400548 157344
rect 400496 157301 400505 157335
rect 400505 157301 400539 157335
rect 400539 157301 400548 157335
rect 400496 157292 400548 157301
rect 422392 157335 422444 157344
rect 422392 157301 422401 157335
rect 422401 157301 422435 157335
rect 422435 157301 422444 157335
rect 422392 157292 422444 157301
rect 466552 157335 466604 157344
rect 466552 157301 466561 157335
rect 466561 157301 466595 157335
rect 466595 157301 466604 157335
rect 466552 157292 466604 157301
rect 324412 157224 324464 157276
rect 346584 157156 346636 157208
rect 292856 155864 292908 155916
rect 265164 154683 265216 154692
rect 265164 154649 265173 154683
rect 265173 154649 265207 154683
rect 265207 154649 265216 154683
rect 265164 154640 265216 154649
rect 266544 154572 266596 154624
rect 266636 154572 266688 154624
rect 370044 154615 370096 154624
rect 370044 154581 370053 154615
rect 370053 154581 370087 154615
rect 370087 154581 370096 154615
rect 370044 154572 370096 154581
rect 376944 154615 376996 154624
rect 376944 154581 376953 154615
rect 376953 154581 376987 154615
rect 376987 154581 376996 154615
rect 376944 154572 376996 154581
rect 382464 154615 382516 154624
rect 382464 154581 382473 154615
rect 382473 154581 382507 154615
rect 382507 154581 382516 154615
rect 382464 154572 382516 154581
rect 397736 154615 397788 154624
rect 397736 154581 397745 154615
rect 397745 154581 397779 154615
rect 397779 154581 397788 154615
rect 397736 154572 397788 154581
rect 242992 154547 243044 154556
rect 242992 154513 243001 154547
rect 243001 154513 243035 154547
rect 243035 154513 243044 154547
rect 242992 154504 243044 154513
rect 331404 154547 331456 154556
rect 331404 154513 331413 154547
rect 331413 154513 331447 154547
rect 331447 154513 331456 154547
rect 331404 154504 331456 154513
rect 375564 154547 375616 154556
rect 375564 154513 375573 154547
rect 375573 154513 375607 154547
rect 375607 154513 375616 154547
rect 375564 154504 375616 154513
rect 381084 154547 381136 154556
rect 381084 154513 381093 154547
rect 381093 154513 381127 154547
rect 381127 154513 381136 154547
rect 381084 154504 381136 154513
rect 386604 154504 386656 154556
rect 386788 154504 386840 154556
rect 392124 154547 392176 154556
rect 392124 154513 392133 154547
rect 392133 154513 392167 154547
rect 392167 154513 392176 154547
rect 392124 154504 392176 154513
rect 254124 153212 254176 153264
rect 254400 153212 254452 153264
rect 480260 153255 480312 153264
rect 480260 153221 480269 153255
rect 480269 153221 480303 153255
rect 480303 153221 480312 153255
rect 480260 153212 480312 153221
rect 240232 153144 240284 153196
rect 240508 153144 240560 153196
rect 281724 153144 281776 153196
rect 281816 153144 281868 153196
rect 334624 153144 334676 153196
rect 254400 153119 254452 153128
rect 254400 153085 254409 153119
rect 254409 153085 254443 153119
rect 254443 153085 254452 153119
rect 254400 153076 254452 153085
rect 356428 151827 356480 151836
rect 356428 151793 356437 151827
rect 356437 151793 356471 151827
rect 356471 151793 356480 151827
rect 356428 151784 356480 151793
rect 236368 151759 236420 151768
rect 236368 151725 236377 151759
rect 236377 151725 236411 151759
rect 236411 151725 236420 151759
rect 236368 151716 236420 151725
rect 334624 151716 334676 151768
rect 271972 148631 272024 148640
rect 271972 148597 271981 148631
rect 271981 148597 272015 148631
rect 272015 148597 272024 148631
rect 271972 148588 272024 148597
rect 265164 147704 265216 147756
rect 433616 147704 433668 147756
rect 233332 147636 233384 147688
rect 233516 147636 233568 147688
rect 309324 147636 309376 147688
rect 318892 147636 318944 147688
rect 319076 147636 319128 147688
rect 364524 147636 364576 147688
rect 370044 147636 370096 147688
rect 400404 147636 400456 147688
rect 400588 147636 400640 147688
rect 422300 147636 422352 147688
rect 422484 147636 422536 147688
rect 243084 147568 243136 147620
rect 265164 147568 265216 147620
rect 292764 147611 292816 147620
rect 292764 147577 292773 147611
rect 292773 147577 292807 147611
rect 292807 147577 292816 147611
rect 292764 147568 292816 147577
rect 309416 147568 309468 147620
rect 364616 147568 364668 147620
rect 466460 147636 466512 147688
rect 466644 147636 466696 147688
rect 370136 147568 370188 147620
rect 375564 147611 375616 147620
rect 375564 147577 375573 147611
rect 375573 147577 375607 147611
rect 375607 147577 375616 147611
rect 375564 147568 375616 147577
rect 381084 147611 381136 147620
rect 381084 147577 381093 147611
rect 381093 147577 381127 147611
rect 381127 147577 381136 147611
rect 381084 147568 381136 147577
rect 392124 147611 392176 147620
rect 392124 147577 392133 147611
rect 392133 147577 392167 147611
rect 392167 147577 392176 147611
rect 392124 147568 392176 147577
rect 433616 147568 433668 147620
rect 451556 147611 451608 147620
rect 451556 147577 451565 147611
rect 451565 147577 451599 147611
rect 451599 147577 451608 147611
rect 451556 147568 451608 147577
rect 331496 147432 331548 147484
rect 393228 145027 393280 145036
rect 393228 144993 393237 145027
rect 393237 144993 393271 145027
rect 393271 144993 393280 145027
rect 393228 144984 393280 144993
rect 252744 144916 252796 144968
rect 252836 144916 252888 144968
rect 283104 144916 283156 144968
rect 308128 144916 308180 144968
rect 308220 144916 308272 144968
rect 397736 144959 397788 144968
rect 397736 144925 397745 144959
rect 397745 144925 397779 144959
rect 397779 144925 397788 144959
rect 397736 144916 397788 144925
rect 243176 144848 243228 144900
rect 243268 144848 243320 144900
rect 271972 144848 272024 144900
rect 272064 144848 272116 144900
rect 283012 144848 283064 144900
rect 292764 144891 292816 144900
rect 292764 144857 292773 144891
rect 292773 144857 292807 144891
rect 292807 144857 292816 144891
rect 292764 144848 292816 144857
rect 294052 144848 294104 144900
rect 294236 144848 294288 144900
rect 295616 144848 295668 144900
rect 295708 144848 295760 144900
rect 298284 144848 298336 144900
rect 298468 144848 298520 144900
rect 347964 144848 348016 144900
rect 348056 144848 348108 144900
rect 352012 144848 352064 144900
rect 352196 144848 352248 144900
rect 353484 144848 353536 144900
rect 353576 144848 353628 144900
rect 357532 144848 357584 144900
rect 357716 144848 357768 144900
rect 359004 144848 359056 144900
rect 359188 144848 359240 144900
rect 364524 144848 364576 144900
rect 364616 144848 364668 144900
rect 370136 144848 370188 144900
rect 370228 144848 370280 144900
rect 375564 144848 375616 144900
rect 375656 144848 375708 144900
rect 400496 144891 400548 144900
rect 400496 144857 400505 144891
rect 400505 144857 400539 144891
rect 400539 144857 400548 144891
rect 400496 144848 400548 144857
rect 422392 144891 422444 144900
rect 422392 144857 422401 144891
rect 422401 144857 422435 144891
rect 422435 144857 422444 144891
rect 422392 144848 422444 144857
rect 427728 144848 427780 144900
rect 428004 144848 428056 144900
rect 466552 144891 466604 144900
rect 466552 144857 466561 144891
rect 466561 144857 466595 144891
rect 466595 144857 466604 144891
rect 466552 144848 466604 144857
rect 381176 144780 381228 144832
rect 254124 143556 254176 143608
rect 397736 143599 397788 143608
rect 397736 143565 397745 143599
rect 397745 143565 397779 143599
rect 397779 143565 397788 143599
rect 397736 143556 397788 143565
rect 252744 143488 252796 143540
rect 252928 143488 252980 143540
rect 254216 143531 254268 143540
rect 254216 143497 254225 143531
rect 254225 143497 254259 143531
rect 254259 143497 254268 143531
rect 254216 143488 254268 143497
rect 259736 143488 259788 143540
rect 266452 143488 266504 143540
rect 266728 143488 266780 143540
rect 287244 143531 287296 143540
rect 287244 143497 287253 143531
rect 287253 143497 287287 143531
rect 287287 143497 287296 143531
rect 287244 143488 287296 143497
rect 305092 143531 305144 143540
rect 305092 143497 305101 143531
rect 305101 143497 305135 143531
rect 305135 143497 305144 143531
rect 305092 143488 305144 143497
rect 309416 143488 309468 143540
rect 309692 143488 309744 143540
rect 321652 143531 321704 143540
rect 321652 143497 321661 143531
rect 321661 143497 321695 143531
rect 321695 143497 321704 143531
rect 321652 143488 321704 143497
rect 393228 143531 393280 143540
rect 393228 143497 393237 143531
rect 393237 143497 393271 143531
rect 393271 143497 393280 143531
rect 393228 143488 393280 143497
rect 480260 143488 480312 143540
rect 480444 143488 480496 143540
rect 236368 143463 236420 143472
rect 236368 143429 236377 143463
rect 236377 143429 236411 143463
rect 236411 143429 236420 143463
rect 236368 143420 236420 143429
rect 334440 142171 334492 142180
rect 334440 142137 334449 142171
rect 334449 142137 334483 142171
rect 334483 142137 334492 142171
rect 334440 142128 334492 142137
rect 283012 142103 283064 142112
rect 283012 142069 283021 142103
rect 283021 142069 283055 142103
rect 283055 142069 283064 142103
rect 283012 142060 283064 142069
rect 408868 140020 408920 140072
rect 409052 140020 409104 140072
rect 277676 138048 277728 138100
rect 376944 137980 376996 138032
rect 382464 137980 382516 138032
rect 416872 137980 416924 138032
rect 451556 137980 451608 138032
rect 472072 137980 472124 138032
rect 277584 137912 277636 137964
rect 400496 137955 400548 137964
rect 400496 137921 400505 137955
rect 400505 137921 400539 137955
rect 400539 137921 400548 137955
rect 400496 137912 400548 137921
rect 416780 137912 416832 137964
rect 422392 137955 422444 137964
rect 422392 137921 422401 137955
rect 422401 137921 422435 137955
rect 422435 137921 422444 137955
rect 422392 137912 422444 137921
rect 451740 137912 451792 137964
rect 466552 137955 466604 137964
rect 466552 137921 466561 137955
rect 466561 137921 466595 137955
rect 466595 137921 466604 137955
rect 466552 137912 466604 137921
rect 471980 137912 472032 137964
rect 376944 137844 376996 137896
rect 382464 137844 382516 137896
rect 292764 135303 292816 135312
rect 292764 135269 292773 135303
rect 292773 135269 292807 135303
rect 292807 135269 292816 135303
rect 292764 135260 292816 135269
rect 365996 135260 366048 135312
rect 381084 135303 381136 135312
rect 381084 135269 381093 135303
rect 381093 135269 381127 135303
rect 381127 135269 381136 135303
rect 381084 135260 381136 135269
rect 243084 135192 243136 135244
rect 243268 135192 243320 135244
rect 271880 135192 271932 135244
rect 271972 135192 272024 135244
rect 321652 135235 321704 135244
rect 321652 135201 321661 135235
rect 321661 135201 321695 135235
rect 321695 135201 321704 135235
rect 321652 135192 321704 135201
rect 365904 135192 365956 135244
rect 367376 135192 367428 135244
rect 367560 135192 367612 135244
rect 298008 134104 298060 134156
rect 301596 134104 301648 134156
rect 383660 134036 383712 134088
rect 385224 134036 385276 134088
rect 287244 133943 287296 133952
rect 287244 133909 287253 133943
rect 287253 133909 287287 133943
rect 287287 133909 287296 133943
rect 287244 133900 287296 133909
rect 305092 133943 305144 133952
rect 305092 133909 305101 133943
rect 305101 133909 305135 133943
rect 305135 133909 305144 133943
rect 305092 133900 305144 133909
rect 393228 133943 393280 133952
rect 393228 133909 393237 133943
rect 393237 133909 393271 133943
rect 393271 133909 393280 133943
rect 393228 133900 393280 133909
rect 521660 133900 521712 133952
rect 526444 133900 526496 133952
rect 243268 133875 243320 133884
rect 243268 133841 243277 133875
rect 243277 133841 243311 133875
rect 243311 133841 243320 133875
rect 243268 133832 243320 133841
rect 292764 133875 292816 133884
rect 292764 133841 292773 133875
rect 292773 133841 292807 133875
rect 292807 133841 292816 133875
rect 292764 133832 292816 133841
rect 334440 133875 334492 133884
rect 334440 133841 334449 133875
rect 334449 133841 334483 133875
rect 334483 133841 334492 133875
rect 334440 133832 334492 133841
rect 353484 133875 353536 133884
rect 353484 133841 353493 133875
rect 353493 133841 353527 133875
rect 353527 133841 353536 133875
rect 353484 133832 353536 133841
rect 356428 133875 356480 133884
rect 356428 133841 356437 133875
rect 356437 133841 356471 133875
rect 356471 133841 356480 133875
rect 356428 133832 356480 133841
rect 386604 133875 386656 133884
rect 386604 133841 386613 133875
rect 386613 133841 386647 133875
rect 386647 133841 386656 133875
rect 386604 133832 386656 133841
rect 259736 133764 259788 133816
rect 283104 132472 283156 132524
rect 267280 132404 267332 132456
rect 233332 128324 233384 128376
rect 233516 128324 233568 128376
rect 318892 128324 318944 128376
rect 319076 128324 319128 128376
rect 330024 128392 330076 128444
rect 422300 128324 422352 128376
rect 422484 128324 422536 128376
rect 451556 128324 451608 128376
rect 451740 128324 451792 128376
rect 329932 128256 329984 128308
rect 236276 125740 236328 125792
rect 305092 125672 305144 125724
rect 236276 125604 236328 125656
rect 240140 125604 240192 125656
rect 240324 125604 240376 125656
rect 347964 125604 348016 125656
rect 364524 125604 364576 125656
rect 365904 125604 365956 125656
rect 365996 125604 366048 125656
rect 400496 125604 400548 125656
rect 400588 125604 400640 125656
rect 270592 125536 270644 125588
rect 270776 125536 270828 125588
rect 271972 125536 272024 125588
rect 272064 125536 272116 125588
rect 292764 125579 292816 125588
rect 292764 125545 292773 125579
rect 292773 125545 292807 125579
rect 292807 125545 292816 125579
rect 292764 125536 292816 125545
rect 310704 125579 310756 125588
rect 310704 125545 310713 125579
rect 310713 125545 310747 125579
rect 310747 125545 310756 125579
rect 310704 125536 310756 125545
rect 342444 125536 342496 125588
rect 342628 125536 342680 125588
rect 348056 125468 348108 125520
rect 369952 125536 370004 125588
rect 370136 125536 370188 125588
rect 371424 125536 371476 125588
rect 371516 125536 371568 125588
rect 381176 125579 381228 125588
rect 381176 125545 381185 125579
rect 381185 125545 381219 125579
rect 381219 125545 381228 125579
rect 381176 125536 381228 125545
rect 433616 125579 433668 125588
rect 433616 125545 433625 125579
rect 433625 125545 433659 125579
rect 433659 125545 433668 125579
rect 433616 125536 433668 125545
rect 364616 125468 364668 125520
rect 259736 124312 259788 124364
rect 243360 124176 243412 124228
rect 254216 124219 254268 124228
rect 254216 124185 254225 124219
rect 254225 124185 254259 124219
rect 254259 124185 254268 124219
rect 254216 124176 254268 124185
rect 259736 124176 259788 124228
rect 304908 124219 304960 124228
rect 304908 124185 304917 124219
rect 304917 124185 304951 124219
rect 304951 124185 304960 124219
rect 304908 124176 304960 124185
rect 334440 124219 334492 124228
rect 334440 124185 334449 124219
rect 334449 124185 334483 124219
rect 334483 124185 334492 124219
rect 334440 124176 334492 124185
rect 353576 124176 353628 124228
rect 356428 124219 356480 124228
rect 356428 124185 356437 124219
rect 356437 124185 356471 124219
rect 356471 124185 356480 124219
rect 356428 124176 356480 124185
rect 397736 124176 397788 124228
rect 397920 124176 397972 124228
rect 240140 124151 240192 124160
rect 240140 124117 240149 124151
rect 240149 124117 240183 124151
rect 240183 124117 240192 124151
rect 249984 124151 250036 124160
rect 240140 124108 240192 124117
rect 249984 124117 249993 124151
rect 249993 124117 250027 124151
rect 250027 124117 250036 124151
rect 249984 124108 250036 124117
rect 271972 124151 272024 124160
rect 271972 124117 271981 124151
rect 271981 124117 272015 124151
rect 272015 124117 272024 124151
rect 271972 124108 272024 124117
rect 287244 124108 287296 124160
rect 292856 124151 292908 124160
rect 292856 124117 292865 124151
rect 292865 124117 292899 124151
rect 292899 124117 292908 124151
rect 292856 124108 292908 124117
rect 295524 124108 295576 124160
rect 295616 124108 295668 124160
rect 309508 124108 309560 124160
rect 309324 123972 309376 124024
rect 327172 124108 327224 124160
rect 327264 124108 327316 124160
rect 342628 124151 342680 124160
rect 342628 124117 342637 124151
rect 342637 124117 342671 124151
rect 342671 124117 342680 124151
rect 342628 124108 342680 124117
rect 365904 124151 365956 124160
rect 365904 124117 365913 124151
rect 365913 124117 365947 124151
rect 365947 124117 365956 124151
rect 365904 124108 365956 124117
rect 407764 124151 407816 124160
rect 407764 124117 407773 124151
rect 407773 124117 407807 124151
rect 407807 124117 407816 124151
rect 407764 124108 407816 124117
rect 466644 124151 466696 124160
rect 466644 124117 466653 124151
rect 466653 124117 466687 124151
rect 466687 124117 466696 124151
rect 466644 124108 466696 124117
rect 345940 123224 345992 123276
rect 354588 123224 354640 123276
rect 454040 123020 454092 123072
rect 458180 123020 458232 123072
rect 514576 123020 514628 123072
rect 516876 123020 516928 123072
rect 475936 122952 475988 123004
rect 478144 122952 478196 123004
rect 386696 122884 386748 122936
rect 425060 122884 425112 122936
rect 434536 122884 434588 122936
rect 524236 122884 524288 122936
rect 526444 122884 526496 122936
rect 266636 122816 266688 122868
rect 266728 122816 266780 122868
rect 267188 122859 267240 122868
rect 267188 122825 267197 122859
rect 267197 122825 267231 122859
rect 267231 122825 267240 122859
rect 267188 122816 267240 122825
rect 259736 122748 259788 122800
rect 259828 122748 259880 122800
rect 327264 122791 327316 122800
rect 327264 122757 327273 122791
rect 327273 122757 327307 122791
rect 327307 122757 327316 122791
rect 327264 122748 327316 122757
rect 2964 122204 3016 122256
rect 6184 122204 6236 122256
rect 386604 121388 386656 121440
rect 265072 120708 265124 120760
rect 265256 120708 265308 120760
rect 329932 120232 329984 120284
rect 252560 119348 252612 119400
rect 321744 118847 321796 118856
rect 321744 118813 321753 118847
rect 321753 118813 321787 118847
rect 321787 118813 321796 118847
rect 321744 118804 321796 118813
rect 324504 118847 324556 118856
rect 324504 118813 324513 118847
rect 324513 118813 324547 118847
rect 324547 118813 324556 118847
rect 324504 118804 324556 118813
rect 298284 118736 298336 118788
rect 357624 118736 357676 118788
rect 451740 118736 451792 118788
rect 231860 118668 231912 118720
rect 232044 118668 232096 118720
rect 244372 118668 244424 118720
rect 308128 118668 308180 118720
rect 332784 118668 332836 118720
rect 336832 118668 336884 118720
rect 346584 118668 346636 118720
rect 244464 118600 244516 118652
rect 310704 118643 310756 118652
rect 310704 118609 310713 118643
rect 310713 118609 310747 118643
rect 310747 118609 310756 118643
rect 310704 118600 310756 118609
rect 416872 118668 416924 118720
rect 422392 118668 422444 118720
rect 357624 118600 357676 118652
rect 365904 118643 365956 118652
rect 365904 118609 365913 118643
rect 365913 118609 365947 118643
rect 365947 118609 365956 118643
rect 365904 118600 365956 118609
rect 416780 118600 416832 118652
rect 472072 118668 472124 118720
rect 422484 118600 422536 118652
rect 451740 118600 451792 118652
rect 471980 118600 472032 118652
rect 308128 118532 308180 118584
rect 332784 118532 332836 118584
rect 336832 118532 336884 118584
rect 346584 118532 346636 118584
rect 236276 117988 236328 118040
rect 236460 117988 236512 118040
rect 266912 117784 266964 117836
rect 267188 117784 267240 117836
rect 381176 115991 381228 116000
rect 381176 115957 381185 115991
rect 381185 115957 381219 115991
rect 381219 115957 381228 115991
rect 381176 115948 381228 115957
rect 400404 115948 400456 116000
rect 400496 115948 400548 116000
rect 433616 115991 433668 116000
rect 433616 115957 433625 115991
rect 433625 115957 433659 115991
rect 433659 115957 433668 115991
rect 433616 115948 433668 115957
rect 254124 115880 254176 115932
rect 254216 115880 254268 115932
rect 277492 115880 277544 115932
rect 277676 115880 277728 115932
rect 305092 115923 305144 115932
rect 305092 115889 305101 115923
rect 305101 115889 305135 115923
rect 305135 115889 305144 115923
rect 305092 115880 305144 115889
rect 271972 115379 272024 115388
rect 271972 115345 271981 115379
rect 271981 115345 272015 115379
rect 272015 115345 272024 115379
rect 271972 115336 272024 115345
rect 393228 114656 393280 114708
rect 294052 114588 294104 114640
rect 240232 114520 240284 114572
rect 243176 114520 243228 114572
rect 243360 114520 243412 114572
rect 249984 114563 250036 114572
rect 249984 114529 249993 114563
rect 249993 114529 250027 114563
rect 250027 114529 250036 114563
rect 249984 114520 250036 114529
rect 283104 114520 283156 114572
rect 283196 114520 283248 114572
rect 287152 114563 287204 114572
rect 287152 114529 287161 114563
rect 287161 114529 287195 114563
rect 287195 114529 287204 114563
rect 287152 114520 287204 114529
rect 353576 114588 353628 114640
rect 356428 114588 356480 114640
rect 369952 114588 370004 114640
rect 294144 114520 294196 114572
rect 321744 114563 321796 114572
rect 321744 114529 321753 114563
rect 321753 114529 321787 114563
rect 321787 114529 321796 114563
rect 321744 114520 321796 114529
rect 324504 114563 324556 114572
rect 324504 114529 324513 114563
rect 324513 114529 324547 114563
rect 324547 114529 324556 114563
rect 324504 114520 324556 114529
rect 342628 114563 342680 114572
rect 342628 114529 342637 114563
rect 342637 114529 342671 114563
rect 342671 114529 342680 114563
rect 342628 114520 342680 114529
rect 348056 114563 348108 114572
rect 348056 114529 348065 114563
rect 348065 114529 348099 114563
rect 348099 114529 348108 114563
rect 348056 114520 348108 114529
rect 353484 114520 353536 114572
rect 408592 114588 408644 114640
rect 408776 114588 408828 114640
rect 356520 114520 356572 114572
rect 370044 114520 370096 114572
rect 393228 114520 393280 114572
rect 407764 114563 407816 114572
rect 407764 114529 407773 114563
rect 407773 114529 407807 114563
rect 407807 114529 407816 114563
rect 407764 114520 407816 114529
rect 466828 114520 466880 114572
rect 254124 114452 254176 114504
rect 254216 114452 254268 114504
rect 397736 114452 397788 114504
rect 408776 114452 408828 114504
rect 292948 113160 293000 113212
rect 327264 113203 327316 113212
rect 327264 113169 327273 113203
rect 327273 113169 327307 113203
rect 327307 113169 327316 113203
rect 327264 113160 327316 113169
rect 348056 113203 348108 113212
rect 348056 113169 348065 113203
rect 348065 113169 348099 113203
rect 348099 113169 348108 113203
rect 348056 113160 348108 113169
rect 236368 113092 236420 113144
rect 295524 113135 295576 113144
rect 295524 113101 295533 113135
rect 295533 113101 295567 113135
rect 295567 113101 295576 113135
rect 295524 113092 295576 113101
rect 336740 110712 336792 110764
rect 346216 110712 346268 110764
rect 425060 110508 425112 110560
rect 434536 110508 434588 110560
rect 521660 110508 521712 110560
rect 526444 110508 526496 110560
rect 243084 109735 243136 109744
rect 243084 109701 243093 109735
rect 243093 109701 243127 109735
rect 243127 109701 243136 109735
rect 243084 109692 243136 109701
rect 282920 109692 282972 109744
rect 283104 109692 283156 109744
rect 294144 109692 294196 109744
rect 294144 109556 294196 109608
rect 364524 109080 364576 109132
rect 364708 109080 364760 109132
rect 233332 109012 233384 109064
rect 233516 109012 233568 109064
rect 422300 109012 422352 109064
rect 422484 109012 422536 109064
rect 252744 106335 252796 106344
rect 252744 106301 252753 106335
rect 252753 106301 252787 106335
rect 252787 106301 252796 106335
rect 252744 106292 252796 106301
rect 305184 106292 305236 106344
rect 319076 106292 319128 106344
rect 330024 106335 330076 106344
rect 330024 106301 330033 106335
rect 330033 106301 330067 106335
rect 330067 106301 330076 106335
rect 330024 106292 330076 106301
rect 342536 106292 342588 106344
rect 342628 106292 342680 106344
rect 370044 106292 370096 106344
rect 240232 106224 240284 106276
rect 241796 106224 241848 106276
rect 241980 106224 242032 106276
rect 281632 106267 281684 106276
rect 281632 106233 281641 106267
rect 281641 106233 281675 106267
rect 281675 106233 281684 106267
rect 281632 106224 281684 106233
rect 309232 106224 309284 106276
rect 309324 106224 309376 106276
rect 324504 106267 324556 106276
rect 324504 106233 324513 106267
rect 324513 106233 324547 106267
rect 324547 106233 324556 106267
rect 324504 106224 324556 106233
rect 357624 106267 357676 106276
rect 357624 106233 357633 106267
rect 357633 106233 357667 106267
rect 357667 106233 357676 106267
rect 357624 106224 357676 106233
rect 243268 106156 243320 106208
rect 319076 106156 319128 106208
rect 392032 106224 392084 106276
rect 392308 106224 392360 106276
rect 422392 106267 422444 106276
rect 422392 106233 422401 106267
rect 422401 106233 422435 106267
rect 422435 106233 422444 106267
rect 422392 106224 422444 106233
rect 427912 106267 427964 106276
rect 427912 106233 427921 106267
rect 427921 106233 427955 106267
rect 427955 106233 427964 106267
rect 427912 106224 427964 106233
rect 433616 106267 433668 106276
rect 433616 106233 433625 106267
rect 433625 106233 433659 106267
rect 433659 106233 433668 106267
rect 433616 106224 433668 106233
rect 370136 106156 370188 106208
rect 327264 104932 327316 104984
rect 397644 104975 397696 104984
rect 397644 104941 397653 104975
rect 397653 104941 397687 104975
rect 397687 104941 397696 104975
rect 397644 104932 397696 104941
rect 271880 104864 271932 104916
rect 271972 104864 272024 104916
rect 292764 104864 292816 104916
rect 292948 104864 293000 104916
rect 327172 104864 327224 104916
rect 347872 104864 347924 104916
rect 348056 104864 348108 104916
rect 408684 104907 408736 104916
rect 408684 104873 408693 104907
rect 408693 104873 408727 104907
rect 408727 104873 408736 104907
rect 408684 104864 408736 104873
rect 282920 104839 282972 104848
rect 282920 104805 282929 104839
rect 282929 104805 282963 104839
rect 282963 104805 282972 104839
rect 282920 104796 282972 104805
rect 309232 104839 309284 104848
rect 309232 104805 309241 104839
rect 309241 104805 309275 104839
rect 309275 104805 309284 104839
rect 309232 104796 309284 104805
rect 319076 104839 319128 104848
rect 319076 104805 319085 104839
rect 319085 104805 319119 104839
rect 319119 104805 319128 104839
rect 319076 104796 319128 104805
rect 393228 104796 393280 104848
rect 397644 104796 397696 104848
rect 400496 104839 400548 104848
rect 400496 104805 400505 104839
rect 400505 104805 400539 104839
rect 400539 104805 400548 104839
rect 400496 104796 400548 104805
rect 407764 104839 407816 104848
rect 407764 104805 407773 104839
rect 407773 104805 407807 104839
rect 407807 104805 407816 104839
rect 407764 104796 407816 104805
rect 480444 104839 480496 104848
rect 480444 104805 480453 104839
rect 480453 104805 480487 104839
rect 480487 104805 480496 104839
rect 480444 104796 480496 104805
rect 397828 104728 397880 104780
rect 364524 103708 364576 103760
rect 364708 103708 364760 103760
rect 236276 103547 236328 103556
rect 236276 103513 236285 103547
rect 236285 103513 236319 103547
rect 236319 103513 236328 103547
rect 236276 103504 236328 103513
rect 295524 103547 295576 103556
rect 295524 103513 295533 103547
rect 295533 103513 295567 103547
rect 295567 103513 295576 103547
rect 295524 103504 295576 103513
rect 386880 103547 386932 103556
rect 386880 103513 386889 103547
rect 386889 103513 386923 103547
rect 386923 103513 386932 103547
rect 386880 103504 386932 103513
rect 254216 103479 254268 103488
rect 254216 103445 254225 103479
rect 254225 103445 254259 103479
rect 254259 103445 254268 103479
rect 254216 103436 254268 103445
rect 353576 103436 353628 103488
rect 356612 103436 356664 103488
rect 370136 103436 370188 103488
rect 370320 103436 370372 103488
rect 356428 103368 356480 103420
rect 236276 103096 236328 103148
rect 236460 103096 236512 103148
rect 298376 102187 298428 102196
rect 298376 102153 298385 102187
rect 298385 102153 298419 102187
rect 298419 102153 298428 102187
rect 298376 102144 298428 102153
rect 266544 102076 266596 102128
rect 231860 101396 231912 101448
rect 232044 101396 232096 101448
rect 281632 101371 281684 101380
rect 281632 101337 281641 101371
rect 281641 101337 281675 101371
rect 281675 101337 281684 101371
rect 281632 101328 281684 101337
rect 408776 100079 408828 100088
rect 408776 100045 408785 100079
rect 408785 100045 408819 100079
rect 408819 100045 408828 100079
rect 408776 100036 408828 100045
rect 244464 99424 244516 99476
rect 277584 99424 277636 99476
rect 298376 99467 298428 99476
rect 298376 99433 298385 99467
rect 298385 99433 298419 99467
rect 298419 99433 298428 99467
rect 298376 99424 298428 99433
rect 288624 99399 288676 99408
rect 288624 99365 288633 99399
rect 288633 99365 288667 99399
rect 288667 99365 288676 99399
rect 288624 99356 288676 99365
rect 308128 99399 308180 99408
rect 308128 99365 308137 99399
rect 308137 99365 308171 99399
rect 308171 99365 308180 99399
rect 308128 99356 308180 99365
rect 310704 99399 310756 99408
rect 310704 99365 310713 99399
rect 310713 99365 310747 99399
rect 310747 99365 310756 99399
rect 310704 99356 310756 99365
rect 416872 99356 416924 99408
rect 472072 99356 472124 99408
rect 244464 99288 244516 99340
rect 271880 99288 271932 99340
rect 272064 99288 272116 99340
rect 277584 99288 277636 99340
rect 416780 99288 416832 99340
rect 422392 99331 422444 99340
rect 422392 99297 422401 99331
rect 422401 99297 422435 99331
rect 422435 99297 422444 99331
rect 422392 99288 422444 99297
rect 427912 99331 427964 99340
rect 427912 99297 427921 99331
rect 427921 99297 427955 99331
rect 427955 99297 427964 99331
rect 427912 99288 427964 99297
rect 433616 99331 433668 99340
rect 433616 99297 433625 99331
rect 433625 99297 433659 99331
rect 433659 99297 433668 99331
rect 433616 99288 433668 99297
rect 471980 99288 472032 99340
rect 393136 98719 393188 98728
rect 393136 98685 393145 98719
rect 393145 98685 393179 98719
rect 393179 98685 393188 98719
rect 393136 98676 393188 98685
rect 240140 96679 240192 96688
rect 240140 96645 240149 96679
rect 240149 96645 240183 96679
rect 240183 96645 240192 96679
rect 240140 96636 240192 96645
rect 288624 96679 288676 96688
rect 288624 96645 288633 96679
rect 288633 96645 288667 96679
rect 288667 96645 288676 96679
rect 288624 96636 288676 96645
rect 308128 96679 308180 96688
rect 308128 96645 308137 96679
rect 308137 96645 308171 96679
rect 308171 96645 308180 96679
rect 308128 96636 308180 96645
rect 310704 96679 310756 96688
rect 310704 96645 310713 96679
rect 310713 96645 310747 96679
rect 310747 96645 310756 96679
rect 310704 96636 310756 96645
rect 324504 96679 324556 96688
rect 324504 96645 324513 96679
rect 324513 96645 324547 96679
rect 324547 96645 324556 96679
rect 324504 96636 324556 96645
rect 357716 96500 357768 96552
rect 259644 95208 259696 95260
rect 259828 95208 259880 95260
rect 266912 95208 266964 95260
rect 267096 95208 267148 95260
rect 282920 95251 282972 95260
rect 282920 95217 282929 95251
rect 282929 95217 282963 95251
rect 282963 95217 282972 95251
rect 282920 95208 282972 95217
rect 295524 95208 295576 95260
rect 319076 95251 319128 95260
rect 319076 95217 319085 95251
rect 319085 95217 319119 95251
rect 319119 95217 319128 95251
rect 319076 95208 319128 95217
rect 327172 95208 327224 95260
rect 327264 95208 327316 95260
rect 400588 95208 400640 95260
rect 466552 95208 466604 95260
rect 466828 95208 466880 95260
rect 480536 95208 480588 95260
rect 236368 95140 236420 95192
rect 240140 95183 240192 95192
rect 240140 95149 240149 95183
rect 240149 95149 240183 95183
rect 240183 95149 240192 95183
rect 240140 95140 240192 95149
rect 287244 95140 287296 95192
rect 295616 95072 295668 95124
rect 351828 95072 351880 95124
rect 352196 95072 352248 95124
rect 386788 93916 386840 93968
rect 254216 93891 254268 93900
rect 254216 93857 254225 93891
rect 254225 93857 254259 93891
rect 254259 93857 254268 93891
rect 254216 93848 254268 93857
rect 353484 93891 353536 93900
rect 353484 93857 353493 93891
rect 353493 93857 353527 93891
rect 353527 93857 353536 93891
rect 353484 93848 353536 93857
rect 386880 93848 386932 93900
rect 294144 93780 294196 93832
rect 298376 93823 298428 93832
rect 298376 93789 298385 93823
rect 298385 93789 298419 93823
rect 298419 93789 298428 93823
rect 298376 93780 298428 93789
rect 364708 93780 364760 93832
rect 375564 93551 375616 93560
rect 375564 93517 375573 93551
rect 375573 93517 375607 93551
rect 375607 93517 375616 93551
rect 375564 93508 375616 93517
rect 266452 92531 266504 92540
rect 266452 92497 266461 92531
rect 266461 92497 266495 92531
rect 266495 92497 266504 92531
rect 266452 92488 266504 92497
rect 242992 91740 243044 91792
rect 243452 91740 243504 91792
rect 342444 89768 342496 89820
rect 381084 89768 381136 89820
rect 233332 89700 233384 89752
rect 233516 89700 233568 89752
rect 259644 89700 259696 89752
rect 356428 89700 356480 89752
rect 422300 89700 422352 89752
rect 422484 89700 422536 89752
rect 427820 89700 427872 89752
rect 428004 89700 428056 89752
rect 309324 89632 309376 89684
rect 342444 89632 342496 89684
rect 259736 89564 259788 89616
rect 359004 89632 359056 89684
rect 359188 89632 359240 89684
rect 408776 89675 408828 89684
rect 408776 89641 408785 89675
rect 408785 89641 408819 89675
rect 408819 89641 408828 89675
rect 408776 89632 408828 89641
rect 356520 89564 356572 89616
rect 298376 88952 298428 89004
rect 365628 87184 365680 87236
rect 373908 87184 373960 87236
rect 267740 87116 267792 87168
rect 273720 87116 273772 87168
rect 328552 87116 328604 87168
rect 338028 87116 338080 87168
rect 340788 87116 340840 87168
rect 354588 87116 354640 87168
rect 415400 87048 415452 87100
rect 424784 87048 424836 87100
rect 475936 87048 475988 87100
rect 476120 87048 476172 87100
rect 572628 87048 572680 87100
rect 576768 87048 576820 87100
rect 267096 86980 267148 87032
rect 331312 86980 331364 87032
rect 331404 86980 331456 87032
rect 334256 86980 334308 87032
rect 334440 86980 334492 87032
rect 380992 87023 381044 87032
rect 380992 86989 381001 87023
rect 381001 86989 381035 87023
rect 381035 86989 381044 87023
rect 380992 86980 381044 86989
rect 407856 86980 407908 87032
rect 425060 86980 425112 87032
rect 434536 86980 434588 87032
rect 466552 86980 466604 87032
rect 466644 86980 466696 87032
rect 241796 86955 241848 86964
rect 241796 86921 241805 86955
rect 241805 86921 241839 86955
rect 241839 86921 241848 86955
rect 241796 86912 241848 86921
rect 267004 86912 267056 86964
rect 288624 86955 288676 86964
rect 288624 86921 288633 86955
rect 288633 86921 288667 86955
rect 288667 86921 288676 86955
rect 288624 86912 288676 86921
rect 305184 86955 305236 86964
rect 305184 86921 305193 86955
rect 305193 86921 305227 86955
rect 305227 86921 305236 86955
rect 305184 86912 305236 86921
rect 308128 86955 308180 86964
rect 308128 86921 308137 86955
rect 308137 86921 308171 86955
rect 308171 86921 308180 86955
rect 308128 86912 308180 86921
rect 310704 86955 310756 86964
rect 310704 86921 310713 86955
rect 310713 86921 310747 86955
rect 310747 86921 310756 86955
rect 310704 86912 310756 86921
rect 324504 86912 324556 86964
rect 324596 86912 324648 86964
rect 342536 86955 342588 86964
rect 342536 86921 342545 86955
rect 342545 86921 342579 86955
rect 342579 86921 342588 86955
rect 342536 86912 342588 86921
rect 346584 86955 346636 86964
rect 346584 86921 346593 86955
rect 346593 86921 346627 86955
rect 346627 86921 346636 86955
rect 346584 86912 346636 86921
rect 382464 86955 382516 86964
rect 382464 86921 382473 86955
rect 382473 86921 382507 86955
rect 382507 86921 382516 86955
rect 382464 86912 382516 86921
rect 422392 86955 422444 86964
rect 422392 86921 422401 86955
rect 422401 86921 422435 86955
rect 422435 86921 422444 86955
rect 422392 86912 422444 86921
rect 270592 86844 270644 86896
rect 270868 86844 270920 86896
rect 357532 86844 357584 86896
rect 357716 86844 357768 86896
rect 240232 85620 240284 85672
rect 287152 85663 287204 85672
rect 287152 85629 287161 85663
rect 287161 85629 287195 85663
rect 287195 85629 287204 85663
rect 287152 85620 287204 85629
rect 236276 85595 236328 85604
rect 236276 85561 236285 85595
rect 236285 85561 236319 85595
rect 236319 85561 236328 85595
rect 236276 85552 236328 85561
rect 295524 85552 295576 85604
rect 295616 85552 295668 85604
rect 327172 85552 327224 85604
rect 327264 85552 327316 85604
rect 347872 85552 347924 85604
rect 348056 85552 348108 85604
rect 352104 85552 352156 85604
rect 352196 85552 352248 85604
rect 375656 85552 375708 85604
rect 249984 85527 250036 85536
rect 249984 85493 249993 85527
rect 249993 85493 250027 85527
rect 250027 85493 250036 85527
rect 249984 85484 250036 85493
rect 254216 85484 254268 85536
rect 287152 85484 287204 85536
rect 334256 85527 334308 85536
rect 334256 85493 334265 85527
rect 334265 85493 334299 85527
rect 334299 85493 334308 85527
rect 334256 85484 334308 85493
rect 380992 85527 381044 85536
rect 380992 85493 381001 85527
rect 381001 85493 381035 85527
rect 381035 85493 381044 85527
rect 380992 85484 381044 85493
rect 407764 85527 407816 85536
rect 407764 85493 407773 85527
rect 407773 85493 407807 85527
rect 407807 85493 407816 85527
rect 407764 85484 407816 85493
rect 408868 85484 408920 85536
rect 466460 85527 466512 85536
rect 466460 85493 466469 85527
rect 466469 85493 466503 85527
rect 466503 85493 466512 85527
rect 466460 85484 466512 85493
rect 472072 85527 472124 85536
rect 472072 85493 472081 85527
rect 472081 85493 472115 85527
rect 472115 85493 472124 85527
rect 472072 85484 472124 85493
rect 480444 85527 480496 85536
rect 480444 85493 480453 85527
rect 480453 85493 480487 85527
rect 480487 85493 480496 85527
rect 480444 85484 480496 85493
rect 236276 85459 236328 85468
rect 236276 85425 236285 85459
rect 236285 85425 236319 85459
rect 236319 85425 236328 85459
rect 236276 85416 236328 85425
rect 272064 84260 272116 84312
rect 271972 84192 272024 84244
rect 294144 84235 294196 84244
rect 294144 84201 294153 84235
rect 294153 84201 294187 84235
rect 294187 84201 294196 84235
rect 294144 84192 294196 84201
rect 298560 84235 298612 84244
rect 298560 84201 298569 84235
rect 298569 84201 298603 84235
rect 298603 84201 298612 84235
rect 364524 84235 364576 84244
rect 298560 84192 298612 84201
rect 364524 84201 364533 84235
rect 364533 84201 364567 84235
rect 364567 84201 364576 84235
rect 364524 84192 364576 84201
rect 259736 84124 259788 84176
rect 353484 84124 353536 84176
rect 356520 84124 356572 84176
rect 357716 84167 357768 84176
rect 357716 84133 357725 84167
rect 357725 84133 357759 84167
rect 357759 84133 357768 84167
rect 357716 84124 357768 84133
rect 359004 84167 359056 84176
rect 359004 84133 359013 84167
rect 359013 84133 359047 84167
rect 359047 84133 359056 84167
rect 359004 84124 359056 84133
rect 353392 84056 353444 84108
rect 356520 83988 356572 84040
rect 271972 82807 272024 82816
rect 271972 82773 271981 82807
rect 271981 82773 272015 82807
rect 272015 82773 272024 82807
rect 271972 82764 272024 82773
rect 356520 82764 356572 82816
rect 243360 80724 243412 80776
rect 433708 80180 433760 80232
rect 309324 80087 309376 80096
rect 309324 80053 309333 80087
rect 309333 80053 309367 80087
rect 309367 80053 309376 80087
rect 309324 80044 309376 80053
rect 332784 80044 332836 80096
rect 336832 80044 336884 80096
rect 365904 80044 365956 80096
rect 376944 80044 376996 80096
rect 387984 80044 388036 80096
rect 255504 80019 255556 80028
rect 255504 79985 255513 80019
rect 255513 79985 255547 80019
rect 255547 79985 255556 80019
rect 255504 79976 255556 79985
rect 342536 80019 342588 80028
rect 342536 79985 342545 80019
rect 342545 79985 342579 80019
rect 342579 79985 342588 80019
rect 342536 79976 342588 79985
rect 346584 80019 346636 80028
rect 346584 79985 346593 80019
rect 346593 79985 346627 80019
rect 346627 79985 346636 80019
rect 346584 79976 346636 79985
rect 332784 79908 332836 79960
rect 336832 79908 336884 79960
rect 365904 79908 365956 79960
rect 376944 79908 376996 79960
rect 387984 79908 388036 79960
rect 249984 79339 250036 79348
rect 249984 79305 249993 79339
rect 249993 79305 250027 79339
rect 250027 79305 250036 79339
rect 249984 79296 250036 79305
rect 334440 79296 334492 79348
rect 3332 79160 3384 79212
rect 7656 79160 7708 79212
rect 266636 77936 266688 77988
rect 359280 77936 359332 77988
rect 386604 77392 386656 77444
rect 348056 77324 348108 77376
rect 352104 77324 352156 77376
rect 392216 77324 392268 77376
rect 416872 77324 416924 77376
rect 416964 77324 417016 77376
rect 232044 77256 232096 77308
rect 241796 77299 241848 77308
rect 241796 77265 241805 77299
rect 241805 77265 241839 77299
rect 241839 77265 241848 77299
rect 241796 77256 241848 77265
rect 270684 77256 270736 77308
rect 270868 77256 270920 77308
rect 281724 77299 281776 77308
rect 281724 77265 281733 77299
rect 281733 77265 281767 77299
rect 281767 77265 281776 77299
rect 281724 77256 281776 77265
rect 288624 77299 288676 77308
rect 288624 77265 288633 77299
rect 288633 77265 288667 77299
rect 288667 77265 288676 77299
rect 288624 77256 288676 77265
rect 305184 77299 305236 77308
rect 305184 77265 305193 77299
rect 305193 77265 305227 77299
rect 305227 77265 305236 77299
rect 305184 77256 305236 77265
rect 308128 77299 308180 77308
rect 308128 77265 308137 77299
rect 308137 77265 308171 77299
rect 308171 77265 308180 77299
rect 308128 77256 308180 77265
rect 309232 77256 309284 77308
rect 310704 77299 310756 77308
rect 310704 77265 310713 77299
rect 310713 77265 310747 77299
rect 310747 77265 310756 77299
rect 310704 77256 310756 77265
rect 347964 77256 348016 77308
rect 386604 77256 386656 77308
rect 392124 77256 392176 77308
rect 422484 77256 422536 77308
rect 433616 77299 433668 77308
rect 433616 77265 433625 77299
rect 433625 77265 433659 77299
rect 433659 77265 433668 77299
rect 433616 77256 433668 77265
rect 232044 77120 232096 77172
rect 466552 77120 466604 77172
rect 480536 77120 480588 77172
rect 427912 76347 427964 76356
rect 427912 76313 427921 76347
rect 427921 76313 427955 76347
rect 427955 76313 427964 76347
rect 427912 76304 427964 76313
rect 398748 76236 398800 76288
rect 405648 76236 405700 76288
rect 309048 76168 309100 76220
rect 317328 76168 317380 76220
rect 514576 76100 514628 76152
rect 516876 76100 516928 76152
rect 475936 76032 475988 76084
rect 478144 76032 478196 76084
rect 283472 75964 283524 76016
rect 290556 75964 290608 76016
rect 346216 75964 346268 76016
rect 370044 75964 370096 76016
rect 370320 75964 370372 76016
rect 408684 76007 408736 76016
rect 408684 75973 408693 76007
rect 408693 75973 408727 76007
rect 408727 75973 408736 76007
rect 408684 75964 408736 75973
rect 524236 75964 524288 76016
rect 526444 75964 526496 76016
rect 236368 75896 236420 75948
rect 240232 75896 240284 75948
rect 240416 75896 240468 75948
rect 281724 75939 281776 75948
rect 281724 75905 281733 75939
rect 281733 75905 281767 75939
rect 281767 75905 281776 75939
rect 281724 75896 281776 75905
rect 287244 75939 287296 75948
rect 287244 75905 287253 75939
rect 287253 75905 287287 75939
rect 287287 75905 287296 75939
rect 287244 75896 287296 75905
rect 319076 75896 319128 75948
rect 319168 75896 319220 75948
rect 327172 75896 327224 75948
rect 327264 75896 327316 75948
rect 346308 75896 346360 75948
rect 381084 75896 381136 75948
rect 382464 75939 382516 75948
rect 382464 75905 382473 75939
rect 382473 75905 382507 75939
rect 382507 75905 382516 75939
rect 382464 75896 382516 75905
rect 407764 75939 407816 75948
rect 407764 75905 407773 75939
rect 407773 75905 407807 75939
rect 407807 75905 407816 75939
rect 407764 75896 407816 75905
rect 270684 75871 270736 75880
rect 270684 75837 270693 75871
rect 270693 75837 270727 75871
rect 270727 75837 270736 75871
rect 270684 75828 270736 75837
rect 375564 75871 375616 75880
rect 375564 75837 375573 75871
rect 375573 75837 375607 75871
rect 375607 75837 375616 75871
rect 375564 75828 375616 75837
rect 408684 75871 408736 75880
rect 408684 75837 408693 75871
rect 408693 75837 408727 75871
rect 408727 75837 408736 75871
rect 408684 75828 408736 75837
rect 267004 74604 267056 74656
rect 255504 74579 255556 74588
rect 255504 74545 255513 74579
rect 255513 74545 255547 74579
rect 255547 74545 255556 74579
rect 255504 74536 255556 74545
rect 266820 74468 266872 74520
rect 357716 74579 357768 74588
rect 357716 74545 357725 74579
rect 357725 74545 357759 74579
rect 357759 74545 357768 74579
rect 357716 74536 357768 74545
rect 334440 74468 334492 74520
rect 364524 74511 364576 74520
rect 364524 74477 364533 74511
rect 364533 74477 364567 74511
rect 364567 74477 364576 74511
rect 364524 74468 364576 74477
rect 271972 73219 272024 73228
rect 271972 73185 271981 73219
rect 271981 73185 272015 73219
rect 272015 73185 272024 73219
rect 271972 73176 272024 73185
rect 356428 73219 356480 73228
rect 356428 73185 356437 73219
rect 356437 73185 356471 73219
rect 356471 73185 356480 73219
rect 356428 73176 356480 73185
rect 359188 73108 359240 73160
rect 359280 73108 359332 73160
rect 294052 72428 294104 72480
rect 294236 72428 294288 72480
rect 259644 71111 259696 71120
rect 259644 71077 259653 71111
rect 259653 71077 259687 71111
rect 259687 71077 259696 71111
rect 259644 71068 259696 71077
rect 244464 70499 244516 70508
rect 244464 70465 244473 70499
rect 244473 70465 244507 70499
rect 244507 70465 244516 70499
rect 244464 70456 244516 70465
rect 277584 70456 277636 70508
rect 305184 70499 305236 70508
rect 305184 70465 305193 70499
rect 305193 70465 305227 70499
rect 305227 70465 305236 70499
rect 305184 70456 305236 70465
rect 416964 70456 417016 70508
rect 277584 70320 277636 70372
rect 416872 70320 416924 70372
rect 236368 67804 236420 67856
rect 331404 67736 331456 67788
rect 309232 67668 309284 67720
rect 240140 67600 240192 67652
rect 240324 67600 240376 67652
rect 243176 67643 243228 67652
rect 243176 67609 243185 67643
rect 243185 67609 243219 67643
rect 243219 67609 243228 67643
rect 243176 67600 243228 67609
rect 244464 67643 244516 67652
rect 244464 67609 244473 67643
rect 244473 67609 244507 67643
rect 244507 67609 244516 67643
rect 244464 67600 244516 67609
rect 254124 67643 254176 67652
rect 254124 67609 254133 67643
rect 254133 67609 254167 67643
rect 254167 67609 254176 67643
rect 254124 67600 254176 67609
rect 292764 67600 292816 67652
rect 292856 67600 292908 67652
rect 305184 67643 305236 67652
rect 305184 67609 305193 67643
rect 305193 67609 305227 67643
rect 305227 67609 305236 67643
rect 305184 67600 305236 67609
rect 376944 67668 376996 67720
rect 309324 67600 309376 67652
rect 310612 67600 310664 67652
rect 310704 67600 310756 67652
rect 318984 67600 319036 67652
rect 319076 67600 319128 67652
rect 331404 67600 331456 67652
rect 376852 67600 376904 67652
rect 400496 67600 400548 67652
rect 400588 67600 400640 67652
rect 422392 67600 422444 67652
rect 422484 67600 422536 67652
rect 428004 67600 428056 67652
rect 472072 67643 472124 67652
rect 472072 67609 472081 67643
rect 472081 67609 472115 67643
rect 472115 67609 472124 67643
rect 472072 67600 472124 67609
rect 231860 67532 231912 67584
rect 232044 67532 232096 67584
rect 236276 67532 236328 67584
rect 281724 67575 281776 67584
rect 281724 67541 281733 67575
rect 281733 67541 281767 67575
rect 281767 67541 281776 67575
rect 281724 67532 281776 67541
rect 381084 67575 381136 67584
rect 381084 67541 381093 67575
rect 381093 67541 381127 67575
rect 381127 67541 381136 67575
rect 381084 67532 381136 67541
rect 416872 67532 416924 67584
rect 417056 67532 417108 67584
rect 480260 67532 480312 67584
rect 480444 67532 480496 67584
rect 370044 66376 370096 66428
rect 265164 66240 265216 66292
rect 265256 66240 265308 66292
rect 270776 66240 270828 66292
rect 249892 66172 249944 66224
rect 249984 66172 250036 66224
rect 283196 66308 283248 66360
rect 287244 66308 287296 66360
rect 352012 66283 352064 66292
rect 352012 66249 352021 66283
rect 352021 66249 352055 66283
rect 352055 66249 352064 66283
rect 352012 66240 352064 66249
rect 370044 66240 370096 66292
rect 292764 66215 292816 66224
rect 292764 66181 292773 66215
rect 292773 66181 292807 66215
rect 292807 66181 292816 66215
rect 292764 66172 292816 66181
rect 293960 66172 294012 66224
rect 294236 66172 294288 66224
rect 324504 66215 324556 66224
rect 324504 66181 324513 66215
rect 324513 66181 324547 66215
rect 324547 66181 324556 66215
rect 324504 66172 324556 66181
rect 346584 66172 346636 66224
rect 346676 66172 346728 66224
rect 408776 66240 408828 66292
rect 393228 66172 393280 66224
rect 407764 66215 407816 66224
rect 407764 66181 407773 66215
rect 407773 66181 407807 66215
rect 407807 66181 407816 66215
rect 407764 66172 407816 66181
rect 393136 66104 393188 66156
rect 334348 64991 334400 65000
rect 334348 64957 334357 64991
rect 334357 64957 334391 64991
rect 334391 64957 334400 64991
rect 334348 64948 334400 64957
rect 266452 64923 266504 64932
rect 266452 64889 266461 64923
rect 266461 64889 266495 64923
rect 266495 64889 266504 64923
rect 266452 64880 266504 64889
rect 357624 64880 357676 64932
rect 357716 64880 357768 64932
rect 364524 64923 364576 64932
rect 364524 64889 364533 64923
rect 364533 64889 364567 64923
rect 364567 64889 364576 64923
rect 364524 64880 364576 64889
rect 249892 64855 249944 64864
rect 249892 64821 249901 64855
rect 249901 64821 249935 64855
rect 249935 64821 249944 64855
rect 249892 64812 249944 64821
rect 255504 64855 255556 64864
rect 255504 64821 255513 64855
rect 255513 64821 255547 64855
rect 255547 64821 255556 64855
rect 255504 64812 255556 64821
rect 271972 64812 272024 64864
rect 272064 64812 272116 64864
rect 310612 64855 310664 64864
rect 310612 64821 310621 64855
rect 310621 64821 310655 64855
rect 310655 64821 310664 64855
rect 310612 64812 310664 64821
rect 331404 64855 331456 64864
rect 331404 64821 331413 64855
rect 331413 64821 331447 64855
rect 331447 64821 331456 64855
rect 331404 64812 331456 64821
rect 334348 64855 334400 64864
rect 334348 64821 334357 64855
rect 334357 64821 334391 64855
rect 334391 64821 334400 64855
rect 334348 64812 334400 64821
rect 356428 64812 356480 64864
rect 356612 64812 356664 64864
rect 240048 64472 240100 64524
rect 248328 64472 248380 64524
rect 267648 63860 267700 63912
rect 275928 63860 275980 63912
rect 355508 63792 355560 63844
rect 360384 63792 360436 63844
rect 393320 63792 393372 63844
rect 405648 63792 405700 63844
rect 346216 63588 346268 63640
rect 346492 63588 346544 63640
rect 521660 63588 521712 63640
rect 526444 63588 526496 63640
rect 337476 63520 337528 63572
rect 344928 63520 344980 63572
rect 356612 63452 356664 63504
rect 359188 63495 359240 63504
rect 359188 63461 359197 63495
rect 359197 63461 359231 63495
rect 359231 63461 359240 63495
rect 359188 63452 359240 63461
rect 281724 61455 281776 61464
rect 281724 61421 281733 61455
rect 281733 61421 281767 61455
rect 281767 61421 281776 61455
rect 281724 61412 281776 61421
rect 386604 61412 386656 61464
rect 386788 61412 386840 61464
rect 259644 60800 259696 60852
rect 270776 60800 270828 60852
rect 347964 60800 348016 60852
rect 259644 60664 259696 60716
rect 270684 60664 270736 60716
rect 347964 60664 348016 60716
rect 433524 60664 433576 60716
rect 433708 60664 433760 60716
rect 471980 60664 472032 60716
rect 472164 60664 472216 60716
rect 240140 57944 240192 57996
rect 240232 57944 240284 57996
rect 244372 57944 244424 57996
rect 244556 57944 244608 57996
rect 298284 57944 298336 57996
rect 308036 57944 308088 57996
rect 308128 57944 308180 57996
rect 381084 57987 381136 57996
rect 381084 57953 381093 57987
rect 381093 57953 381127 57987
rect 381127 57953 381136 57987
rect 381084 57944 381136 57953
rect 387892 57876 387944 57928
rect 387984 57876 388036 57928
rect 416964 57876 417016 57928
rect 433708 57876 433760 57928
rect 466644 57876 466696 57928
rect 472164 57876 472216 57928
rect 480352 57876 480404 57928
rect 480536 57876 480588 57928
rect 298376 57808 298428 57860
rect 287244 56695 287296 56704
rect 287244 56661 287253 56695
rect 287253 56661 287287 56695
rect 287287 56661 287296 56695
rect 287244 56652 287296 56661
rect 283104 56627 283156 56636
rect 283104 56593 283113 56627
rect 283113 56593 283147 56627
rect 283147 56593 283156 56627
rect 283104 56584 283156 56593
rect 324504 56627 324556 56636
rect 324504 56593 324513 56627
rect 324513 56593 324547 56627
rect 324547 56593 324556 56627
rect 324504 56584 324556 56593
rect 375564 56584 375616 56636
rect 407764 56627 407816 56636
rect 407764 56593 407773 56627
rect 407773 56593 407807 56627
rect 407807 56593 407816 56627
rect 407764 56584 407816 56593
rect 240232 56559 240284 56568
rect 240232 56525 240241 56559
rect 240241 56525 240275 56559
rect 240275 56525 240284 56559
rect 240232 56516 240284 56525
rect 249892 56559 249944 56568
rect 249892 56525 249901 56559
rect 249901 56525 249935 56559
rect 249935 56525 249944 56559
rect 249892 56516 249944 56525
rect 281724 56516 281776 56568
rect 287244 56559 287296 56568
rect 287244 56525 287253 56559
rect 287253 56525 287287 56559
rect 287287 56525 287296 56559
rect 287244 56516 287296 56525
rect 329932 56516 329984 56568
rect 330024 56516 330076 56568
rect 353484 56516 353536 56568
rect 353668 56516 353720 56568
rect 397828 56516 397880 56568
rect 375564 56491 375616 56500
rect 375564 56457 375573 56491
rect 375573 56457 375607 56491
rect 375607 56457 375616 56491
rect 375564 56448 375616 56457
rect 255504 55267 255556 55276
rect 255504 55233 255513 55267
rect 255513 55233 255547 55267
rect 255547 55233 255556 55267
rect 255504 55224 255556 55233
rect 266820 55224 266872 55276
rect 267004 55224 267056 55276
rect 310888 55224 310940 55276
rect 298376 55156 298428 55208
rect 298468 55156 298520 55208
rect 329932 55199 329984 55208
rect 329932 55165 329941 55199
rect 329941 55165 329975 55199
rect 329975 55165 329984 55199
rect 329932 55156 329984 55165
rect 342536 55156 342588 55208
rect 367284 55156 367336 55208
rect 367376 55156 367428 55208
rect 267004 55131 267056 55140
rect 267004 55097 267013 55131
rect 267013 55097 267047 55131
rect 267047 55097 267056 55131
rect 267004 55088 267056 55097
rect 359188 53839 359240 53848
rect 359188 53805 359197 53839
rect 359197 53805 359231 53839
rect 359231 53805 359240 53839
rect 359188 53796 359240 53805
rect 272064 51756 272116 51808
rect 375656 51688 375708 51740
rect 249892 51187 249944 51196
rect 249892 51153 249901 51187
rect 249901 51153 249935 51187
rect 249935 51153 249944 51187
rect 249892 51144 249944 51153
rect 261024 51076 261076 51128
rect 305184 51144 305236 51196
rect 321744 51187 321796 51196
rect 321744 51153 321753 51187
rect 321753 51153 321787 51187
rect 321787 51153 321796 51187
rect 321744 51144 321796 51153
rect 309324 51076 309376 51128
rect 327264 51076 327316 51128
rect 382464 51076 382516 51128
rect 305092 51008 305144 51060
rect 261024 50940 261076 50992
rect 392216 51076 392268 51128
rect 408684 51076 408736 51128
rect 392124 51008 392176 51060
rect 408776 51008 408828 51060
rect 309416 50940 309468 50992
rect 327264 50940 327316 50992
rect 236368 48356 236420 48408
rect 233424 48288 233476 48340
rect 233516 48288 233568 48340
rect 236276 48288 236328 48340
rect 331496 48288 331548 48340
rect 332784 48356 332836 48408
rect 352104 48356 352156 48408
rect 359188 48356 359240 48408
rect 416872 48399 416924 48408
rect 416872 48365 416881 48399
rect 416881 48365 416915 48399
rect 416915 48365 416924 48399
rect 416872 48356 416924 48365
rect 334440 48288 334492 48340
rect 352012 48288 352064 48340
rect 382372 48331 382424 48340
rect 382372 48297 382381 48331
rect 382381 48297 382415 48331
rect 382415 48297 382424 48331
rect 382372 48288 382424 48297
rect 393136 48288 393188 48340
rect 393228 48288 393280 48340
rect 422392 48288 422444 48340
rect 422484 48288 422536 48340
rect 433616 48331 433668 48340
rect 433616 48297 433625 48331
rect 433625 48297 433659 48331
rect 433659 48297 433668 48331
rect 433616 48288 433668 48297
rect 466552 48331 466604 48340
rect 466552 48297 466561 48331
rect 466561 48297 466595 48331
rect 466595 48297 466604 48331
rect 466552 48288 466604 48297
rect 472072 48331 472124 48340
rect 472072 48297 472081 48331
rect 472081 48297 472115 48331
rect 472115 48297 472124 48331
rect 472072 48288 472124 48297
rect 332692 48220 332744 48272
rect 380992 48220 381044 48272
rect 381176 48220 381228 48272
rect 386696 48220 386748 48272
rect 386788 48220 386840 48272
rect 392124 48263 392176 48272
rect 392124 48229 392133 48263
rect 392133 48229 392167 48263
rect 392167 48229 392176 48263
rect 392124 48220 392176 48229
rect 416872 48220 416924 48272
rect 417056 48220 417108 48272
rect 400588 47175 400640 47184
rect 400588 47141 400597 47175
rect 400597 47141 400631 47175
rect 400631 47141 400640 47175
rect 400588 47132 400640 47141
rect 249892 47039 249944 47048
rect 249892 47005 249901 47039
rect 249901 47005 249935 47039
rect 249935 47005 249944 47039
rect 249892 46996 249944 47005
rect 270684 46996 270736 47048
rect 287244 47039 287296 47048
rect 287244 47005 287253 47039
rect 287253 47005 287287 47039
rect 287287 47005 287296 47039
rect 287244 46996 287296 47005
rect 292856 46996 292908 47048
rect 321744 47039 321796 47048
rect 321744 47005 321753 47039
rect 321753 47005 321787 47039
rect 321787 47005 321796 47039
rect 321744 46996 321796 47005
rect 240232 46971 240284 46980
rect 240232 46937 240241 46971
rect 240241 46937 240275 46971
rect 240275 46937 240284 46971
rect 240232 46928 240284 46937
rect 270592 46928 270644 46980
rect 271972 46971 272024 46980
rect 271972 46937 271981 46971
rect 271981 46937 272015 46971
rect 272015 46937 272024 46971
rect 271972 46928 272024 46937
rect 281632 46971 281684 46980
rect 281632 46937 281641 46971
rect 281641 46937 281675 46971
rect 281675 46937 281684 46971
rect 281632 46928 281684 46937
rect 330024 46928 330076 46980
rect 347964 46928 348016 46980
rect 348148 46928 348200 46980
rect 370044 46928 370096 46980
rect 370136 46928 370188 46980
rect 397736 46971 397788 46980
rect 397736 46937 397745 46971
rect 397745 46937 397779 46971
rect 397779 46937 397788 46971
rect 397736 46928 397788 46937
rect 451372 46928 451424 46980
rect 451648 46928 451700 46980
rect 231952 46903 232004 46912
rect 231952 46869 231961 46903
rect 231961 46869 231995 46903
rect 231995 46869 232004 46903
rect 231952 46860 232004 46869
rect 236276 46903 236328 46912
rect 236276 46869 236285 46903
rect 236285 46869 236319 46903
rect 236319 46869 236328 46903
rect 236276 46860 236328 46869
rect 244464 46903 244516 46912
rect 244464 46869 244473 46903
rect 244473 46869 244507 46903
rect 244507 46869 244516 46903
rect 244464 46860 244516 46869
rect 249892 46903 249944 46912
rect 249892 46869 249901 46903
rect 249901 46869 249935 46903
rect 249935 46869 249944 46903
rect 249892 46860 249944 46869
rect 288532 46860 288584 46912
rect 288624 46860 288676 46912
rect 309416 46860 309468 46912
rect 321652 46860 321704 46912
rect 321744 46860 321796 46912
rect 407764 46903 407816 46912
rect 407764 46869 407773 46903
rect 407773 46869 407807 46903
rect 407807 46869 407816 46903
rect 407764 46860 407816 46869
rect 255596 45568 255648 45620
rect 255780 45568 255832 45620
rect 267096 45568 267148 45620
rect 342444 45611 342496 45620
rect 342444 45577 342453 45611
rect 342453 45577 342487 45611
rect 342487 45577 342496 45611
rect 342444 45568 342496 45577
rect 356520 45611 356572 45620
rect 356520 45577 356529 45611
rect 356529 45577 356563 45611
rect 356563 45577 356572 45611
rect 356520 45568 356572 45577
rect 359096 45611 359148 45620
rect 359096 45577 359105 45611
rect 359105 45577 359139 45611
rect 359139 45577 359148 45611
rect 359096 45568 359148 45577
rect 400588 45611 400640 45620
rect 400588 45577 400597 45611
rect 400597 45577 400631 45611
rect 400631 45577 400640 45611
rect 400588 45568 400640 45577
rect 283196 45500 283248 45552
rect 292856 45543 292908 45552
rect 292856 45509 292865 45543
rect 292865 45509 292899 45543
rect 292899 45509 292908 45543
rect 292856 45500 292908 45509
rect 353576 45543 353628 45552
rect 353576 45509 353585 45543
rect 353585 45509 353619 45543
rect 353619 45509 353628 45543
rect 353576 45500 353628 45509
rect 408684 45500 408736 45552
rect 408776 45500 408828 45552
rect 400680 45475 400732 45484
rect 400680 45441 400689 45475
rect 400689 45441 400723 45475
rect 400723 45441 400732 45475
rect 400680 45432 400732 45441
rect 330024 44115 330076 44124
rect 330024 44081 330033 44115
rect 330033 44081 330067 44115
rect 330067 44081 330076 44115
rect 330024 44072 330076 44081
rect 271972 42916 272024 42968
rect 267096 42075 267148 42084
rect 267096 42041 267105 42075
rect 267105 42041 267139 42075
rect 267139 42041 267148 42075
rect 267096 42032 267148 42041
rect 332692 42032 332744 42084
rect 332876 42032 332928 42084
rect 357624 41420 357676 41472
rect 471980 41352 472032 41404
rect 472164 41352 472216 41404
rect 451372 41284 451424 41336
rect 451740 41284 451792 41336
rect 356520 40740 356572 40792
rect 267740 40332 267792 40384
rect 277308 40332 277360 40384
rect 402980 40332 403032 40384
rect 412456 40332 412508 40384
rect 252744 40171 252796 40180
rect 252744 40137 252753 40171
rect 252753 40137 252787 40171
rect 252787 40137 252796 40171
rect 252744 40128 252796 40137
rect 324504 40171 324556 40180
rect 324504 40137 324513 40171
rect 324513 40137 324547 40171
rect 324547 40137 324556 40171
rect 324504 40128 324556 40137
rect 311808 40060 311860 40112
rect 317328 40060 317380 40112
rect 521660 40060 521712 40112
rect 526444 40060 526496 40112
rect 480260 38700 480312 38752
rect 480536 38700 480588 38752
rect 376852 38632 376904 38684
rect 376944 38632 376996 38684
rect 382372 38632 382424 38684
rect 382464 38632 382516 38684
rect 472164 38607 472216 38616
rect 472164 38573 472173 38607
rect 472173 38573 472207 38607
rect 472207 38573 472216 38607
rect 472164 38564 472216 38573
rect 232044 37272 232096 37324
rect 236368 37272 236420 37324
rect 244556 37272 244608 37324
rect 249892 37315 249944 37324
rect 249892 37281 249901 37315
rect 249901 37281 249935 37315
rect 249935 37281 249944 37315
rect 249892 37272 249944 37281
rect 287244 37272 287296 37324
rect 287336 37272 287388 37324
rect 295524 37272 295576 37324
rect 295708 37272 295760 37324
rect 309324 37315 309376 37324
rect 309324 37281 309333 37315
rect 309333 37281 309367 37315
rect 309367 37281 309376 37315
rect 309324 37272 309376 37281
rect 310612 37272 310664 37324
rect 310796 37272 310848 37324
rect 331404 37272 331456 37324
rect 331496 37272 331548 37324
rect 334348 37272 334400 37324
rect 334440 37272 334492 37324
rect 352012 37272 352064 37324
rect 352104 37272 352156 37324
rect 407764 37315 407816 37324
rect 407764 37281 407773 37315
rect 407773 37281 407807 37315
rect 407807 37281 407816 37315
rect 407764 37272 407816 37281
rect 353576 37247 353628 37256
rect 353576 37213 353585 37247
rect 353585 37213 353619 37247
rect 353619 37213 353628 37247
rect 353576 37204 353628 37213
rect 400680 37179 400732 37188
rect 400680 37145 400689 37179
rect 400689 37145 400723 37179
rect 400723 37145 400732 37179
rect 400680 37136 400732 37145
rect 364616 35980 364668 36032
rect 282920 35955 282972 35964
rect 282920 35921 282929 35955
rect 282929 35921 282963 35955
rect 282963 35921 282972 35955
rect 282920 35912 282972 35921
rect 292856 35955 292908 35964
rect 292856 35921 292865 35955
rect 292865 35921 292899 35955
rect 292899 35921 292908 35955
rect 292856 35912 292908 35921
rect 347872 35912 347924 35964
rect 348148 35912 348200 35964
rect 356612 35955 356664 35964
rect 356612 35921 356621 35955
rect 356621 35921 356655 35955
rect 356655 35921 356664 35955
rect 356612 35912 356664 35921
rect 357532 35955 357584 35964
rect 357532 35921 357541 35955
rect 357541 35921 357575 35955
rect 357575 35921 357584 35955
rect 357532 35912 357584 35921
rect 364524 35912 364576 35964
rect 367376 35912 367428 35964
rect 367468 35912 367520 35964
rect 370044 35912 370096 35964
rect 370136 35912 370188 35964
rect 392216 35912 392268 35964
rect 3516 35844 3568 35896
rect 7564 35844 7616 35896
rect 232044 35844 232096 35896
rect 358912 35844 358964 35896
rect 359096 35844 359148 35896
rect 375564 35844 375616 35896
rect 375748 35844 375800 35896
rect 342444 32376 342496 32428
rect 240232 31875 240284 31884
rect 240232 31841 240241 31875
rect 240241 31841 240275 31875
rect 240275 31841 240284 31875
rect 240232 31832 240284 31841
rect 408776 31764 408828 31816
rect 416964 31764 417016 31816
rect 451740 31764 451792 31816
rect 480260 31764 480312 31816
rect 408684 31696 408736 31748
rect 416872 31696 416924 31748
rect 451648 31696 451700 31748
rect 252836 31628 252888 31680
rect 480352 31628 480404 31680
rect 472164 31195 472216 31204
rect 472164 31161 472173 31195
rect 472173 31161 472207 31195
rect 472207 31161 472216 31195
rect 472164 31152 472216 31161
rect 356612 31084 356664 31136
rect 278780 29180 278832 29232
rect 283104 29180 283156 29232
rect 466276 29180 466328 29232
rect 473268 29180 473320 29232
rect 572628 29180 572680 29232
rect 576768 29180 576820 29232
rect 261024 29044 261076 29096
rect 386788 29044 386840 29096
rect 521660 29044 521712 29096
rect 525892 29044 525944 29096
rect 244372 28976 244424 29028
rect 244556 28976 244608 29028
rect 249892 28976 249944 29028
rect 249984 28976 250036 29028
rect 260932 28976 260984 29028
rect 267096 29019 267148 29028
rect 267096 28985 267105 29019
rect 267105 28985 267139 29019
rect 267139 28985 267148 29019
rect 267096 28976 267148 28985
rect 270684 28976 270736 29028
rect 270776 28976 270828 29028
rect 272064 29019 272116 29028
rect 272064 28985 272073 29019
rect 272073 28985 272107 29019
rect 272107 28985 272116 29019
rect 272064 28976 272116 28985
rect 321652 28976 321704 29028
rect 321744 28976 321796 29028
rect 324504 29019 324556 29028
rect 324504 28985 324513 29019
rect 324513 28985 324547 29019
rect 324547 28985 324556 29019
rect 324504 28976 324556 28985
rect 381084 28976 381136 29028
rect 381176 28976 381228 29028
rect 386696 28976 386748 29028
rect 387892 28976 387944 29028
rect 388076 28976 388128 29028
rect 393136 28976 393188 29028
rect 393228 28976 393280 29028
rect 243084 28908 243136 28960
rect 243176 28908 243228 28960
rect 252836 28951 252888 28960
rect 252836 28917 252845 28951
rect 252845 28917 252879 28951
rect 252879 28917 252888 28951
rect 252836 28908 252888 28917
rect 254216 28908 254268 28960
rect 254308 28908 254360 28960
rect 259552 28908 259604 28960
rect 259736 28908 259788 28960
rect 265164 28908 265216 28960
rect 265256 28908 265308 28960
rect 266544 28908 266596 28960
rect 266636 28908 266688 28960
rect 281724 28951 281776 28960
rect 281724 28917 281733 28951
rect 281733 28917 281767 28951
rect 281767 28917 281776 28951
rect 281724 28908 281776 28917
rect 288440 28908 288492 28960
rect 288624 28908 288676 28960
rect 293960 28908 294012 28960
rect 294144 28908 294196 28960
rect 371240 28908 371292 28960
rect 371424 28908 371476 28960
rect 427912 28908 427964 28960
rect 400496 28840 400548 28892
rect 400680 28840 400732 28892
rect 422392 27616 422444 27668
rect 422484 27616 422536 27668
rect 266636 27591 266688 27600
rect 266636 27557 266645 27591
rect 266645 27557 266679 27591
rect 266679 27557 266688 27591
rect 266636 27548 266688 27557
rect 270776 27548 270828 27600
rect 318984 27591 319036 27600
rect 318984 27557 318993 27591
rect 318993 27557 319027 27591
rect 319027 27557 319036 27591
rect 318984 27548 319036 27557
rect 324504 27548 324556 27600
rect 327172 27548 327224 27600
rect 327264 27548 327316 27600
rect 331312 27548 331364 27600
rect 331404 27548 331456 27600
rect 346492 27591 346544 27600
rect 346492 27557 346501 27591
rect 346501 27557 346535 27591
rect 346535 27557 346544 27591
rect 346492 27548 346544 27557
rect 376852 27548 376904 27600
rect 377036 27548 377088 27600
rect 382372 27548 382424 27600
rect 382648 27548 382700 27600
rect 393228 27591 393280 27600
rect 393228 27557 393237 27591
rect 393237 27557 393271 27591
rect 393271 27557 393280 27591
rect 393228 27548 393280 27557
rect 407764 27591 407816 27600
rect 407764 27557 407773 27591
rect 407773 27557 407807 27591
rect 407807 27557 407816 27591
rect 407764 27548 407816 27557
rect 480352 27591 480404 27600
rect 480352 27557 480361 27591
rect 480361 27557 480395 27591
rect 480395 27557 480404 27591
rect 480352 27548 480404 27557
rect 240232 26367 240284 26376
rect 240232 26333 240241 26367
rect 240241 26333 240275 26367
rect 240275 26333 240284 26367
rect 240232 26324 240284 26333
rect 356520 26367 356572 26376
rect 356520 26333 356529 26367
rect 356529 26333 356563 26367
rect 356563 26333 356572 26367
rect 356520 26324 356572 26333
rect 231860 26299 231912 26308
rect 231860 26265 231869 26299
rect 231869 26265 231903 26299
rect 231903 26265 231912 26299
rect 231860 26256 231912 26265
rect 330116 26256 330168 26308
rect 236368 26231 236420 26240
rect 236368 26197 236377 26231
rect 236377 26197 236411 26231
rect 236411 26197 236420 26231
rect 236368 26188 236420 26197
rect 240232 26188 240284 26240
rect 347872 26231 347924 26240
rect 347872 26197 347881 26231
rect 347881 26197 347915 26231
rect 347915 26197 347924 26231
rect 347872 26188 347924 26197
rect 357532 26231 357584 26240
rect 357532 26197 357541 26231
rect 357541 26197 357575 26231
rect 357575 26197 357584 26231
rect 357532 26188 357584 26197
rect 358912 26188 358964 26240
rect 364800 26231 364852 26240
rect 364800 26197 364809 26231
rect 364809 26197 364843 26231
rect 364843 26197 364852 26231
rect 364800 26188 364852 26197
rect 392216 26231 392268 26240
rect 392216 26197 392225 26231
rect 392225 26197 392259 26231
rect 392259 26197 392268 26231
rect 392216 26188 392268 26197
rect 231768 26120 231820 26172
rect 231860 26120 231912 26172
rect 240324 26120 240376 26172
rect 359004 26120 359056 26172
rect 365720 22720 365772 22772
rect 365996 22720 366048 22772
rect 422116 22516 422168 22568
rect 422392 22516 422444 22568
rect 472164 22287 472216 22296
rect 472164 22253 472173 22287
rect 472173 22253 472207 22287
rect 472207 22253 472216 22287
rect 472164 22244 472216 22253
rect 380808 22176 380860 22228
rect 381176 22176 381228 22228
rect 277584 22108 277636 22160
rect 277492 22040 277544 22092
rect 416780 22040 416832 22092
rect 416964 22040 417016 22092
rect 244372 19388 244424 19440
rect 347964 19388 348016 19440
rect 427820 19431 427872 19440
rect 427820 19397 427829 19431
rect 427829 19397 427863 19431
rect 427863 19397 427872 19431
rect 427820 19388 427872 19397
rect 252836 19363 252888 19372
rect 252836 19329 252845 19363
rect 252845 19329 252879 19363
rect 252879 19329 252888 19363
rect 252836 19320 252888 19329
rect 260932 19320 260984 19372
rect 261024 19320 261076 19372
rect 281724 19363 281776 19372
rect 281724 19329 281733 19363
rect 281733 19329 281767 19363
rect 281767 19329 281776 19363
rect 281724 19320 281776 19329
rect 342352 19363 342404 19372
rect 342352 19329 342361 19363
rect 342361 19329 342395 19363
rect 342395 19329 342404 19363
rect 342352 19320 342404 19329
rect 472164 19363 472216 19372
rect 472164 19329 472173 19363
rect 472173 19329 472207 19363
rect 472207 19329 472216 19363
rect 472164 19320 472216 19329
rect 254308 19252 254360 19304
rect 255596 19252 255648 19304
rect 288532 19295 288584 19304
rect 288532 19261 288541 19295
rect 288541 19261 288575 19295
rect 288575 19261 288584 19295
rect 288532 19252 288584 19261
rect 305092 19295 305144 19304
rect 305092 19261 305101 19295
rect 305101 19261 305135 19295
rect 305135 19261 305144 19295
rect 305092 19252 305144 19261
rect 308036 19295 308088 19304
rect 308036 19261 308045 19295
rect 308045 19261 308079 19295
rect 308079 19261 308088 19295
rect 308036 19252 308088 19261
rect 397644 19252 397696 19304
rect 427820 19295 427872 19304
rect 427820 19261 427829 19295
rect 427829 19261 427863 19295
rect 427863 19261 427872 19295
rect 427820 19252 427872 19261
rect 266636 19227 266688 19236
rect 266636 19193 266645 19227
rect 266645 19193 266679 19227
rect 266679 19193 266688 19227
rect 266636 19184 266688 19193
rect 254308 19116 254360 19168
rect 255596 19116 255648 19168
rect 272064 18028 272116 18080
rect 270684 18003 270736 18012
rect 270684 17969 270693 18003
rect 270693 17969 270727 18003
rect 270727 17969 270736 18003
rect 270684 17960 270736 17969
rect 271972 17960 272024 18012
rect 318984 18003 319036 18012
rect 318984 17969 318993 18003
rect 318993 17969 319027 18003
rect 319027 17969 319036 18003
rect 318984 17960 319036 17969
rect 324412 18003 324464 18012
rect 324412 17969 324421 18003
rect 324421 17969 324455 18003
rect 324455 17969 324464 18003
rect 324412 17960 324464 17969
rect 346492 18003 346544 18012
rect 346492 17969 346501 18003
rect 346501 17969 346535 18003
rect 346535 17969 346544 18003
rect 346492 17960 346544 17969
rect 393228 18003 393280 18012
rect 393228 17969 393237 18003
rect 393237 17969 393271 18003
rect 393271 17969 393280 18003
rect 393228 17960 393280 17969
rect 480352 18003 480404 18012
rect 480352 17969 480361 18003
rect 480361 17969 480395 18003
rect 480395 17969 480404 18003
rect 480352 17960 480404 17969
rect 330116 17935 330168 17944
rect 330116 17901 330125 17935
rect 330125 17901 330159 17935
rect 330159 17901 330168 17935
rect 330116 17892 330168 17901
rect 334348 17935 334400 17944
rect 334348 17901 334357 17935
rect 334357 17901 334391 17935
rect 334391 17901 334400 17935
rect 334348 17892 334400 17901
rect 364800 17459 364852 17468
rect 364800 17425 364809 17459
rect 364809 17425 364843 17459
rect 364843 17425 364852 17459
rect 364800 17416 364852 17425
rect 347688 16804 347740 16856
rect 355968 16804 356020 16856
rect 514576 16736 514628 16788
rect 516048 16736 516100 16788
rect 318708 16668 318760 16720
rect 319628 16668 319680 16720
rect 334072 16668 334124 16720
rect 338120 16668 338172 16720
rect 524236 16668 524288 16720
rect 526444 16668 526496 16720
rect 236368 16643 236420 16652
rect 236368 16609 236377 16643
rect 236377 16609 236411 16643
rect 236411 16609 236420 16643
rect 236368 16600 236420 16609
rect 244280 16643 244332 16652
rect 244280 16609 244289 16643
rect 244289 16609 244323 16643
rect 244323 16609 244332 16643
rect 244280 16600 244332 16609
rect 392216 16643 392268 16652
rect 392216 16609 392225 16643
rect 392225 16609 392259 16643
rect 392259 16609 392268 16643
rect 392216 16600 392268 16609
rect 125416 16328 125468 16380
rect 292764 16328 292816 16380
rect 121368 16260 121420 16312
rect 291292 16260 291344 16312
rect 114468 16192 114520 16244
rect 287244 16192 287296 16244
rect 110328 16124 110380 16176
rect 285772 16124 285824 16176
rect 107568 16056 107620 16108
rect 284392 16056 284444 16108
rect 103428 15988 103480 16040
rect 281724 15988 281776 16040
rect 31668 15920 31720 15972
rect 245752 15920 245804 15972
rect 28908 15852 28960 15904
rect 243084 15852 243136 15904
rect 336556 15172 336608 15224
rect 336832 15172 336884 15224
rect 356336 15172 356388 15224
rect 356428 15172 356480 15224
rect 129648 15104 129700 15156
rect 295524 15104 295576 15156
rect 99288 15036 99340 15088
rect 280252 15036 280304 15088
rect 96528 14968 96580 15020
rect 278872 14968 278924 15020
rect 92388 14900 92440 14952
rect 276112 14900 276164 14952
rect 89628 14832 89680 14884
rect 274732 14832 274784 14884
rect 85488 14764 85540 14816
rect 273352 14764 273404 14816
rect 82728 14696 82780 14748
rect 270684 14696 270736 14748
rect 78588 14628 78640 14680
rect 269212 14628 269264 14680
rect 392032 14628 392084 14680
rect 392216 14628 392268 14680
rect 74448 14560 74500 14612
rect 267832 14560 267884 14612
rect 71688 14492 71740 14544
rect 265164 14492 265216 14544
rect 23388 14424 23440 14476
rect 241704 14424 241756 14476
rect 244188 14424 244240 14476
rect 354772 14424 354824 14476
rect 160008 14356 160060 14408
rect 311992 14356 312044 14408
rect 157248 14288 157300 14340
rect 309324 14288 309376 14340
rect 165528 14220 165580 14272
rect 313464 14220 313516 14272
rect 168288 14152 168340 14204
rect 316132 14152 316184 14204
rect 117228 14084 117280 14136
rect 246304 14084 246356 14136
rect 240048 14016 240100 14068
rect 352196 14016 352248 14068
rect 202788 13744 202840 13796
rect 334164 13744 334216 13796
rect 159916 13676 159968 13728
rect 310704 13676 310756 13728
rect 155868 13608 155920 13660
rect 309140 13608 309192 13660
rect 153108 13540 153160 13592
rect 307852 13540 307904 13592
rect 150348 13472 150400 13524
rect 306472 13472 306524 13524
rect 148968 13404 149020 13456
rect 151728 13336 151780 13388
rect 307944 13336 307996 13388
rect 146208 13268 146260 13320
rect 303620 13268 303672 13320
rect 144828 13200 144880 13252
rect 303712 13200 303764 13252
rect 132408 13132 132460 13184
rect 296904 13132 296956 13184
rect 19248 13064 19300 13116
rect 238852 13064 238904 13116
rect 382648 13064 382700 13116
rect 200028 12996 200080 13048
rect 331312 12996 331364 13048
rect 206928 12928 206980 12980
rect 335452 12928 335504 12980
rect 213828 12860 213880 12912
rect 339684 12860 339736 12912
rect 211068 12792 211120 12844
rect 336832 12792 336884 12844
rect 217968 12724 218020 12776
rect 340972 12724 341024 12776
rect 220728 12656 220780 12708
rect 342352 12656 342404 12708
rect 252836 12520 252888 12572
rect 293960 12495 294012 12504
rect 293960 12461 293969 12495
rect 293969 12461 294003 12495
rect 294003 12461 294012 12495
rect 293960 12452 294012 12461
rect 347964 12452 348016 12504
rect 370044 12452 370096 12504
rect 393228 12452 393280 12504
rect 400496 12452 400548 12504
rect 184848 12384 184900 12436
rect 323124 12384 323176 12436
rect 347872 12384 347924 12436
rect 369952 12384 370004 12436
rect 393044 12384 393096 12436
rect 400404 12384 400456 12436
rect 180708 12316 180760 12368
rect 321744 12316 321796 12368
rect 176568 12248 176620 12300
rect 320272 12248 320324 12300
rect 173808 12180 173860 12232
rect 317604 12180 317656 12232
rect 169668 12112 169720 12164
rect 316040 12112 316092 12164
rect 166908 12044 166960 12096
rect 314752 12044 314804 12096
rect 162768 11976 162820 12028
rect 313372 11976 313424 12028
rect 142068 11908 142120 11960
rect 302424 11908 302476 11960
rect 416964 11908 417016 11960
rect 126888 11840 126940 11892
rect 128268 11772 128320 11824
rect 295340 11772 295392 11824
rect 416964 11772 417016 11824
rect 13636 11704 13688 11756
rect 236184 11704 236236 11756
rect 252744 11747 252796 11756
rect 252744 11713 252753 11747
rect 252753 11713 252787 11747
rect 252787 11713 252796 11747
rect 252744 11704 252796 11713
rect 187608 11636 187660 11688
rect 325792 11636 325844 11688
rect 191748 11568 191800 11620
rect 327264 11568 327316 11620
rect 194508 11500 194560 11552
rect 328644 11500 328696 11552
rect 198648 11432 198700 11484
rect 331220 11432 331272 11484
rect 201500 11364 201552 11416
rect 332876 11364 332928 11416
rect 205548 11296 205600 11348
rect 143448 10956 143500 11008
rect 302332 10956 302384 11008
rect 140688 10888 140740 10940
rect 301044 10888 301096 10940
rect 124128 10820 124180 10872
rect 292580 10820 292632 10872
rect 119988 10752 120040 10804
rect 291200 10752 291252 10804
rect 117136 10684 117188 10736
rect 113088 10616 113140 10668
rect 287060 10616 287112 10668
rect 289912 10616 289964 10668
rect 367192 10616 367244 10668
rect 105176 10548 105228 10600
rect 283012 10548 283064 10600
rect 289820 10548 289872 10600
rect 367376 10548 367428 10600
rect 108764 10480 108816 10532
rect 285680 10480 285732 10532
rect 287612 10480 287664 10532
rect 365720 10480 365772 10532
rect 101588 10412 101640 10464
rect 281540 10412 281592 10464
rect 299664 10412 299716 10464
rect 379612 10412 379664 10464
rect 99196 10344 99248 10396
rect 280160 10344 280212 10396
rect 300952 10344 301004 10396
rect 383752 10344 383804 10396
rect 64788 10276 64840 10328
rect 262312 10276 262364 10328
rect 292948 10276 293000 10328
rect 378324 10276 378376 10328
rect 147588 10208 147640 10260
rect 305000 10208 305052 10260
rect 151636 10140 151688 10192
rect 306380 10140 306432 10192
rect 154488 10072 154540 10124
rect 158628 10004 158680 10056
rect 310520 10004 310572 10056
rect 161388 9936 161440 9988
rect 311900 9936 311952 9988
rect 377036 9936 377088 9988
rect 246764 9868 246816 9920
rect 356244 9868 356296 9920
rect 250352 9800 250404 9852
rect 253848 9732 253900 9784
rect 360292 9732 360344 9784
rect 249984 9664 250036 9716
rect 250076 9664 250128 9716
rect 254032 9664 254084 9716
rect 254308 9664 254360 9716
rect 255320 9664 255372 9716
rect 255596 9664 255648 9716
rect 257436 9664 257488 9716
rect 361764 9664 361816 9716
rect 375472 9664 375524 9716
rect 375748 9664 375800 9716
rect 397552 9707 397604 9716
rect 397552 9673 397561 9707
rect 397561 9673 397595 9707
rect 397595 9673 397604 9707
rect 397552 9664 397604 9673
rect 407856 9664 407908 9716
rect 422116 9664 422168 9716
rect 422392 9664 422444 9716
rect 427912 9664 427964 9716
rect 203892 9596 203944 9648
rect 333980 9596 334032 9648
rect 346492 9639 346544 9648
rect 346492 9605 346501 9639
rect 346501 9605 346535 9639
rect 346535 9605 346544 9639
rect 346492 9596 346544 9605
rect 369952 9639 370004 9648
rect 369952 9605 369961 9639
rect 369961 9605 369995 9639
rect 369995 9605 370004 9639
rect 369952 9596 370004 9605
rect 371240 9639 371292 9648
rect 371240 9605 371249 9639
rect 371249 9605 371283 9639
rect 371283 9605 371292 9639
rect 371240 9596 371292 9605
rect 393044 9639 393096 9648
rect 393044 9605 393053 9639
rect 393053 9605 393087 9639
rect 393087 9605 393096 9639
rect 393044 9596 393096 9605
rect 200396 9528 200448 9580
rect 332600 9528 332652 9580
rect 196808 9460 196860 9512
rect 193220 9392 193272 9444
rect 328736 9392 328788 9444
rect 189632 9324 189684 9376
rect 327080 9324 327132 9376
rect 186044 9256 186096 9308
rect 324412 9256 324464 9308
rect 182548 9188 182600 9240
rect 323216 9188 323268 9240
rect 178960 9120 179012 9172
rect 321560 9120 321612 9172
rect 322572 9120 322624 9172
rect 361672 9256 361724 9308
rect 327080 9188 327132 9240
rect 392032 9188 392084 9240
rect 325516 9120 325568 9172
rect 390652 9120 390704 9172
rect 175372 9052 175424 9104
rect 319076 9052 319128 9104
rect 328552 9052 328604 9104
rect 394792 9052 394844 9104
rect 171784 8984 171836 9036
rect 317696 8984 317748 9036
rect 323584 8984 323636 9036
rect 389272 8984 389324 9036
rect 132592 8916 132644 8968
rect 296812 8916 296864 8968
rect 334716 8916 334768 8968
rect 401692 8916 401744 8968
rect 210976 8848 211028 8900
rect 338212 8848 338264 8900
rect 207480 8780 207532 8832
rect 335360 8780 335412 8832
rect 214656 8712 214708 8764
rect 339776 8712 339828 8764
rect 221740 8644 221792 8696
rect 343732 8644 343784 8696
rect 218152 8576 218204 8628
rect 340880 8576 340932 8628
rect 225328 8508 225380 8560
rect 345204 8508 345256 8560
rect 228916 8440 228968 8492
rect 232504 8372 232556 8424
rect 349252 8372 349304 8424
rect 236000 8304 236052 8356
rect 350724 8304 350776 8356
rect 358912 8304 358964 8356
rect 359004 8304 359056 8356
rect 364432 8304 364484 8356
rect 364800 8304 364852 8356
rect 56416 8236 56468 8288
rect 258356 8236 258408 8288
rect 274088 8236 274140 8288
rect 52828 8168 52880 8220
rect 256792 8168 256844 8220
rect 270500 8168 270552 8220
rect 368572 8168 368624 8220
rect 49332 8100 49384 8152
rect 254032 8100 254084 8152
rect 267004 8100 267056 8152
rect 367100 8100 367152 8152
rect 44548 8032 44600 8084
rect 252652 8032 252704 8084
rect 263416 8032 263468 8084
rect 364432 8032 364484 8084
rect 40960 7964 41012 8016
rect 249984 7964 250036 8016
rect 259828 7964 259880 8016
rect 363052 7964 363104 8016
rect 37372 7896 37424 7948
rect 248512 7896 248564 7948
rect 256240 7896 256292 7948
rect 361580 7896 361632 7948
rect 33876 7828 33928 7880
rect 247224 7828 247276 7880
rect 252652 7828 252704 7880
rect 358912 7828 358964 7880
rect 30288 7760 30340 7812
rect 244280 7760 244332 7812
rect 249156 7760 249208 7812
rect 357440 7760 357492 7812
rect 26700 7692 26752 7744
rect 242900 7692 242952 7744
rect 245568 7692 245620 7744
rect 356152 7692 356204 7744
rect 8852 7624 8904 7676
rect 233332 7624 233384 7676
rect 234804 7624 234856 7676
rect 350632 7624 350684 7676
rect 4068 7556 4120 7608
rect 230664 7556 230716 7608
rect 231308 7556 231360 7608
rect 347872 7556 347924 7608
rect 351828 7556 351880 7608
rect 405832 7556 405884 7608
rect 477592 7556 477644 7608
rect 478696 7556 478748 7608
rect 87328 7488 87380 7540
rect 274640 7488 274692 7540
rect 277676 7488 277728 7540
rect 372712 7488 372764 7540
rect 90916 7420 90968 7472
rect 276020 7420 276072 7472
rect 281264 7420 281316 7472
rect 374092 7420 374144 7472
rect 94504 7352 94556 7404
rect 277492 7352 277544 7404
rect 284760 7352 284812 7404
rect 375472 7352 375524 7404
rect 138480 7284 138532 7336
rect 300860 7284 300912 7336
rect 347964 7284 348016 7336
rect 397552 7284 397604 7336
rect 141976 7216 142028 7268
rect 302516 7216 302568 7268
rect 346492 7216 346544 7268
rect 396172 7216 396224 7268
rect 224132 7148 224184 7200
rect 345112 7148 345164 7200
rect 227720 7080 227772 7132
rect 346400 7080 346452 7132
rect 238392 7012 238444 7064
rect 351920 7012 351972 7064
rect 241980 6944 242032 6996
rect 353392 6944 353444 6996
rect 163504 6808 163556 6860
rect 313556 6808 313608 6860
rect 349068 6808 349120 6860
rect 408776 6808 408828 6860
rect 83832 6740 83884 6792
rect 271880 6740 271932 6792
rect 320180 6740 320232 6792
rect 325608 6740 325660 6792
rect 386512 6740 386564 6792
rect 80244 6672 80296 6724
rect 270592 6672 270644 6724
rect 318800 6672 318852 6724
rect 380808 6672 380860 6724
rect 76656 6604 76708 6656
rect 269120 6604 269172 6656
rect 320180 6604 320232 6656
rect 385132 6604 385184 6656
rect 73068 6536 73120 6588
rect 266360 6536 266412 6588
rect 312176 6536 312228 6588
rect 389364 6536 389416 6588
rect 69480 6468 69532 6520
rect 264980 6468 265032 6520
rect 308588 6468 308640 6520
rect 387892 6468 387944 6520
rect 62396 6400 62448 6452
rect 260932 6400 260984 6452
rect 305000 6400 305052 6452
rect 386420 6400 386472 6452
rect 65984 6332 66036 6384
rect 263692 6332 263744 6384
rect 290740 6332 290792 6384
rect 378232 6332 378284 6384
rect 58808 6264 58860 6316
rect 259460 6264 259512 6316
rect 287152 6264 287204 6316
rect 55220 6196 55272 6248
rect 258264 6196 258316 6248
rect 283656 6196 283708 6248
rect 375380 6196 375432 6248
rect 379980 6196 380032 6248
rect 425152 6196 425204 6248
rect 51632 6128 51684 6180
rect 255320 6128 255372 6180
rect 279976 6128 280028 6180
rect 372804 6128 372856 6180
rect 372896 6128 372948 6180
rect 421104 6128 421156 6180
rect 167092 6060 167144 6112
rect 314568 6060 314620 6112
rect 314660 6060 314712 6112
rect 170588 5992 170640 6044
rect 317420 5992 317472 6044
rect 322940 5992 322992 6044
rect 354956 5992 355008 6044
rect 411352 5992 411404 6044
rect 174176 5924 174228 5976
rect 177764 5856 177816 5908
rect 316592 5924 316644 5976
rect 369860 5924 369912 5976
rect 318892 5856 318944 5908
rect 325332 5856 325384 5908
rect 360200 5856 360252 5908
rect 362132 5856 362184 5908
rect 415584 5856 415636 5908
rect 181352 5788 181404 5840
rect 322664 5788 322716 5840
rect 364340 5788 364392 5840
rect 369216 5788 369268 5840
rect 419632 5788 419684 5840
rect 184848 5720 184900 5772
rect 324320 5720 324372 5772
rect 188436 5652 188488 5704
rect 325700 5652 325752 5704
rect 192024 5584 192076 5636
rect 328460 5584 328512 5636
rect 195612 5516 195664 5568
rect 329840 5516 329892 5568
rect 137284 5448 137336 5500
rect 299480 5448 299532 5500
rect 315764 5448 315816 5500
rect 391940 5448 391992 5500
rect 401324 5448 401376 5500
rect 436192 5448 436244 5500
rect 133788 5380 133840 5432
rect 298100 5380 298152 5432
rect 301412 5380 301464 5432
rect 383844 5380 383896 5432
rect 397828 5380 397880 5432
rect 433616 5380 433668 5432
rect 130200 5312 130252 5364
rect 296720 5312 296772 5364
rect 297916 5312 297968 5364
rect 394240 5312 394292 5364
rect 432144 5312 432196 5364
rect 67180 5244 67232 5296
rect 263784 5244 263836 5296
rect 294328 5244 294380 5296
rect 380900 5244 380952 5296
rect 390652 5244 390704 5296
rect 430672 5244 430724 5296
rect 21916 5176 21968 5228
rect 240232 5176 240284 5228
rect 251456 5176 251508 5228
rect 358820 5176 358872 5228
rect 387064 5176 387116 5228
rect 427912 5176 427964 5228
rect 17316 5108 17368 5160
rect 237472 5108 237524 5160
rect 247960 5108 248012 5160
rect 356428 5108 356480 5160
rect 383568 5108 383620 5160
rect 426716 5108 426768 5160
rect 12440 5040 12492 5092
rect 236092 5040 236144 5092
rect 244372 5040 244424 5092
rect 354680 5040 354732 5092
rect 376392 5040 376444 5092
rect 422392 5040 422444 5092
rect 7656 4972 7708 5024
rect 233240 4972 233292 5024
rect 240784 4972 240836 5024
rect 353300 4972 353352 5024
rect 365720 4972 365772 5024
rect 416964 4972 417016 5024
rect 2872 4904 2924 4956
rect 230756 4904 230808 4956
rect 237196 4904 237248 4956
rect 350540 4904 350592 4956
rect 358544 4904 358596 4956
rect 414112 4904 414164 4956
rect 503536 4904 503588 4956
rect 529756 4904 529808 4956
rect 1676 4836 1728 4888
rect 230480 4836 230532 4888
rect 233700 4836 233752 4888
rect 349160 4836 349212 4888
rect 351368 4836 351420 4888
rect 410064 4836 410116 4888
rect 509148 4836 509200 4888
rect 540520 4836 540572 4888
rect 572 4768 624 4820
rect 229100 4768 229152 4820
rect 230112 4768 230164 4820
rect 347780 4768 347832 4820
rect 347872 4768 347924 4820
rect 408500 4768 408552 4820
rect 506296 4768 506348 4820
rect 536932 4768 536984 4820
rect 215852 4700 215904 4752
rect 339500 4700 339552 4752
rect 340696 4700 340748 4752
rect 404544 4700 404596 4752
rect 404912 4700 404964 4752
rect 437756 4700 437808 4752
rect 222936 4632 222988 4684
rect 343640 4632 343692 4684
rect 344284 4632 344336 4684
rect 405924 4632 405976 4684
rect 226524 4564 226576 4616
rect 345020 4564 345072 4616
rect 356060 4564 356112 4616
rect 362960 4564 363012 4616
rect 208676 4496 208728 4548
rect 283564 4496 283616 4548
rect 319260 4496 319312 4548
rect 393504 4496 393556 4548
rect 212264 4428 212316 4480
rect 284944 4428 284996 4480
rect 322848 4428 322900 4480
rect 394884 4428 394936 4480
rect 326436 4360 326488 4412
rect 397460 4360 397512 4412
rect 330024 4292 330076 4344
rect 399024 4292 399076 4344
rect 333612 4224 333664 4276
rect 400404 4224 400456 4276
rect 407856 4224 407908 4276
rect 124220 4156 124272 4208
rect 125416 4156 125468 4208
rect 140872 4156 140924 4208
rect 142068 4156 142120 4208
rect 150440 4156 150492 4208
rect 151636 4156 151688 4208
rect 158720 4156 158772 4208
rect 159916 4156 159968 4208
rect 209872 4156 209924 4208
rect 211068 4156 211120 4208
rect 42156 4088 42208 4140
rect 50344 4088 50396 4140
rect 57612 4088 57664 4140
rect 255964 4088 256016 4140
rect 276480 4088 276532 4140
rect 314660 4156 314712 4208
rect 337108 4156 337160 4208
rect 403072 4156 403124 4208
rect 314568 4088 314620 4140
rect 316684 4088 316736 4140
rect 321652 4088 321704 4140
rect 322756 4088 322808 4140
rect 331220 4088 331272 4140
rect 332508 4088 332560 4140
rect 346676 4088 346728 4140
rect 50528 4020 50580 4072
rect 253204 4020 253256 4072
rect 262220 4020 262272 4072
rect 322664 4020 322716 4072
rect 339500 4020 339552 4072
rect 405004 4156 405056 4208
rect 34980 3952 35032 4004
rect 46204 3952 46256 4004
rect 46940 3952 46992 4004
rect 252744 3952 252796 4004
rect 271696 3952 271748 4004
rect 283472 3952 283524 4004
rect 300308 3952 300360 4004
rect 363696 3952 363748 4004
rect 364524 3952 364576 4004
rect 366456 3952 366508 4004
rect 408408 4020 408460 4072
rect 412088 4088 412140 4140
rect 412548 4088 412600 4140
rect 414664 4088 414716 4140
rect 415676 4088 415728 4140
rect 416688 4088 416740 4140
rect 419172 4088 419224 4140
rect 420276 4088 420328 4140
rect 420368 4088 420420 4140
rect 420828 4088 420880 4140
rect 421564 4088 421616 4140
rect 422208 4088 422260 4140
rect 422760 4088 422812 4140
rect 423588 4088 423640 4140
rect 429936 4088 429988 4140
rect 430488 4088 430540 4140
rect 430580 4088 430632 4140
rect 431132 4088 431184 4140
rect 431868 4088 431920 4140
rect 433524 4088 433576 4140
rect 434628 4088 434680 4140
rect 437020 4088 437072 4140
rect 442356 4088 442408 4140
rect 451280 4088 451332 4140
rect 453396 4088 453448 4140
rect 469128 4088 469180 4140
rect 469864 4088 469916 4140
rect 470324 4088 470376 4140
rect 470784 4088 470836 4140
rect 472164 4088 472216 4140
rect 472716 4088 472768 4140
rect 473360 4088 473412 4140
rect 473912 4088 473964 4140
rect 474648 4088 474700 4140
rect 475108 4088 475160 4140
rect 478788 4088 478840 4140
rect 482284 4088 482336 4140
rect 493968 4088 494020 4140
rect 513196 4088 513248 4140
rect 517428 4088 517480 4140
rect 557172 4088 557224 4140
rect 558184 4088 558236 4140
rect 576216 4088 576268 4140
rect 410892 4020 410944 4072
rect 413376 4020 413428 4072
rect 414480 4020 414532 4072
rect 416136 4020 416188 4072
rect 438952 4020 439004 4072
rect 440608 4020 440660 4072
rect 445024 4020 445076 4072
rect 445392 4020 445444 4072
rect 451924 4020 451976 4072
rect 454868 4020 454920 4072
rect 456064 4020 456116 4072
rect 477408 4020 477460 4072
rect 479892 4020 479944 4072
rect 492588 4020 492640 4072
rect 509608 4020 509660 4072
rect 510528 4020 510580 4072
rect 518808 4020 518860 4072
rect 559564 4020 559616 4072
rect 409144 3952 409196 4004
rect 424416 3952 424468 4004
rect 427544 3952 427596 4004
rect 45744 3884 45796 3936
rect 251824 3884 251876 3936
rect 258632 3884 258684 3936
rect 322572 3884 322624 3936
rect 325240 3884 325292 3936
rect 391204 3884 391256 3936
rect 396724 3884 396776 3936
rect 400220 3884 400272 3936
rect 432420 3884 432472 3936
rect 448520 3952 448572 4004
rect 456156 3952 456208 4004
rect 462964 3952 463016 4004
rect 493876 3952 493928 4004
rect 512000 3952 512052 4004
rect 520096 3952 520148 4004
rect 561956 3952 562008 4004
rect 442264 3884 442316 3936
rect 496084 3884 496136 3936
rect 515588 3884 515640 3936
rect 520188 3884 520240 3936
rect 564348 3884 564400 3936
rect 565084 3884 565136 3936
rect 579804 3884 579856 3936
rect 38568 3816 38620 3868
rect 248420 3816 248472 3868
rect 255044 3816 255096 3868
rect 39764 3748 39816 3800
rect 249800 3748 249852 3800
rect 272892 3748 272944 3800
rect 316592 3748 316644 3800
rect 32680 3680 32732 3732
rect 245660 3680 245712 3732
rect 264612 3680 264664 3732
rect 287704 3680 287756 3732
rect 299112 3680 299164 3732
rect 300952 3680 301004 3732
rect 307392 3680 307444 3732
rect 309784 3680 309836 3732
rect 316960 3816 317012 3868
rect 327080 3816 327132 3868
rect 332416 3816 332468 3868
rect 318064 3748 318116 3800
rect 389824 3748 389876 3800
rect 400864 3816 400916 3868
rect 402520 3816 402572 3868
rect 403716 3816 403768 3868
rect 437664 3816 437716 3868
rect 448980 3816 449032 3868
rect 453304 3816 453356 3868
rect 467932 3816 467984 3868
rect 470692 3816 470744 3868
rect 482836 3816 482888 3868
rect 490564 3816 490616 3868
rect 496728 3816 496780 3868
rect 509884 3816 509936 3868
rect 520280 3816 520332 3868
rect 521568 3816 521620 3868
rect 566740 3816 566792 3868
rect 395344 3748 395396 3800
rect 399024 3748 399076 3800
rect 434812 3748 434864 3800
rect 438216 3748 438268 3800
rect 447784 3748 447836 3800
rect 459652 3748 459704 3800
rect 464344 3748 464396 3800
rect 489184 3748 489236 3800
rect 497740 3748 497792 3800
rect 500868 3748 500920 3800
rect 525064 3748 525116 3800
rect 525616 3748 525668 3800
rect 572628 3748 572680 3800
rect 325332 3680 325384 3732
rect 352564 3680 352616 3732
rect 353208 3680 353260 3732
rect 378416 3680 378468 3732
rect 385868 3680 385920 3732
rect 433340 3680 433392 3732
rect 434536 3680 434588 3732
rect 446404 3680 446456 3732
rect 450176 3680 450228 3732
rect 451188 3680 451240 3732
rect 466828 3680 466880 3732
rect 467748 3680 467800 3732
rect 485688 3680 485740 3732
rect 495348 3680 495400 3732
rect 498844 3680 498896 3732
rect 519084 3680 519136 3732
rect 522948 3680 523000 3732
rect 569040 3680 569092 3732
rect 25504 3612 25556 3664
rect 239588 3612 239640 3664
rect 240048 3612 240100 3664
rect 243176 3612 243228 3664
rect 244188 3612 244240 3664
rect 269304 3612 269356 3664
rect 289820 3612 289872 3664
rect 291936 3612 291988 3664
rect 299664 3612 299716 3664
rect 303804 3612 303856 3664
rect 382924 3612 382976 3664
rect 388260 3612 388312 3664
rect 389088 3612 389140 3664
rect 391848 3612 391900 3664
rect 408316 3612 408368 3664
rect 408592 3612 408644 3664
rect 426624 3612 426676 3664
rect 429292 3612 429344 3664
rect 443000 3612 443052 3664
rect 456984 3612 457036 3664
rect 458456 3612 458508 3664
rect 464436 3612 464488 3664
rect 484308 3612 484360 3664
rect 492956 3612 493008 3664
rect 499488 3612 499540 3664
rect 522672 3612 522724 3664
rect 524328 3612 524380 3664
rect 571432 3612 571484 3664
rect 18328 3544 18380 3596
rect 19248 3544 19300 3596
rect 19524 3544 19576 3596
rect 24124 3544 24176 3596
rect 24308 3544 24360 3596
rect 241520 3544 241572 3596
rect 275284 3544 275336 3596
rect 276664 3544 276716 3596
rect 16028 3476 16080 3528
rect 237564 3476 237616 3528
rect 241796 3476 241848 3528
rect 265808 3476 265860 3528
rect 287612 3476 287664 3528
rect 289544 3544 289596 3596
rect 296720 3544 296772 3596
rect 381544 3544 381596 3596
rect 389456 3544 389508 3596
rect 439412 3544 439464 3596
rect 455604 3544 455656 3596
rect 457260 3544 457312 3596
rect 465080 3544 465132 3596
rect 484216 3544 484268 3596
rect 494152 3544 494204 3596
rect 499396 3544 499448 3596
rect 523868 3544 523920 3596
rect 525524 3544 525576 3596
rect 289912 3476 289964 3528
rect 376024 3476 376076 3528
rect 382372 3476 382424 3528
rect 426348 3476 426400 3528
rect 428464 3476 428516 3528
rect 452476 3476 452528 3528
rect 460204 3476 460256 3528
rect 465632 3476 465684 3528
rect 466368 3476 466420 3528
rect 487068 3476 487120 3528
rect 498936 3476 498988 3528
rect 500776 3476 500828 3528
rect 526260 3476 526312 3528
rect 528468 3476 528520 3528
rect 569224 3476 569276 3528
rect 570236 3476 570288 3528
rect 573364 3544 573416 3596
rect 582196 3544 582248 3596
rect 573824 3476 573876 3528
rect 5264 3408 5316 3460
rect 10324 3408 10376 3460
rect 14832 3408 14884 3460
rect 236368 3408 236420 3460
rect 261024 3408 261076 3460
rect 356060 3408 356112 3460
rect 36176 3340 36228 3392
rect 39304 3340 39356 3392
rect 11244 3272 11296 3324
rect 17224 3272 17276 3324
rect 20720 3272 20772 3324
rect 28264 3272 28316 3324
rect 43352 3204 43404 3256
rect 54024 3272 54076 3324
rect 57244 3272 57296 3324
rect 60004 3340 60056 3392
rect 60648 3340 60700 3392
rect 63592 3340 63644 3392
rect 64788 3340 64840 3392
rect 70676 3340 70728 3392
rect 71688 3340 71740 3392
rect 61384 3272 61436 3324
rect 64788 3204 64840 3256
rect 257344 3340 257396 3392
rect 268108 3340 268160 3392
rect 278872 3340 278924 3392
rect 280068 3340 280120 3392
rect 282460 3340 282512 3392
rect 294604 3340 294656 3392
rect 295524 3340 295576 3392
rect 318800 3340 318852 3392
rect 324044 3340 324096 3392
rect 346492 3340 346544 3392
rect 353760 3340 353812 3392
rect 396632 3340 396684 3392
rect 408408 3408 408460 3460
rect 408500 3408 408552 3460
rect 409788 3408 409840 3460
rect 71872 3272 71924 3324
rect 258724 3272 258776 3324
rect 306196 3272 306248 3324
rect 325608 3272 325660 3324
rect 347964 3272 348016 3324
rect 360936 3272 360988 3324
rect 77852 3204 77904 3256
rect 78588 3204 78640 3256
rect 81440 3204 81492 3256
rect 82728 3204 82780 3256
rect 27896 3136 27948 3188
rect 28908 3136 28960 3188
rect 29092 3136 29144 3188
rect 32404 3136 32456 3188
rect 61200 3136 61252 3188
rect 66904 3136 66956 3188
rect 82636 3136 82688 3188
rect 84844 3204 84896 3256
rect 84936 3204 84988 3256
rect 85488 3204 85540 3256
rect 88524 3204 88576 3256
rect 89628 3204 89680 3256
rect 261484 3204 261536 3256
rect 288348 3204 288400 3256
rect 292948 3204 293000 3256
rect 302608 3204 302660 3256
rect 320180 3204 320232 3256
rect 328828 3204 328880 3256
rect 363604 3204 363656 3256
rect 370412 3204 370464 3256
rect 407304 3340 407356 3392
rect 409696 3340 409748 3392
rect 406108 3272 406160 3324
rect 411904 3204 411956 3256
rect 416780 3272 416832 3324
rect 417424 3272 417476 3324
rect 417976 3272 418028 3324
rect 444564 3408 444616 3460
rect 446588 3408 446640 3460
rect 459744 3408 459796 3460
rect 488356 3408 488408 3460
rect 501236 3408 501288 3460
rect 502248 3408 502300 3460
rect 528652 3408 528704 3460
rect 529848 3408 529900 3460
rect 581000 3408 581052 3460
rect 424324 3340 424376 3392
rect 425152 3340 425204 3392
rect 432328 3340 432380 3392
rect 89812 3136 89864 3188
rect 262864 3136 262916 3188
rect 285956 3136 286008 3188
rect 286968 3136 287020 3188
rect 293132 3136 293184 3188
rect 293868 3136 293920 3188
rect 309784 3136 309836 3188
rect 323584 3136 323636 3188
rect 327632 3136 327684 3188
rect 343088 3136 343140 3188
rect 381176 3136 381228 3188
rect 423956 3204 424008 3256
rect 424968 3204 425020 3256
rect 431224 3136 431276 3188
rect 441804 3272 441856 3324
rect 449164 3340 449216 3392
rect 482928 3340 482980 3392
rect 489368 3340 489420 3392
rect 492496 3340 492548 3392
rect 508412 3340 508464 3392
rect 514668 3340 514720 3392
rect 552388 3340 552440 3392
rect 556804 3340 556856 3392
rect 565544 3340 565596 3392
rect 578608 3340 578660 3392
rect 447784 3272 447836 3324
rect 448428 3272 448480 3324
rect 464436 3272 464488 3324
rect 464988 3272 465040 3324
rect 481548 3272 481600 3324
rect 486976 3272 487028 3324
rect 488448 3272 488500 3324
rect 502432 3272 502484 3324
rect 516784 3272 516836 3324
rect 451556 3204 451608 3256
rect 485044 3204 485096 3256
rect 488172 3204 488224 3256
rect 489828 3204 489880 3256
rect 504824 3204 504876 3256
rect 511816 3204 511868 3256
rect 540244 3272 540296 3324
rect 542912 3272 542964 3324
rect 547236 3272 547288 3324
rect 550088 3272 550140 3324
rect 435364 3136 435416 3188
rect 493324 3136 493376 3188
rect 496544 3136 496596 3188
rect 511908 3136 511960 3188
rect 540336 3204 540388 3256
rect 544108 3204 544160 3256
rect 545764 3204 545816 3256
rect 554780 3204 554832 3256
rect 95700 3068 95752 3120
rect 96528 3068 96580 3120
rect 10048 3000 10100 3052
rect 15844 3000 15896 3052
rect 68284 3000 68336 3052
rect 71044 3000 71096 3052
rect 93308 3000 93360 3052
rect 97264 3068 97316 3120
rect 98092 3068 98144 3120
rect 99196 3068 99248 3120
rect 102784 3068 102836 3120
rect 103428 3068 103480 3120
rect 103980 3068 104032 3120
rect 104808 3068 104860 3120
rect 106372 3068 106424 3120
rect 107568 3068 107620 3120
rect 111156 3068 111208 3120
rect 111708 3068 111760 3120
rect 96896 3000 96948 3052
rect 264244 3068 264296 3120
rect 313372 3068 313424 3120
rect 325516 3068 325568 3120
rect 335912 3068 335964 3120
rect 366364 3068 366416 3120
rect 368020 3068 368072 3120
rect 375196 3068 375248 3120
rect 79048 2932 79100 2984
rect 86132 2932 86184 2984
rect 75460 2864 75512 2916
rect 106924 2932 106976 2984
rect 100484 2864 100536 2916
rect 264336 3000 264388 3052
rect 320456 3000 320508 3052
rect 328552 3000 328604 3052
rect 338304 3000 338356 3052
rect 339408 3000 339460 3052
rect 350264 3000 350316 3052
rect 374552 3000 374604 3052
rect 378784 3000 378836 3052
rect 408592 3000 408644 3052
rect 410616 3068 410668 3120
rect 416780 3068 416832 3120
rect 416872 3068 416924 3120
rect 438124 3068 438176 3120
rect 444196 3068 444248 3120
rect 446496 3068 446548 3120
rect 501604 3068 501656 3120
rect 506020 3068 506072 3120
rect 507768 3068 507820 3120
rect 538128 3068 538180 3120
rect 545304 3136 545356 3188
rect 547144 3136 547196 3188
rect 548892 3136 548944 3188
rect 549904 3136 549956 3188
rect 558368 3272 558420 3324
rect 547696 3068 547748 3120
rect 413284 3000 413336 3052
rect 413376 3000 413428 3052
rect 506388 3000 506440 3052
rect 535736 3000 535788 3052
rect 546500 3000 546552 3052
rect 112352 2932 112404 2984
rect 113088 2932 113140 2984
rect 113548 2932 113600 2984
rect 114468 2932 114520 2984
rect 115940 2932 115992 2984
rect 116952 2932 117004 2984
rect 119436 2932 119488 2984
rect 119988 2932 120040 2984
rect 120632 2932 120684 2984
rect 121368 2932 121420 2984
rect 114744 2864 114796 2916
rect 105544 2796 105596 2848
rect 107568 2796 107620 2848
rect 266912 2932 266964 2984
rect 341892 2932 341944 2984
rect 351828 2932 351880 2984
rect 363328 2932 363380 2984
rect 371608 2932 371660 2984
rect 372528 2932 372580 2984
rect 377588 2932 377640 2984
rect 413468 2932 413520 2984
rect 427084 2932 427136 2984
rect 505008 2932 505060 2984
rect 533436 2932 533488 2984
rect 268384 2864 268436 2916
rect 384672 2864 384724 2916
rect 408592 2864 408644 2916
rect 416044 2864 416096 2916
rect 462044 2864 462096 2916
rect 466736 2864 466788 2916
rect 503720 2864 503772 2916
rect 531044 2864 531096 2916
rect 543004 2864 543056 2916
rect 551192 3068 551244 3120
rect 571984 3000 572036 3052
rect 577412 3000 577464 3052
rect 121828 2796 121880 2848
rect 269764 2796 269816 2848
rect 310980 2796 311032 2848
rect 385684 2796 385736 2848
rect 395436 2796 395488 2848
rect 420184 2796 420236 2848
rect 471520 2796 471572 2848
rect 471888 2796 471940 2848
rect 516692 2796 516744 2848
rect 527456 2796 527508 2848
rect 529204 2796 529256 2848
rect 541716 2796 541768 2848
rect 374000 1912 374052 1964
rect 375288 1912 375340 1964
rect 480352 960 480404 1012
rect 481088 960 481140 1012
rect 345480 688 345532 740
rect 346308 688 346360 740
rect 139676 552 139728 604
rect 140688 552 140740 604
rect 172980 552 173032 604
rect 173808 552 173860 604
rect 180156 552 180208 604
rect 180708 552 180760 604
rect 205088 552 205140 604
rect 205548 552 205600 604
rect 206284 552 206336 604
rect 206928 552 206980 604
rect 220544 552 220596 604
rect 220728 552 220780 604
rect 393044 595 393096 604
rect 393044 561 393053 595
rect 393053 561 393087 595
rect 393087 561 393096 595
rect 393044 552 393096 561
rect 435824 552 435876 604
rect 436008 552 436060 604
rect 453672 552 453724 604
rect 453948 552 454000 604
rect 499764 552 499816 604
rect 500132 552 500184 604
rect 506664 552 506716 604
rect 507216 552 507268 604
rect 513564 552 513616 604
rect 514392 552 514444 604
rect 520372 552 520424 604
rect 521476 552 521528 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 8114 700360 8170 700369
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 105464 700602 105492 703520
rect 137848 700670 137876 703520
rect 154132 700738 154160 703520
rect 170324 700806 170352 703520
rect 202800 700874 202828 703520
rect 218992 701010 219020 703520
rect 218980 701004 219032 701010
rect 218980 700946 219032 700952
rect 202788 700868 202840 700874
rect 202788 700810 202840 700816
rect 170312 700800 170364 700806
rect 170312 700742 170364 700748
rect 154120 700732 154172 700738
rect 154120 700674 154172 700680
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 105452 700596 105504 700602
rect 105452 700538 105504 700544
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 8114 700295 8170 700304
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 235184 699718 235212 703520
rect 267660 700194 267688 703520
rect 267648 700188 267700 700194
rect 267648 700130 267700 700136
rect 283852 699990 283880 703520
rect 283840 699984 283892 699990
rect 283840 699926 283892 699932
rect 300136 699718 300164 703520
rect 332520 699922 332548 703520
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 348804 699786 348832 703520
rect 355968 700936 356020 700942
rect 355968 700878 356020 700884
rect 353208 700256 353260 700262
rect 353208 700198 353260 700204
rect 348792 699780 348844 699786
rect 348792 699722 348844 699728
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 235920 643822 235948 699654
rect 300780 643958 300808 699654
rect 344928 696992 344980 696998
rect 344928 696934 344980 696940
rect 342168 673532 342220 673538
rect 342168 673474 342220 673480
rect 336648 650072 336700 650078
rect 336648 650014 336700 650020
rect 300768 643952 300820 643958
rect 300768 643894 300820 643900
rect 235908 643816 235960 643822
rect 235908 643758 235960 643764
rect 331036 643068 331088 643074
rect 331036 643010 331088 643016
rect 323124 643000 323176 643006
rect 3514 642968 3570 642977
rect 323124 642942 323176 642948
rect 3514 642903 3570 642912
rect 315212 642932 315264 642938
rect 3240 642524 3292 642530
rect 3240 642466 3292 642472
rect 3148 624980 3200 624986
rect 3148 624922 3200 624928
rect 3160 624889 3188 624922
rect 3146 624880 3202 624889
rect 3146 624815 3202 624824
rect 2780 610564 2832 610570
rect 2780 610506 2832 610512
rect 2792 610473 2820 610506
rect 2778 610464 2834 610473
rect 2778 610399 2834 610408
rect 3148 596080 3200 596086
rect 3146 596048 3148 596057
rect 3200 596048 3202 596057
rect 3146 595983 3202 595992
rect 3148 567588 3200 567594
rect 3148 567530 3200 567536
rect 3160 567361 3188 567530
rect 3146 567352 3202 567361
rect 3146 567287 3202 567296
rect 2780 553104 2832 553110
rect 2778 553072 2780 553081
rect 2832 553072 2834 553081
rect 2778 553007 2834 553016
rect 3252 538665 3280 642466
rect 3332 642252 3384 642258
rect 3332 642194 3384 642200
rect 3238 538656 3294 538665
rect 3238 538591 3294 538600
rect 3240 510400 3292 510406
rect 3240 510342 3292 510348
rect 3252 509969 3280 510342
rect 3238 509960 3294 509969
rect 3238 509895 3294 509904
rect 2780 496460 2832 496466
rect 2780 496402 2832 496408
rect 2792 495553 2820 496402
rect 2778 495544 2834 495553
rect 2778 495479 2834 495488
rect 3240 481296 3292 481302
rect 3240 481238 3292 481244
rect 3252 481137 3280 481238
rect 3238 481128 3294 481137
rect 3238 481063 3294 481072
rect 3148 452464 3200 452470
rect 3146 452432 3148 452441
rect 3200 452432 3202 452441
rect 3146 452367 3202 452376
rect 2780 438048 2832 438054
rect 2778 438016 2780 438025
rect 2832 438016 2834 438025
rect 2778 437951 2834 437960
rect 3240 424312 3292 424318
rect 3240 424254 3292 424260
rect 3252 423745 3280 424254
rect 3238 423736 3294 423745
rect 3238 423671 3294 423680
rect 3344 395049 3372 642194
rect 3422 638208 3478 638217
rect 3422 638143 3478 638152
rect 3330 395040 3386 395049
rect 3330 394975 3386 394984
rect 3240 380656 3292 380662
rect 3238 380624 3240 380633
rect 3292 380624 3294 380633
rect 3238 380559 3294 380568
rect 2780 366784 2832 366790
rect 2780 366726 2832 366732
rect 2792 366217 2820 366726
rect 2778 366208 2834 366217
rect 2778 366143 2834 366152
rect 3332 337544 3384 337550
rect 3330 337512 3332 337521
rect 3384 337512 3386 337521
rect 3330 337447 3386 337456
rect 3146 324320 3202 324329
rect 3146 324255 3202 324264
rect 3160 323105 3188 324255
rect 3146 323096 3202 323105
rect 3146 323031 3202 323040
rect 2780 308848 2832 308854
rect 2778 308816 2780 308825
rect 2832 308816 2834 308825
rect 2778 308751 2834 308760
rect 3332 294976 3384 294982
rect 3332 294918 3384 294924
rect 3344 294409 3372 294918
rect 3330 294400 3386 294409
rect 3330 294335 3386 294344
rect 3148 280152 3200 280158
rect 3146 280120 3148 280129
rect 3200 280120 3202 280129
rect 3146 280055 3202 280064
rect 3146 252512 3202 252521
rect 3146 252447 3202 252456
rect 3160 251297 3188 252447
rect 3146 251288 3202 251297
rect 3146 251223 3202 251232
rect 2780 237176 2832 237182
rect 2780 237118 2832 237124
rect 2792 237017 2820 237118
rect 2778 237008 2834 237017
rect 2778 236943 2834 236952
rect 3330 180704 3386 180713
rect 3330 180639 3386 180648
rect 3344 179489 3372 180639
rect 3330 179480 3386 179489
rect 3330 179415 3386 179424
rect 2780 165164 2832 165170
rect 2780 165106 2832 165112
rect 2792 165073 2820 165106
rect 2778 165064 2834 165073
rect 2778 164999 2834 165008
rect 3330 151736 3386 151745
rect 3330 151671 3386 151680
rect 3344 150793 3372 151671
rect 3330 150784 3386 150793
rect 3330 150719 3386 150728
rect 2964 122256 3016 122262
rect 2964 122198 3016 122204
rect 2976 122097 3004 122198
rect 2962 122088 3018 122097
rect 2962 122023 3018 122032
rect 3332 79212 3384 79218
rect 3332 79154 3384 79160
rect 3344 78985 3372 79154
rect 3330 78976 3386 78985
rect 3330 78911 3386 78920
rect 3436 7177 3464 638143
rect 3528 50153 3556 642903
rect 315212 642874 315264 642880
rect 296812 642864 296864 642870
rect 296812 642806 296864 642812
rect 270500 642728 270552 642734
rect 270500 642670 270552 642676
rect 5448 642660 5500 642666
rect 5448 642602 5500 642608
rect 5356 642592 5408 642598
rect 5356 642534 5408 642540
rect 5172 642388 5224 642394
rect 5172 642330 5224 642336
rect 4988 642116 5040 642122
rect 4988 642058 5040 642064
rect 4068 641980 4120 641986
rect 4068 641922 4120 641928
rect 3976 641912 4028 641918
rect 3976 641854 4028 641860
rect 3884 641844 3936 641850
rect 3884 641786 3936 641792
rect 3792 641776 3844 641782
rect 3792 641718 3844 641724
rect 3608 638988 3660 638994
rect 3608 638930 3660 638936
rect 3620 64569 3648 638930
rect 3698 638344 3754 638353
rect 3698 638279 3754 638288
rect 3712 93265 3740 638279
rect 3804 107681 3832 641718
rect 3896 136377 3924 641786
rect 3988 193905 4016 641854
rect 4080 222601 4108 641922
rect 4804 640552 4856 640558
rect 4804 640494 4856 640500
rect 4066 222592 4122 222601
rect 4066 222527 4122 222536
rect 3974 193896 4030 193905
rect 3974 193831 4030 193840
rect 4816 165170 4844 640494
rect 4894 638480 4950 638489
rect 4894 638415 4950 638424
rect 4908 237182 4936 638415
rect 5000 308854 5028 642058
rect 5078 638616 5134 638625
rect 5078 638551 5134 638560
rect 5092 366790 5120 638551
rect 5184 496466 5212 642330
rect 5262 638752 5318 638761
rect 5262 638687 5318 638696
rect 5172 496460 5224 496466
rect 5172 496402 5224 496408
rect 5276 438054 5304 638687
rect 5368 553110 5396 642534
rect 5460 610570 5488 642602
rect 8024 642456 8076 642462
rect 8024 642398 8076 642404
rect 7932 642320 7984 642326
rect 7932 642262 7984 642268
rect 6368 642184 6420 642190
rect 6368 642126 6420 642132
rect 6276 642048 6328 642054
rect 6276 641990 6328 641996
rect 6184 640484 6236 640490
rect 6184 640426 6236 640432
rect 5448 610564 5500 610570
rect 5448 610506 5500 610512
rect 5356 553104 5408 553110
rect 5356 553046 5408 553052
rect 5264 438048 5316 438054
rect 5264 437990 5316 437996
rect 5080 366784 5132 366790
rect 5080 366726 5132 366732
rect 4988 308848 5040 308854
rect 4988 308790 5040 308796
rect 4896 237176 4948 237182
rect 4896 237118 4948 237124
rect 4804 165164 4856 165170
rect 4804 165106 4856 165112
rect 3882 136368 3938 136377
rect 3882 136303 3938 136312
rect 6196 122262 6224 640426
rect 6288 280158 6316 641990
rect 6380 380662 6408 642126
rect 7840 640688 7892 640694
rect 7840 640630 7892 640636
rect 7748 640620 7800 640626
rect 7748 640562 7800 640568
rect 7656 640416 7708 640422
rect 7656 640358 7708 640364
rect 7564 640348 7616 640354
rect 7564 640290 7616 640296
rect 6736 639260 6788 639266
rect 6736 639202 6788 639208
rect 6644 639192 6696 639198
rect 6644 639134 6696 639140
rect 6552 639124 6604 639130
rect 6552 639066 6604 639072
rect 6460 639056 6512 639062
rect 6460 638998 6512 639004
rect 6472 452470 6500 638998
rect 6564 510406 6592 639066
rect 6656 567594 6684 639134
rect 6748 624986 6776 639202
rect 6918 638480 6974 638489
rect 6918 638415 6974 638424
rect 6932 638081 6960 638415
rect 6918 638072 6974 638081
rect 6918 638007 6974 638016
rect 6736 624980 6788 624986
rect 6736 624922 6788 624928
rect 6644 567588 6696 567594
rect 6644 567530 6696 567536
rect 6552 510400 6604 510406
rect 6552 510342 6604 510348
rect 6460 452464 6512 452470
rect 6460 452406 6512 452412
rect 6368 380656 6420 380662
rect 6368 380598 6420 380604
rect 6276 280152 6328 280158
rect 6276 280094 6328 280100
rect 6184 122256 6236 122262
rect 6184 122198 6236 122204
rect 3790 107672 3846 107681
rect 3790 107607 3846 107616
rect 3698 93256 3754 93265
rect 3698 93191 3754 93200
rect 3606 64560 3662 64569
rect 3606 64495 3662 64504
rect 3514 50144 3570 50153
rect 3514 50079 3570 50088
rect 7576 35902 7604 640290
rect 7668 79218 7696 640358
rect 7760 294982 7788 640562
rect 7852 337550 7880 640630
rect 7944 424318 7972 642262
rect 8036 481302 8064 642398
rect 265164 640756 265216 640762
rect 265164 640698 265216 640704
rect 265176 639948 265204 640698
rect 270512 639948 270540 642670
rect 288898 642016 288954 642025
rect 288898 641951 288954 641960
rect 286232 640892 286284 640898
rect 286232 640834 286284 640840
rect 278320 640824 278372 640830
rect 278320 640766 278372 640772
rect 278332 639948 278360 640766
rect 286244 639948 286272 640834
rect 288912 639948 288940 641951
rect 294144 640960 294196 640966
rect 294144 640902 294196 640908
rect 294156 639948 294184 640902
rect 296824 639948 296852 642806
rect 309968 642796 310020 642802
rect 309968 642738 310020 642744
rect 302056 641028 302108 641034
rect 302056 640970 302108 640976
rect 302068 639948 302096 640970
rect 309980 639948 310008 642738
rect 312544 641096 312596 641102
rect 312544 641038 312596 641044
rect 312556 639948 312584 641038
rect 315224 639948 315252 642874
rect 317786 642832 317842 642841
rect 317786 642767 317842 642776
rect 317800 639948 317828 642767
rect 320456 641164 320508 641170
rect 320456 641106 320508 641112
rect 320468 639948 320496 641106
rect 323136 639948 323164 642942
rect 331048 639948 331076 643010
rect 336660 639962 336688 650014
rect 342180 640098 342208 673474
rect 344940 640098 344968 696934
rect 347688 685908 347740 685914
rect 347688 685850 347740 685856
rect 347700 640098 347728 685850
rect 349436 643748 349488 643754
rect 349436 643690 349488 643696
rect 341812 640070 342208 640098
rect 344572 640070 344968 640098
rect 347148 640070 347728 640098
rect 341812 639962 341840 640070
rect 344572 639962 344600 640070
rect 347148 639962 347176 640070
rect 336306 639934 336688 639962
rect 341550 639934 341840 639962
rect 344218 639934 344600 639962
rect 346794 639934 347176 639962
rect 349448 639948 349476 643690
rect 353220 640098 353248 700198
rect 355980 640098 356008 700878
rect 362868 700120 362920 700126
rect 362868 700062 362920 700068
rect 360108 700052 360160 700058
rect 360108 699994 360160 700000
rect 357348 643884 357400 643890
rect 357348 643826 357400 643832
rect 352576 640070 353248 640098
rect 355336 640070 356008 640098
rect 352576 639962 352604 640070
rect 355336 639962 355364 640070
rect 352038 639934 352604 639962
rect 354706 639934 355364 639962
rect 357360 639948 357388 643826
rect 360120 639962 360148 699994
rect 362880 639962 362908 700062
rect 364996 699718 365024 703520
rect 393320 701004 393372 701010
rect 393320 700946 393372 700952
rect 390560 700868 390612 700874
rect 390560 700810 390612 700816
rect 383660 700188 383712 700194
rect 383660 700130 383712 700136
rect 375380 699916 375432 699922
rect 375380 699858 375432 699864
rect 371148 699848 371200 699854
rect 371148 699790 371200 699796
rect 364984 699712 365036 699718
rect 364984 699654 365036 699660
rect 365628 699712 365680 699718
rect 365628 699654 365680 699660
rect 368388 699712 368440 699718
rect 368388 699654 368440 699660
rect 365168 644020 365220 644026
rect 365168 643962 365220 643968
rect 359950 639934 360148 639962
rect 362618 639934 362908 639962
rect 365180 639948 365208 643962
rect 365640 643142 365668 699654
rect 365628 643136 365680 643142
rect 365628 643078 365680 643084
rect 333888 639872 333940 639878
rect 325726 639810 326016 639826
rect 333638 639820 333888 639826
rect 368400 639826 368428 699654
rect 371160 639826 371188 699790
rect 373080 643136 373132 643142
rect 373080 643078 373132 643084
rect 373092 639948 373120 643078
rect 375392 639962 375420 699858
rect 378140 699780 378192 699786
rect 378140 699722 378192 699728
rect 378152 639962 378180 699722
rect 380992 643952 381044 643958
rect 380992 643894 381044 643900
rect 375392 639934 375774 639962
rect 378152 639934 378350 639962
rect 381004 639948 381032 643894
rect 383672 639948 383700 700130
rect 385040 699984 385092 699990
rect 385040 699926 385092 699932
rect 385052 640098 385080 699926
rect 388904 643816 388956 643822
rect 388904 643758 388956 643764
rect 385052 640070 385632 640098
rect 385604 639962 385632 640070
rect 385604 639934 386262 639962
rect 388916 639948 388944 643758
rect 333638 639814 333940 639820
rect 325726 639804 326028 639810
rect 325726 639798 325976 639804
rect 333638 639798 333928 639814
rect 367862 639798 368428 639826
rect 370530 639798 371188 639826
rect 390572 639826 390600 700810
rect 393332 639962 393360 700946
rect 396080 700800 396132 700806
rect 396080 700742 396132 700748
rect 396092 639962 396120 700742
rect 397472 699718 397500 703520
rect 401600 700732 401652 700738
rect 401600 700674 401652 700680
rect 398840 700664 398892 700670
rect 398840 700606 398892 700612
rect 397460 699712 397512 699718
rect 397460 699654 397512 699660
rect 398852 640098 398880 700606
rect 398852 640070 399156 640098
rect 399128 639962 399156 640070
rect 401612 639962 401640 700674
rect 404360 700596 404412 700602
rect 404360 700538 404412 700544
rect 404372 639962 404400 700538
rect 409880 700528 409932 700534
rect 409880 700470 409932 700476
rect 407120 700460 407172 700466
rect 407120 700402 407172 700408
rect 407132 639962 407160 700402
rect 409892 639962 409920 700470
rect 411260 700392 411312 700398
rect 411260 700334 411312 700340
rect 393332 639934 394174 639962
rect 396092 639934 396842 639962
rect 399128 639934 399418 639962
rect 401612 639934 402086 639962
rect 404372 639934 404662 639962
rect 407132 639934 407330 639962
rect 409892 639934 409998 639962
rect 411272 639826 411300 700334
rect 413664 699854 413692 703520
rect 414018 700360 414074 700369
rect 414018 700295 414074 700304
rect 416780 700324 416832 700330
rect 413652 699848 413704 699854
rect 413652 699790 413704 699796
rect 414032 639826 414060 700295
rect 416780 700266 416832 700272
rect 416792 639826 416820 700266
rect 429856 688634 429884 703520
rect 462332 700058 462360 703520
rect 478524 700126 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700120 478564 700126
rect 478512 700062 478564 700068
rect 462320 700052 462372 700058
rect 462320 699994 462372 700000
rect 429384 688628 429436 688634
rect 429384 688570 429436 688576
rect 429844 688628 429896 688634
rect 429844 688570 429896 688576
rect 429396 685930 429424 688570
rect 494900 686089 494928 703446
rect 527192 700262 527220 703520
rect 543476 700942 543504 703520
rect 543464 700936 543516 700942
rect 543464 700878 543516 700884
rect 527180 700256 527232 700262
rect 527180 700198 527232 700204
rect 559668 688634 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 559104 688628 559156 688634
rect 559104 688570 559156 688576
rect 559656 688628 559708 688634
rect 559656 688570 559708 688576
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 429304 685902 429424 685930
rect 494242 685944 494298 685953
rect 429304 684486 429332 685902
rect 559116 685930 559144 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 494242 685879 494298 685888
rect 559024 685902 559144 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 429292 684480 429344 684486
rect 429292 684422 429344 684428
rect 419540 681760 419592 681766
rect 419540 681702 419592 681708
rect 419552 639826 419580 681702
rect 494256 678994 494284 685879
rect 559024 684486 559052 685902
rect 580172 685850 580224 685856
rect 559012 684480 559064 684486
rect 559012 684422 559064 684428
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 425060 667956 425112 667962
rect 425060 667898 425112 667904
rect 422300 652792 422352 652798
rect 422300 652734 422352 652740
rect 422312 639826 422340 652734
rect 425072 639826 425100 667898
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 429672 659682 429700 666538
rect 429488 659654 429700 659682
rect 494164 659682 494192 666538
rect 559392 659682 559420 666538
rect 494164 659654 494284 659682
rect 429488 656878 429516 659654
rect 429476 656872 429528 656878
rect 429476 656814 429528 656820
rect 494256 654158 494284 659654
rect 559208 659654 559420 659682
rect 559208 656878 559236 659654
rect 559196 656872 559248 656878
rect 559196 656814 559248 656820
rect 494060 654152 494112 654158
rect 494244 654152 494296 654158
rect 494112 654100 494244 654106
rect 494060 654094 494296 654100
rect 494072 654078 494284 654094
rect 429568 647284 429620 647290
rect 429568 647226 429620 647232
rect 429580 644026 429608 647226
rect 429568 644020 429620 644026
rect 429568 643962 429620 643968
rect 494256 643890 494284 654078
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 559288 647284 559340 647290
rect 559288 647226 559340 647232
rect 494244 643884 494296 643890
rect 494244 643826 494296 643832
rect 559300 643754 559328 647226
rect 559288 643748 559340 643754
rect 559288 643690 559340 643696
rect 530400 643068 530452 643074
rect 530400 643010 530452 643016
rect 517794 642968 517850 642977
rect 517794 642903 517850 642912
rect 473082 642696 473138 642705
rect 433616 642660 433668 642666
rect 473082 642631 473138 642640
rect 433616 642602 433668 642608
rect 428108 639946 428398 639962
rect 433628 639948 433656 642602
rect 441528 642592 441580 642598
rect 441528 642534 441580 642540
rect 438860 642524 438912 642530
rect 438860 642466 438912 642472
rect 436112 639946 436310 639962
rect 438872 639948 438900 642466
rect 441540 639948 441568 642534
rect 446772 642456 446824 642462
rect 446772 642398 446824 642404
rect 443840 639946 444222 639962
rect 446784 639948 446812 642398
rect 449440 642388 449492 642394
rect 449440 642330 449492 642336
rect 449452 639948 449480 642330
rect 454684 642320 454736 642326
rect 454684 642262 454736 642268
rect 451752 639946 452042 639962
rect 454696 639948 454724 642262
rect 459928 642252 459980 642258
rect 459928 642194 459980 642200
rect 459940 639948 459968 642194
rect 465172 642184 465224 642190
rect 465172 642126 465224 642132
rect 465184 639948 465212 642126
rect 470508 642116 470560 642122
rect 470508 642058 470560 642064
rect 467840 640688 467892 640694
rect 467840 640630 467892 640636
rect 467852 639948 467880 640630
rect 470520 639948 470548 642058
rect 473096 639948 473124 642631
rect 478326 642560 478382 642569
rect 478326 642495 478382 642504
rect 475752 640620 475804 640626
rect 475752 640562 475804 640568
rect 475764 639948 475792 640562
rect 478340 639948 478368 642495
rect 483662 642424 483718 642433
rect 483662 642359 483718 642368
rect 480996 642048 481048 642054
rect 480996 641990 481048 641996
rect 481008 639948 481036 641990
rect 483676 639948 483704 642359
rect 491482 642288 491538 642297
rect 491482 642223 491538 642232
rect 486240 641980 486292 641986
rect 486240 641922 486292 641928
rect 486252 639948 486280 641922
rect 491496 639948 491524 642223
rect 494150 642152 494206 642161
rect 494150 642087 494206 642096
rect 494164 639948 494192 642087
rect 496820 641912 496872 641918
rect 496820 641854 496872 641860
rect 504638 641880 504694 641889
rect 496832 639948 496860 641854
rect 502064 641844 502116 641850
rect 504638 641815 504694 641824
rect 502064 641786 502116 641792
rect 499396 640552 499448 640558
rect 499396 640494 499448 640500
rect 499408 639948 499436 640494
rect 502076 639948 502104 641786
rect 504652 639948 504680 641815
rect 512552 641776 512604 641782
rect 512552 641718 512604 641724
rect 507308 640484 507360 640490
rect 507308 640426 507360 640432
rect 507320 639948 507348 640426
rect 512564 639948 512592 641718
rect 515220 640416 515272 640422
rect 515220 640358 515272 640364
rect 515232 639948 515260 640358
rect 517808 639948 517836 642903
rect 529572 640960 529624 640966
rect 529572 640902 529624 640908
rect 529480 640892 529532 640898
rect 529480 640834 529532 640840
rect 523132 640348 523184 640354
rect 523132 640290 523184 640296
rect 520292 639946 520490 639962
rect 523144 639948 523172 640290
rect 428096 639940 428398 639946
rect 428148 639934 428398 639940
rect 436100 639940 436310 639946
rect 428096 639882 428148 639888
rect 436152 639934 436310 639940
rect 443828 639940 444222 639946
rect 436100 639882 436152 639888
rect 443880 639934 444222 639940
rect 451740 639940 452042 639946
rect 443828 639882 443880 639888
rect 451792 639934 452042 639940
rect 520280 639940 520490 639946
rect 451740 639882 451792 639888
rect 520332 639934 520490 639940
rect 520280 639882 520332 639888
rect 390572 639798 391506 639826
rect 411272 639798 412574 639826
rect 414032 639798 415242 639826
rect 416792 639798 417818 639826
rect 419552 639798 420486 639826
rect 422312 639798 423154 639826
rect 425072 639798 425730 639826
rect 325976 639746 326028 639752
rect 328460 639736 328512 639742
rect 307326 639674 307616 639690
rect 328460 639678 328512 639684
rect 338028 639736 338080 639742
rect 339224 639736 339276 639742
rect 338028 639678 338080 639684
rect 338882 639684 339224 639690
rect 338882 639678 339276 639684
rect 398102 639704 398158 639713
rect 307326 639668 307628 639674
rect 307326 639662 307576 639668
rect 307576 639610 307628 639616
rect 299480 639600 299532 639606
rect 291502 639538 291792 639554
rect 299414 639548 299480 639554
rect 299414 639542 299532 639548
rect 291502 639532 291804 639538
rect 291502 639526 291752 639532
rect 299414 639526 299520 639542
rect 291752 639474 291804 639480
rect 284024 639464 284076 639470
rect 275770 639402 275968 639418
rect 283682 639412 284024 639418
rect 328472 639418 328500 639678
rect 283682 639406 284076 639412
rect 275770 639396 275980 639402
rect 275770 639390 275928 639396
rect 283682 639390 284064 639406
rect 328394 639390 328500 639418
rect 275928 639338 275980 639344
rect 268200 639328 268252 639334
rect 231398 639296 231454 639305
rect 231058 639254 231398 639282
rect 233974 639296 234030 639305
rect 233634 639254 233974 639282
rect 231398 639231 231454 639240
rect 236550 639296 236606 639305
rect 236302 639254 236550 639282
rect 233974 639231 234030 639240
rect 239126 639296 239182 639305
rect 238878 639254 239126 639282
rect 236550 639231 236606 639240
rect 241886 639296 241942 639305
rect 241546 639254 241886 639282
rect 239126 639231 239182 639240
rect 241886 639231 241942 639240
rect 244002 639296 244058 639305
rect 246946 639296 247002 639305
rect 244058 639254 244214 639282
rect 246790 639254 246946 639282
rect 244002 639231 244058 639240
rect 246946 639231 247002 639240
rect 249154 639296 249210 639305
rect 252282 639296 252338 639305
rect 249210 639254 249458 639282
rect 252034 639254 252282 639282
rect 249154 639231 249210 639240
rect 254950 639296 255006 639305
rect 254702 639254 254950 639282
rect 252282 639231 252338 639240
rect 257710 639296 257766 639305
rect 257370 639254 257710 639282
rect 254950 639231 255006 639240
rect 260286 639296 260342 639305
rect 259946 639254 260286 639282
rect 257710 639231 257766 639240
rect 262862 639296 262918 639305
rect 262614 639254 262862 639282
rect 260286 639231 260342 639240
rect 267858 639276 268200 639282
rect 338040 639305 338068 639678
rect 338882 639662 339264 639678
rect 398102 639639 398158 639648
rect 420182 639704 420238 639713
rect 420182 639639 420238 639648
rect 398116 639441 398144 639639
rect 398102 639432 398158 639441
rect 398102 639367 398158 639376
rect 420196 639305 420224 639639
rect 273166 639296 273222 639305
rect 267858 639270 268252 639276
rect 267858 639254 268240 639270
rect 273102 639254 273166 639282
rect 262862 639231 262918 639240
rect 281170 639296 281226 639305
rect 281014 639254 281170 639282
rect 273166 639231 273222 639240
rect 304906 639296 304962 639305
rect 304658 639254 304906 639282
rect 281170 639231 281226 639240
rect 304906 639231 304962 639240
rect 338026 639296 338082 639305
rect 338026 639231 338082 639240
rect 420182 639296 420238 639305
rect 420182 639231 420238 639240
rect 430762 639296 430818 639305
rect 457166 639296 457222 639305
rect 430818 639254 431066 639282
rect 430762 639231 430818 639240
rect 462318 639296 462374 639305
rect 457222 639254 457378 639282
rect 457166 639231 457222 639240
rect 488630 639296 488686 639305
rect 462374 639254 462622 639282
rect 462318 639231 462374 639240
rect 509790 639296 509846 639305
rect 488686 639254 488934 639282
rect 488630 639231 488686 639240
rect 525430 639296 525486 639305
rect 509846 639254 510002 639282
rect 509790 639231 509846 639240
rect 528098 639296 528154 639305
rect 525486 639254 525734 639282
rect 525430 639231 525486 639240
rect 528154 639254 528402 639282
rect 528098 639231 528154 639240
rect 8114 638888 8170 638897
rect 8114 638823 8170 638832
rect 17406 638888 17462 638897
rect 17406 638823 17462 638832
rect 26146 638888 26202 638897
rect 26146 638823 26202 638832
rect 36726 638888 36782 638897
rect 36726 638823 36782 638832
rect 45466 638888 45522 638897
rect 45466 638823 45522 638832
rect 56046 638888 56102 638897
rect 56046 638823 56102 638832
rect 64786 638888 64842 638897
rect 64786 638823 64842 638832
rect 75366 638888 75422 638897
rect 75366 638823 75422 638832
rect 84106 638888 84162 638897
rect 84106 638823 84162 638832
rect 94686 638888 94742 638897
rect 94686 638823 94742 638832
rect 103426 638888 103482 638897
rect 103426 638823 103482 638832
rect 114006 638888 114062 638897
rect 114006 638823 114062 638832
rect 122746 638888 122802 638897
rect 122746 638823 122802 638832
rect 133326 638888 133382 638897
rect 133326 638823 133382 638832
rect 142066 638888 142122 638897
rect 142066 638823 142122 638832
rect 152646 638888 152702 638897
rect 152646 638823 152702 638832
rect 161386 638888 161442 638897
rect 161386 638823 161442 638832
rect 171966 638888 172022 638897
rect 171966 638823 172022 638832
rect 180706 638888 180762 638897
rect 180706 638823 180762 638832
rect 191286 638888 191342 638897
rect 191286 638823 191342 638832
rect 200026 638888 200082 638897
rect 200026 638823 200082 638832
rect 210606 638888 210662 638897
rect 210606 638823 210662 638832
rect 219990 638888 220046 638897
rect 219990 638823 220046 638832
rect 8128 596086 8156 638823
rect 17222 638480 17278 638489
rect 17222 638415 17278 638424
rect 17236 638081 17264 638415
rect 17420 638081 17448 638823
rect 26160 638081 26188 638823
rect 26238 638480 26294 638489
rect 36542 638480 36598 638489
rect 26294 638438 26372 638466
rect 26238 638415 26294 638424
rect 26344 638081 26372 638438
rect 36542 638415 36598 638424
rect 36556 638081 36584 638415
rect 36740 638081 36768 638823
rect 45480 638081 45508 638823
rect 45558 638480 45614 638489
rect 55862 638480 55918 638489
rect 45614 638438 45692 638466
rect 45558 638415 45614 638424
rect 45664 638081 45692 638438
rect 55862 638415 55918 638424
rect 55876 638081 55904 638415
rect 56060 638081 56088 638823
rect 64800 638081 64828 638823
rect 64878 638480 64934 638489
rect 75182 638480 75238 638489
rect 64934 638438 65012 638466
rect 64878 638415 64934 638424
rect 64984 638081 65012 638438
rect 75182 638415 75238 638424
rect 75196 638081 75224 638415
rect 75380 638081 75408 638823
rect 84120 638081 84148 638823
rect 84198 638480 84254 638489
rect 94502 638480 94558 638489
rect 84254 638438 84332 638466
rect 84198 638415 84254 638424
rect 84304 638081 84332 638438
rect 94502 638415 94558 638424
rect 94516 638081 94544 638415
rect 94700 638081 94728 638823
rect 103440 638081 103468 638823
rect 103518 638480 103574 638489
rect 113822 638480 113878 638489
rect 103574 638438 103652 638466
rect 103518 638415 103574 638424
rect 103624 638081 103652 638438
rect 113822 638415 113878 638424
rect 113836 638081 113864 638415
rect 114020 638081 114048 638823
rect 122760 638081 122788 638823
rect 122838 638480 122894 638489
rect 133142 638480 133198 638489
rect 122894 638438 122972 638466
rect 122838 638415 122894 638424
rect 122944 638081 122972 638438
rect 133142 638415 133198 638424
rect 133156 638081 133184 638415
rect 133340 638081 133368 638823
rect 142080 638081 142108 638823
rect 142158 638480 142214 638489
rect 152462 638480 152518 638489
rect 142214 638438 142292 638466
rect 142158 638415 142214 638424
rect 142264 638081 142292 638438
rect 152462 638415 152518 638424
rect 152476 638081 152504 638415
rect 152660 638081 152688 638823
rect 161400 638081 161428 638823
rect 161478 638480 161534 638489
rect 171782 638480 171838 638489
rect 161534 638438 161612 638466
rect 161478 638415 161534 638424
rect 161584 638081 161612 638438
rect 171782 638415 171838 638424
rect 171796 638081 171824 638415
rect 171980 638081 172008 638823
rect 180720 638081 180748 638823
rect 180798 638480 180854 638489
rect 191102 638480 191158 638489
rect 180854 638438 180932 638466
rect 180798 638415 180854 638424
rect 180904 638081 180932 638438
rect 191102 638415 191158 638424
rect 191116 638081 191144 638415
rect 191300 638081 191328 638823
rect 200040 638081 200068 638823
rect 200118 638480 200174 638489
rect 210422 638480 210478 638489
rect 200174 638438 200252 638466
rect 200118 638415 200174 638424
rect 200224 638081 200252 638438
rect 210422 638415 210478 638424
rect 210436 638081 210464 638415
rect 210620 638081 210648 638823
rect 220004 638081 220032 638823
rect 220082 638480 220138 638489
rect 220082 638415 220138 638424
rect 17222 638072 17278 638081
rect 17222 638007 17278 638016
rect 17406 638072 17462 638081
rect 17406 638007 17462 638016
rect 26146 638072 26202 638081
rect 26146 638007 26202 638016
rect 26330 638072 26386 638081
rect 26330 638007 26386 638016
rect 36542 638072 36598 638081
rect 36542 638007 36598 638016
rect 36726 638072 36782 638081
rect 36726 638007 36782 638016
rect 45466 638072 45522 638081
rect 45466 638007 45522 638016
rect 45650 638072 45706 638081
rect 45650 638007 45706 638016
rect 55862 638072 55918 638081
rect 55862 638007 55918 638016
rect 56046 638072 56102 638081
rect 56046 638007 56102 638016
rect 64786 638072 64842 638081
rect 64786 638007 64842 638016
rect 64970 638072 65026 638081
rect 64970 638007 65026 638016
rect 75182 638072 75238 638081
rect 75182 638007 75238 638016
rect 75366 638072 75422 638081
rect 75366 638007 75422 638016
rect 84106 638072 84162 638081
rect 84106 638007 84162 638016
rect 84290 638072 84346 638081
rect 84290 638007 84346 638016
rect 94502 638072 94558 638081
rect 94502 638007 94558 638016
rect 94686 638072 94742 638081
rect 94686 638007 94742 638016
rect 103426 638072 103482 638081
rect 103426 638007 103482 638016
rect 103610 638072 103666 638081
rect 103610 638007 103666 638016
rect 113822 638072 113878 638081
rect 113822 638007 113878 638016
rect 114006 638072 114062 638081
rect 114006 638007 114062 638016
rect 122746 638072 122802 638081
rect 122746 638007 122802 638016
rect 122930 638072 122986 638081
rect 122930 638007 122986 638016
rect 133142 638072 133198 638081
rect 133142 638007 133198 638016
rect 133326 638072 133382 638081
rect 133326 638007 133382 638016
rect 142066 638072 142122 638081
rect 142066 638007 142122 638016
rect 142250 638072 142306 638081
rect 142250 638007 142306 638016
rect 152462 638072 152518 638081
rect 152462 638007 152518 638016
rect 152646 638072 152702 638081
rect 152646 638007 152702 638016
rect 161386 638072 161442 638081
rect 161386 638007 161442 638016
rect 161570 638072 161626 638081
rect 161570 638007 161626 638016
rect 171782 638072 171838 638081
rect 171782 638007 171838 638016
rect 171966 638072 172022 638081
rect 171966 638007 172022 638016
rect 180706 638072 180762 638081
rect 180706 638007 180762 638016
rect 180890 638072 180946 638081
rect 180890 638007 180946 638016
rect 191102 638072 191158 638081
rect 191102 638007 191158 638016
rect 191286 638072 191342 638081
rect 191286 638007 191342 638016
rect 200026 638072 200082 638081
rect 200026 638007 200082 638016
rect 200210 638072 200266 638081
rect 200210 638007 200266 638016
rect 210422 638072 210478 638081
rect 210422 638007 210478 638016
rect 210606 638072 210662 638081
rect 210606 638007 210662 638016
rect 219990 638072 220046 638081
rect 219990 638007 220046 638016
rect 220096 637945 220124 638415
rect 220082 637936 220138 637945
rect 220082 637871 220138 637880
rect 8116 596080 8168 596086
rect 8116 596022 8168 596028
rect 8024 481296 8076 481302
rect 8024 481238 8076 481244
rect 7932 424312 7984 424318
rect 7932 424254 7984 424260
rect 529492 346338 529520 640834
rect 529584 393310 529612 640902
rect 529756 639872 529808 639878
rect 529756 639814 529808 639820
rect 529664 639804 529716 639810
rect 529664 639746 529716 639752
rect 529676 580990 529704 639746
rect 529768 627910 529796 639814
rect 530306 638888 530362 638897
rect 530306 638823 530362 638832
rect 529756 627904 529808 627910
rect 529756 627846 529808 627852
rect 530320 604450 530348 638823
rect 530308 604444 530360 604450
rect 530308 604386 530360 604392
rect 530412 593366 530440 643010
rect 531228 643000 531280 643006
rect 531228 642942 531280 642948
rect 531044 642932 531096 642938
rect 531044 642874 531096 642880
rect 530768 642864 530820 642870
rect 530768 642806 530820 642812
rect 530492 641164 530544 641170
rect 530492 641106 530544 641112
rect 530400 593360 530452 593366
rect 530400 593302 530452 593308
rect 529664 580984 529716 580990
rect 529664 580926 529716 580932
rect 530504 557530 530532 641106
rect 530584 640824 530636 640830
rect 530584 640766 530636 640772
rect 530492 557524 530544 557530
rect 530492 557466 530544 557472
rect 529572 393304 529624 393310
rect 529572 393246 529624 393252
rect 529664 346384 529716 346390
rect 529492 346332 529664 346338
rect 529492 346326 529716 346332
rect 529492 346310 529704 346326
rect 240520 340190 240994 340218
rect 242360 340190 242834 340218
rect 261312 340190 261878 340218
rect 266832 340190 267306 340218
rect 283300 340190 283866 340218
rect 288820 340190 289386 340218
rect 294524 340190 294906 340218
rect 331692 340190 332258 340218
rect 334820 340190 335294 340218
rect 337212 340190 337778 340218
rect 364812 340190 365286 340218
rect 367848 340190 368414 340218
rect 370332 340190 370806 340218
rect 371528 340190 372002 340218
rect 377048 340190 377522 340218
rect 381280 340190 381846 340218
rect 388088 340190 388562 340218
rect 392320 340190 392886 340218
rect 397840 340190 398406 340218
rect 408880 340190 409354 340218
rect 457272 340190 457746 340218
rect 487738 340190 488304 340218
rect 493258 340190 493824 340218
rect 514050 340190 514616 340218
rect 229112 340054 230046 340082
rect 230492 340054 230598 340082
rect 230768 340054 231242 340082
rect 231504 340054 231794 340082
rect 71044 338088 71096 338094
rect 71044 338030 71096 338036
rect 66904 338020 66956 338026
rect 66904 337962 66956 337968
rect 57244 337952 57296 337958
rect 57244 337894 57296 337900
rect 50344 337884 50396 337890
rect 50344 337826 50396 337832
rect 46204 337816 46256 337822
rect 46204 337758 46256 337764
rect 39304 337748 39356 337754
rect 39304 337690 39356 337696
rect 32404 337680 32456 337686
rect 32404 337622 32456 337628
rect 28264 337612 28316 337618
rect 28264 337554 28316 337560
rect 7840 337544 7892 337550
rect 7840 337486 7892 337492
rect 17224 337544 17276 337550
rect 17224 337486 17276 337492
rect 15844 337408 15896 337414
rect 10322 337376 10378 337385
rect 15844 337350 15896 337356
rect 10322 337311 10378 337320
rect 7748 294976 7800 294982
rect 7748 294918 7800 294924
rect 7656 79212 7708 79218
rect 7656 79154 7708 79160
rect 3516 35896 3568 35902
rect 3514 35864 3516 35873
rect 7564 35896 7616 35902
rect 3568 35864 3570 35873
rect 7564 35838 7616 35844
rect 3514 35799 3570 35808
rect 8852 7676 8904 7682
rect 8852 7618 8904 7624
rect 4068 7608 4120 7614
rect 4068 7550 4120 7556
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4830
rect 2884 480 2912 4898
rect 4080 480 4108 7550
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 8864 480 8892 7618
rect 10336 3466 10364 337311
rect 13636 11756 13688 11762
rect 13636 11698 13688 11704
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11244 3324 11296 3330
rect 11244 3266 11296 3272
rect 10048 3052 10100 3058
rect 10048 2994 10100 3000
rect 10060 480 10088 2994
rect 11256 480 11284 3266
rect 12452 480 12480 5034
rect 13648 480 13676 11698
rect 14832 3460 14884 3466
rect 14832 3402 14884 3408
rect 14844 480 14872 3402
rect 15856 3058 15884 337350
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 16040 480 16068 3470
rect 17236 3330 17264 337486
rect 24124 337476 24176 337482
rect 24124 337418 24176 337424
rect 23388 14476 23440 14482
rect 23388 14418 23440 14424
rect 19248 13116 19300 13122
rect 19248 13058 19300 13064
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17224 3324 17276 3330
rect 17224 3266 17276 3272
rect 17328 1034 17356 5102
rect 19260 3602 19288 13058
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 19248 3596 19300 3602
rect 19248 3538 19300 3544
rect 19524 3596 19576 3602
rect 19524 3538 19576 3544
rect 17236 1006 17356 1034
rect 17236 480 17264 1006
rect 18340 480 18368 3538
rect 19536 480 19564 3538
rect 20720 3324 20772 3330
rect 20720 3266 20772 3272
rect 20732 480 20760 3266
rect 21928 480 21956 5170
rect 23400 3482 23428 14418
rect 24136 3602 24164 337418
rect 26700 7744 26752 7750
rect 26700 7686 26752 7692
rect 25504 3664 25556 3670
rect 25504 3606 25556 3612
rect 24124 3596 24176 3602
rect 24124 3538 24176 3544
rect 24308 3596 24360 3602
rect 24308 3538 24360 3544
rect 23124 3454 23428 3482
rect 23124 480 23152 3454
rect 24320 480 24348 3538
rect 25516 480 25544 3606
rect 26712 480 26740 7686
rect 28276 3330 28304 337554
rect 31668 15972 31720 15978
rect 31668 15914 31720 15920
rect 28908 15904 28960 15910
rect 28908 15846 28960 15852
rect 28264 3324 28316 3330
rect 28264 3266 28316 3272
rect 28920 3194 28948 15846
rect 30288 7812 30340 7818
rect 30288 7754 30340 7760
rect 27896 3188 27948 3194
rect 27896 3130 27948 3136
rect 28908 3188 28960 3194
rect 28908 3130 28960 3136
rect 29092 3188 29144 3194
rect 29092 3130 29144 3136
rect 27908 480 27936 3130
rect 29104 480 29132 3130
rect 30300 480 30328 7754
rect 31680 626 31708 15914
rect 32416 3194 32444 337622
rect 37372 7948 37424 7954
rect 37372 7890 37424 7896
rect 33876 7880 33928 7886
rect 33876 7822 33928 7828
rect 32680 3732 32732 3738
rect 32680 3674 32732 3680
rect 32404 3188 32456 3194
rect 32404 3130 32456 3136
rect 31496 598 31708 626
rect 31496 480 31524 598
rect 32692 480 32720 3674
rect 33888 480 33916 7822
rect 34980 4004 35032 4010
rect 34980 3946 35032 3952
rect 34992 480 35020 3946
rect 36176 3392 36228 3398
rect 36176 3334 36228 3340
rect 36188 480 36216 3334
rect 37384 480 37412 7890
rect 38568 3868 38620 3874
rect 38568 3810 38620 3816
rect 38580 480 38608 3810
rect 39316 3398 39344 337690
rect 44548 8084 44600 8090
rect 44548 8026 44600 8032
rect 40960 8016 41012 8022
rect 40960 7958 41012 7964
rect 39764 3800 39816 3806
rect 39764 3742 39816 3748
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 39776 480 39804 3742
rect 40972 480 41000 7958
rect 42156 4140 42208 4146
rect 42156 4082 42208 4088
rect 42168 480 42196 4082
rect 43352 3256 43404 3262
rect 43352 3198 43404 3204
rect 43364 480 43392 3198
rect 44560 480 44588 8026
rect 46216 4010 46244 337758
rect 49332 8152 49384 8158
rect 49332 8094 49384 8100
rect 48134 6216 48190 6225
rect 48134 6151 48190 6160
rect 46204 4004 46256 4010
rect 46204 3946 46256 3952
rect 46940 4004 46992 4010
rect 46940 3946 46992 3952
rect 45744 3936 45796 3942
rect 45744 3878 45796 3884
rect 45756 480 45784 3878
rect 46952 480 46980 3946
rect 48148 480 48176 6151
rect 49344 480 49372 8094
rect 50356 4146 50384 337826
rect 56416 8288 56468 8294
rect 56416 8230 56468 8236
rect 52828 8220 52880 8226
rect 52828 8162 52880 8168
rect 51632 6180 51684 6186
rect 51632 6122 51684 6128
rect 50344 4140 50396 4146
rect 50344 4082 50396 4088
rect 50528 4072 50580 4078
rect 50528 4014 50580 4020
rect 50540 480 50568 4014
rect 51644 480 51672 6122
rect 52840 480 52868 8162
rect 55220 6248 55272 6254
rect 55220 6190 55272 6196
rect 54024 3324 54076 3330
rect 54024 3266 54076 3272
rect 54036 480 54064 3266
rect 55232 480 55260 6190
rect 56428 480 56456 8230
rect 57256 3330 57284 337894
rect 61384 337340 61436 337346
rect 61384 337282 61436 337288
rect 60646 10296 60702 10305
rect 60646 10231 60702 10240
rect 58808 6316 58860 6322
rect 58808 6258 58860 6264
rect 57612 4140 57664 4146
rect 57612 4082 57664 4088
rect 57244 3324 57296 3330
rect 57244 3266 57296 3272
rect 57624 480 57652 4082
rect 58820 480 58848 6258
rect 60660 3398 60688 10231
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60016 480 60044 3334
rect 61396 3330 61424 337282
rect 64788 10328 64840 10334
rect 64788 10270 64840 10276
rect 62396 6452 62448 6458
rect 62396 6394 62448 6400
rect 61384 3324 61436 3330
rect 61384 3266 61436 3272
rect 61200 3188 61252 3194
rect 61200 3130 61252 3136
rect 61212 480 61240 3130
rect 62408 480 62436 6394
rect 64800 3398 64828 10270
rect 65984 6384 66036 6390
rect 65984 6326 66036 6332
rect 63592 3392 63644 3398
rect 63592 3334 63644 3340
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 63604 480 63632 3334
rect 64788 3256 64840 3262
rect 64788 3198 64840 3204
rect 64800 480 64828 3198
rect 65996 480 66024 6326
rect 66916 3194 66944 337962
rect 69480 6520 69532 6526
rect 69480 6462 69532 6468
rect 67180 5296 67232 5302
rect 67180 5238 67232 5244
rect 66904 3188 66956 3194
rect 66904 3130 66956 3136
rect 67192 480 67220 5238
rect 68284 3052 68336 3058
rect 68284 2994 68336 3000
rect 68296 480 68324 2994
rect 69492 480 69520 6462
rect 70676 3392 70728 3398
rect 70676 3334 70728 3340
rect 70688 480 70716 3334
rect 71056 3058 71084 338030
rect 228180 337544 228232 337550
rect 228180 337486 228232 337492
rect 228192 337414 228220 337486
rect 228180 337408 228232 337414
rect 228180 337350 228232 337356
rect 84844 337272 84896 337278
rect 84844 337214 84896 337220
rect 82728 14748 82780 14754
rect 82728 14690 82780 14696
rect 78588 14680 78640 14686
rect 78588 14622 78640 14628
rect 74448 14612 74500 14618
rect 74448 14554 74500 14560
rect 71688 14544 71740 14550
rect 71688 14486 71740 14492
rect 71700 3398 71728 14486
rect 73068 6588 73120 6594
rect 73068 6530 73120 6536
rect 71688 3392 71740 3398
rect 71688 3334 71740 3340
rect 71872 3324 71924 3330
rect 71872 3266 71924 3272
rect 71044 3052 71096 3058
rect 71044 2994 71096 3000
rect 71884 480 71912 3266
rect 73080 480 73108 6530
rect 74460 3380 74488 14554
rect 76656 6656 76708 6662
rect 76656 6598 76708 6604
rect 74276 3352 74488 3380
rect 74276 480 74304 3352
rect 75460 2916 75512 2922
rect 75460 2858 75512 2864
rect 75472 480 75500 2858
rect 76668 480 76696 6598
rect 78600 3262 78628 14622
rect 80244 6724 80296 6730
rect 80244 6666 80296 6672
rect 77852 3256 77904 3262
rect 77852 3198 77904 3204
rect 78588 3256 78640 3262
rect 78588 3198 78640 3204
rect 77864 480 77892 3198
rect 79048 2984 79100 2990
rect 79048 2926 79100 2932
rect 79060 480 79088 2926
rect 80256 480 80284 6666
rect 82740 3262 82768 14690
rect 83832 6792 83884 6798
rect 83832 6734 83884 6740
rect 81440 3256 81492 3262
rect 81440 3198 81492 3204
rect 82728 3256 82780 3262
rect 82728 3198 82780 3204
rect 81452 480 81480 3198
rect 82636 3188 82688 3194
rect 82636 3130 82688 3136
rect 82648 480 82676 3130
rect 83844 480 83872 6734
rect 84856 3262 84884 337214
rect 97264 337204 97316 337210
rect 97264 337146 97316 337152
rect 96528 15020 96580 15026
rect 96528 14962 96580 14968
rect 92388 14952 92440 14958
rect 92388 14894 92440 14900
rect 89628 14884 89680 14890
rect 89628 14826 89680 14832
rect 85488 14816 85540 14822
rect 85488 14758 85540 14764
rect 85500 3262 85528 14758
rect 87328 7540 87380 7546
rect 87328 7482 87380 7488
rect 84844 3256 84896 3262
rect 84844 3198 84896 3204
rect 84936 3256 84988 3262
rect 84936 3198 84988 3204
rect 85488 3256 85540 3262
rect 85488 3198 85540 3204
rect 84948 480 84976 3198
rect 86132 2984 86184 2990
rect 86132 2926 86184 2932
rect 86144 480 86172 2926
rect 87340 480 87368 7482
rect 89640 3262 89668 14826
rect 90916 7472 90968 7478
rect 90916 7414 90968 7420
rect 88524 3256 88576 3262
rect 88524 3198 88576 3204
rect 89628 3256 89680 3262
rect 89628 3198 89680 3204
rect 88536 480 88564 3198
rect 89812 3188 89864 3194
rect 89812 3130 89864 3136
rect 89824 1578 89852 3130
rect 89732 1550 89852 1578
rect 89732 480 89760 1550
rect 90928 480 90956 7414
rect 92400 3482 92428 14894
rect 94504 7404 94556 7410
rect 94504 7346 94556 7352
rect 92124 3454 92428 3482
rect 92124 480 92152 3454
rect 93308 3052 93360 3058
rect 93308 2994 93360 3000
rect 93320 480 93348 2994
rect 94516 480 94544 7346
rect 96540 3126 96568 14962
rect 97276 3126 97304 337146
rect 104808 337136 104860 337142
rect 104808 337078 104860 337084
rect 103428 16040 103480 16046
rect 103428 15982 103480 15988
rect 99288 15088 99340 15094
rect 99288 15030 99340 15036
rect 99196 10396 99248 10402
rect 99196 10338 99248 10344
rect 99208 3126 99236 10338
rect 95700 3120 95752 3126
rect 95700 3062 95752 3068
rect 96528 3120 96580 3126
rect 96528 3062 96580 3068
rect 97264 3120 97316 3126
rect 97264 3062 97316 3068
rect 98092 3120 98144 3126
rect 98092 3062 98144 3068
rect 99196 3120 99248 3126
rect 99196 3062 99248 3068
rect 95712 480 95740 3062
rect 96896 3052 96948 3058
rect 96896 2994 96948 3000
rect 96908 480 96936 2994
rect 98104 480 98132 3062
rect 99300 480 99328 15030
rect 101588 10464 101640 10470
rect 101588 10406 101640 10412
rect 100484 2916 100536 2922
rect 100484 2858 100536 2864
rect 100496 480 100524 2858
rect 101600 480 101628 10406
rect 103440 3126 103468 15982
rect 104820 3126 104848 337078
rect 111708 337068 111760 337074
rect 111708 337010 111760 337016
rect 105544 336864 105596 336870
rect 105544 336806 105596 336812
rect 105176 10600 105228 10606
rect 105176 10542 105228 10548
rect 102784 3120 102836 3126
rect 102784 3062 102836 3068
rect 103428 3120 103480 3126
rect 103428 3062 103480 3068
rect 103980 3120 104032 3126
rect 103980 3062 104032 3068
rect 104808 3120 104860 3126
rect 104808 3062 104860 3068
rect 102796 480 102824 3062
rect 103992 480 104020 3062
rect 105188 480 105216 10542
rect 105556 2854 105584 336806
rect 106924 336796 106976 336802
rect 106924 336738 106976 336744
rect 106372 3120 106424 3126
rect 106372 3062 106424 3068
rect 105544 2848 105596 2854
rect 105544 2790 105596 2796
rect 106384 480 106412 3062
rect 106936 2990 106964 336738
rect 110328 16176 110380 16182
rect 110328 16118 110380 16124
rect 107568 16108 107620 16114
rect 107568 16050 107620 16056
rect 107580 3126 107608 16050
rect 108764 10532 108816 10538
rect 108764 10474 108816 10480
rect 107568 3120 107620 3126
rect 107568 3062 107620 3068
rect 106924 2984 106976 2990
rect 106924 2926 106976 2932
rect 107568 2848 107620 2854
rect 107568 2790 107620 2796
rect 107580 480 107608 2790
rect 108776 480 108804 10474
rect 110340 3346 110368 16118
rect 109972 3318 110368 3346
rect 109972 480 110000 3318
rect 111720 3126 111748 337010
rect 118608 337000 118660 337006
rect 118608 336942 118660 336948
rect 114468 16244 114520 16250
rect 114468 16186 114520 16192
rect 113088 10668 113140 10674
rect 113088 10610 113140 10616
rect 111156 3120 111208 3126
rect 111156 3062 111208 3068
rect 111708 3120 111760 3126
rect 111708 3062 111760 3068
rect 111168 480 111196 3062
rect 113100 2990 113128 10610
rect 114480 2990 114508 16186
rect 117228 14136 117280 14142
rect 117228 14078 117280 14084
rect 117136 10736 117188 10742
rect 117136 10678 117188 10684
rect 117148 3618 117176 10678
rect 116964 3590 117176 3618
rect 116964 2990 116992 3590
rect 117240 3482 117268 14078
rect 117148 3454 117268 3482
rect 112352 2984 112404 2990
rect 112352 2926 112404 2932
rect 113088 2984 113140 2990
rect 113088 2926 113140 2932
rect 113548 2984 113600 2990
rect 113548 2926 113600 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 115940 2984 115992 2990
rect 115940 2926 115992 2932
rect 116952 2984 117004 2990
rect 116952 2926 117004 2932
rect 112364 480 112392 2926
rect 113560 480 113588 2926
rect 114744 2916 114796 2922
rect 114744 2858 114796 2864
rect 114756 480 114784 2858
rect 115952 480 115980 2926
rect 117148 480 117176 3454
rect 118620 3346 118648 336942
rect 125508 336932 125560 336938
rect 125508 336874 125560 336880
rect 125416 16380 125468 16386
rect 125416 16322 125468 16328
rect 121368 16312 121420 16318
rect 121368 16254 121420 16260
rect 119988 10804 120040 10810
rect 119988 10746 120040 10752
rect 118252 3318 118648 3346
rect 118252 480 118280 3318
rect 120000 2990 120028 10746
rect 121380 2990 121408 16254
rect 124128 10872 124180 10878
rect 124128 10814 124180 10820
rect 124140 3482 124168 10814
rect 125428 4214 125456 16322
rect 124220 4208 124272 4214
rect 124220 4150 124272 4156
rect 125416 4208 125468 4214
rect 125416 4150 125468 4156
rect 123036 3454 124168 3482
rect 119436 2984 119488 2990
rect 119436 2926 119488 2932
rect 119988 2984 120040 2990
rect 119988 2926 120040 2932
rect 120632 2984 120684 2990
rect 120632 2926 120684 2932
rect 121368 2984 121420 2990
rect 121368 2926 121420 2932
rect 119448 480 119476 2926
rect 120644 480 120672 2926
rect 121828 2848 121880 2854
rect 121828 2790 121880 2796
rect 121840 480 121868 2790
rect 123036 480 123064 3454
rect 124232 480 124260 4150
rect 125520 3482 125548 336874
rect 129648 15156 129700 15162
rect 129648 15098 129700 15104
rect 126888 11892 126940 11898
rect 126888 11834 126940 11840
rect 126900 3482 126928 11834
rect 128268 11824 128320 11830
rect 128268 11766 128320 11772
rect 128280 3482 128308 11766
rect 129660 3482 129688 15098
rect 160008 14408 160060 14414
rect 160008 14350 160060 14356
rect 157248 14340 157300 14346
rect 157248 14282 157300 14288
rect 155868 13660 155920 13666
rect 155868 13602 155920 13608
rect 153108 13592 153160 13598
rect 153108 13534 153160 13540
rect 150348 13524 150400 13530
rect 150348 13466 150400 13472
rect 148968 13456 149020 13462
rect 148968 13398 149020 13404
rect 146208 13320 146260 13326
rect 146208 13262 146260 13268
rect 144828 13252 144880 13258
rect 144828 13194 144880 13200
rect 132408 13184 132460 13190
rect 132408 13126 132460 13132
rect 130200 5364 130252 5370
rect 130200 5306 130252 5312
rect 125428 3454 125548 3482
rect 126624 3454 126928 3482
rect 127820 3454 128308 3482
rect 129016 3454 129688 3482
rect 125428 480 125456 3454
rect 126624 480 126652 3454
rect 127820 480 127848 3454
rect 129016 480 129044 3454
rect 130212 480 130240 5306
rect 132420 3482 132448 13126
rect 142068 11960 142120 11966
rect 142068 11902 142120 11908
rect 140688 10940 140740 10946
rect 140688 10882 140740 10888
rect 132592 8968 132644 8974
rect 132592 8910 132644 8916
rect 136086 8936 136142 8945
rect 131408 3454 132448 3482
rect 131408 480 131436 3454
rect 132604 480 132632 8910
rect 136086 8871 136142 8880
rect 134890 7576 134946 7585
rect 134890 7511 134946 7520
rect 133788 5432 133840 5438
rect 133788 5374 133840 5380
rect 133800 480 133828 5374
rect 134904 480 134932 7511
rect 136100 480 136128 8871
rect 138480 7336 138532 7342
rect 138480 7278 138532 7284
rect 137284 5500 137336 5506
rect 137284 5442 137336 5448
rect 137296 480 137324 5442
rect 138492 480 138520 7278
rect 140700 610 140728 10882
rect 141976 7268 142028 7274
rect 141976 7210 142028 7216
rect 140872 4208 140924 4214
rect 140872 4150 140924 4156
rect 139676 604 139728 610
rect 139676 546 139728 552
rect 140688 604 140740 610
rect 140688 546 140740 552
rect 139688 480 139716 546
rect 140884 480 140912 4150
rect 141988 3482 142016 7210
rect 142080 4214 142108 11902
rect 143448 11008 143500 11014
rect 143448 10950 143500 10956
rect 142068 4208 142120 4214
rect 142068 4150 142120 4156
rect 141988 3454 142108 3482
rect 142080 480 142108 3454
rect 143460 3346 143488 10950
rect 144840 3346 144868 13194
rect 146220 3346 146248 13262
rect 147588 10260 147640 10266
rect 147588 10202 147640 10208
rect 147600 3346 147628 10202
rect 148980 3346 149008 13398
rect 150360 3346 150388 13466
rect 151728 13388 151780 13394
rect 151728 13330 151780 13336
rect 151636 10192 151688 10198
rect 151636 10134 151688 10140
rect 151648 4214 151676 10134
rect 150440 4208 150492 4214
rect 150440 4150 150492 4156
rect 151636 4208 151688 4214
rect 151636 4150 151688 4156
rect 143276 3318 143488 3346
rect 144472 3318 144868 3346
rect 145668 3318 146248 3346
rect 146864 3318 147628 3346
rect 148060 3318 149008 3346
rect 149256 3318 150388 3346
rect 143276 480 143304 3318
rect 144472 480 144500 3318
rect 145668 480 145696 3318
rect 146864 480 146892 3318
rect 148060 480 148088 3318
rect 149256 480 149284 3318
rect 150452 480 150480 4150
rect 151740 3482 151768 13330
rect 151556 3454 151768 3482
rect 151556 480 151584 3454
rect 153120 3346 153148 13534
rect 154488 10124 154540 10130
rect 154488 10066 154540 10072
rect 154500 3346 154528 10066
rect 155880 3346 155908 13602
rect 157260 3346 157288 14282
rect 159916 13728 159968 13734
rect 159916 13670 159968 13676
rect 158628 10056 158680 10062
rect 158628 9998 158680 10004
rect 158640 3346 158668 9998
rect 159928 4214 159956 13670
rect 158720 4208 158772 4214
rect 158720 4150 158772 4156
rect 159916 4208 159968 4214
rect 159916 4150 159968 4156
rect 152752 3318 153148 3346
rect 153948 3318 154528 3346
rect 155144 3318 155908 3346
rect 156340 3318 157288 3346
rect 157536 3318 158668 3346
rect 152752 480 152780 3318
rect 153948 480 153976 3318
rect 155144 480 155172 3318
rect 156340 480 156368 3318
rect 157536 480 157564 3318
rect 158732 480 158760 4150
rect 160020 3482 160048 14350
rect 165528 14272 165580 14278
rect 165528 14214 165580 14220
rect 162768 12028 162820 12034
rect 162768 11970 162820 11976
rect 161388 9988 161440 9994
rect 161388 9930 161440 9936
rect 159928 3454 160048 3482
rect 159928 480 159956 3454
rect 161400 3346 161428 9930
rect 162780 3346 162808 11970
rect 163504 6860 163556 6866
rect 163504 6802 163556 6808
rect 161124 3318 161428 3346
rect 162320 3318 162808 3346
rect 161124 480 161152 3318
rect 162320 480 162348 3318
rect 163516 480 163544 6802
rect 165540 3346 165568 14214
rect 168288 14204 168340 14210
rect 168288 14146 168340 14152
rect 166908 12096 166960 12102
rect 166908 12038 166960 12044
rect 166920 3346 166948 12038
rect 167092 6112 167144 6118
rect 167092 6054 167144 6060
rect 164712 3318 165568 3346
rect 165908 3318 166948 3346
rect 164712 480 164740 3318
rect 165908 480 165936 3318
rect 167104 480 167132 6054
rect 168300 3482 168328 14146
rect 202788 13796 202840 13802
rect 202788 13738 202840 13744
rect 200028 13048 200080 13054
rect 200028 12990 200080 12996
rect 184848 12436 184900 12442
rect 184848 12378 184900 12384
rect 180708 12368 180760 12374
rect 180708 12310 180760 12316
rect 176568 12300 176620 12306
rect 176568 12242 176620 12248
rect 173808 12232 173860 12238
rect 173808 12174 173860 12180
rect 169668 12164 169720 12170
rect 169668 12106 169720 12112
rect 168208 3454 168328 3482
rect 168208 480 168236 3454
rect 169680 3346 169708 12106
rect 171784 9036 171836 9042
rect 171784 8978 171836 8984
rect 170588 6044 170640 6050
rect 170588 5986 170640 5992
rect 169404 3318 169708 3346
rect 169404 480 169432 3318
rect 170600 480 170628 5986
rect 171796 480 171824 8978
rect 173820 610 173848 12174
rect 175372 9104 175424 9110
rect 175372 9046 175424 9052
rect 174176 5976 174228 5982
rect 174176 5918 174228 5924
rect 172980 604 173032 610
rect 172980 546 173032 552
rect 173808 604 173860 610
rect 173808 546 173860 552
rect 172992 480 173020 546
rect 174188 480 174216 5918
rect 175384 480 175412 9046
rect 176580 480 176608 12242
rect 178960 9172 179012 9178
rect 178960 9114 179012 9120
rect 177764 5908 177816 5914
rect 177764 5850 177816 5856
rect 177776 480 177804 5850
rect 178972 480 179000 9114
rect 180720 610 180748 12310
rect 182548 9240 182600 9246
rect 182548 9182 182600 9188
rect 181352 5840 181404 5846
rect 181352 5782 181404 5788
rect 180156 604 180208 610
rect 180156 546 180208 552
rect 180708 604 180760 610
rect 180708 546 180760 552
rect 180168 480 180196 546
rect 181364 480 181392 5782
rect 182560 480 182588 9182
rect 184860 5930 184888 12378
rect 187608 11688 187660 11694
rect 187608 11630 187660 11636
rect 186044 9308 186096 9314
rect 186044 9250 186096 9256
rect 183756 5902 184888 5930
rect 183756 480 183784 5902
rect 184848 5772 184900 5778
rect 184848 5714 184900 5720
rect 184860 480 184888 5714
rect 186056 480 186084 9250
rect 187620 3482 187648 11630
rect 191748 11620 191800 11626
rect 191748 11562 191800 11568
rect 189632 9376 189684 9382
rect 189632 9318 189684 9324
rect 188436 5704 188488 5710
rect 188436 5646 188488 5652
rect 187252 3454 187648 3482
rect 187252 480 187280 3454
rect 188448 480 188476 5646
rect 189644 480 189672 9318
rect 191760 3482 191788 11562
rect 194508 11552 194560 11558
rect 194508 11494 194560 11500
rect 193220 9444 193272 9450
rect 193220 9386 193272 9392
rect 192024 5636 192076 5642
rect 192024 5578 192076 5584
rect 190840 3454 191788 3482
rect 190840 480 190868 3454
rect 192036 480 192064 5578
rect 193232 480 193260 9386
rect 194520 3482 194548 11494
rect 198648 11484 198700 11490
rect 198648 11426 198700 11432
rect 196808 9512 196860 9518
rect 196808 9454 196860 9460
rect 195612 5568 195664 5574
rect 195612 5510 195664 5516
rect 194428 3454 194548 3482
rect 194428 480 194456 3454
rect 195624 480 195652 5510
rect 196820 480 196848 9454
rect 198660 3482 198688 11426
rect 200040 3482 200068 12990
rect 201500 11416 201552 11422
rect 201500 11358 201552 11364
rect 200396 9580 200448 9586
rect 200396 9522 200448 9528
rect 198016 3454 198688 3482
rect 199212 3454 200068 3482
rect 198016 480 198044 3454
rect 199212 480 199240 3454
rect 200408 480 200436 9522
rect 201512 480 201540 11358
rect 202800 3482 202828 13738
rect 206928 12980 206980 12986
rect 206928 12922 206980 12928
rect 205548 11348 205600 11354
rect 205548 11290 205600 11296
rect 203892 9648 203944 9654
rect 203892 9590 203944 9596
rect 202708 3454 202828 3482
rect 202708 480 202736 3454
rect 203904 480 203932 9590
rect 205560 610 205588 11290
rect 206940 610 206968 12922
rect 213828 12912 213880 12918
rect 213828 12854 213880 12860
rect 211068 12844 211120 12850
rect 211068 12786 211120 12792
rect 210976 8900 211028 8906
rect 210976 8842 211028 8848
rect 207480 8832 207532 8838
rect 207480 8774 207532 8780
rect 205088 604 205140 610
rect 205088 546 205140 552
rect 205548 604 205600 610
rect 205548 546 205600 552
rect 206284 604 206336 610
rect 206284 546 206336 552
rect 206928 604 206980 610
rect 206928 546 206980 552
rect 205100 480 205128 546
rect 206296 480 206324 546
rect 207492 480 207520 8774
rect 208676 4548 208728 4554
rect 208676 4490 208728 4496
rect 208688 480 208716 4490
rect 209872 4208 209924 4214
rect 209872 4150 209924 4156
rect 209884 480 209912 4150
rect 210988 3482 211016 8842
rect 211080 4214 211108 12786
rect 212264 4480 212316 4486
rect 212264 4422 212316 4428
rect 211068 4208 211120 4214
rect 211068 4150 211120 4156
rect 210988 3454 211108 3482
rect 211080 480 211108 3454
rect 212276 480 212304 4422
rect 213840 3482 213868 12854
rect 217968 12776 218020 12782
rect 217968 12718 218020 12724
rect 214656 8764 214708 8770
rect 214656 8706 214708 8712
rect 213472 3454 213868 3482
rect 213472 480 213500 3454
rect 214668 480 214696 8706
rect 215852 4752 215904 4758
rect 215852 4694 215904 4700
rect 215864 480 215892 4694
rect 217980 3482 218008 12718
rect 220728 12708 220780 12714
rect 220728 12650 220780 12656
rect 218152 8628 218204 8634
rect 218152 8570 218204 8576
rect 217060 3454 218008 3482
rect 217060 480 217088 3454
rect 218164 480 218192 8570
rect 219346 4856 219402 4865
rect 219346 4791 219402 4800
rect 219360 480 219388 4791
rect 220740 610 220768 12650
rect 221740 8696 221792 8702
rect 221740 8638 221792 8644
rect 220544 604 220596 610
rect 220544 546 220596 552
rect 220728 604 220780 610
rect 220728 546 220780 552
rect 220556 480 220584 546
rect 221752 480 221780 8638
rect 225328 8560 225380 8566
rect 225328 8502 225380 8508
rect 224132 7200 224184 7206
rect 224132 7142 224184 7148
rect 222936 4684 222988 4690
rect 222936 4626 222988 4632
rect 222948 480 222976 4626
rect 224144 480 224172 7142
rect 225340 480 225368 8502
rect 228916 8492 228968 8498
rect 228916 8434 228968 8440
rect 227720 7132 227772 7138
rect 227720 7074 227772 7080
rect 226524 4616 226576 4622
rect 226524 4558 226576 4564
rect 226536 480 226564 4558
rect 227732 480 227760 7074
rect 228928 480 228956 8434
rect 229112 4826 229140 340054
rect 230492 4894 230520 340054
rect 230664 335640 230716 335646
rect 230664 335582 230716 335588
rect 230676 7614 230704 335582
rect 230664 7608 230716 7614
rect 230664 7550 230716 7556
rect 230768 4962 230796 340054
rect 231504 335646 231532 340054
rect 232424 337385 232452 340068
rect 232608 340054 233082 340082
rect 233252 340054 233634 340082
rect 233804 340054 234278 340082
rect 232410 337376 232466 337385
rect 232410 337311 232466 337320
rect 231492 335640 231544 335646
rect 231492 335582 231544 335588
rect 232608 333282 232636 340054
rect 232240 333254 232636 333282
rect 232240 328438 232268 333254
rect 232228 328432 232280 328438
rect 232228 328374 232280 328380
rect 232320 328432 232372 328438
rect 232320 328374 232372 328380
rect 232332 324290 232360 328374
rect 232320 324284 232372 324290
rect 232320 324226 232372 324232
rect 232424 314702 232452 314733
rect 232412 314696 232464 314702
rect 232332 314644 232412 314650
rect 232332 314638 232464 314644
rect 232332 314622 232452 314638
rect 232332 313274 232360 314622
rect 232320 313268 232372 313274
rect 232320 313210 232372 313216
rect 232320 294908 232372 294914
rect 232320 294850 232372 294856
rect 232332 293962 232360 294850
rect 232320 293956 232372 293962
rect 232320 293898 232372 293904
rect 232412 293956 232464 293962
rect 232412 293898 232464 293904
rect 232424 292534 232452 293898
rect 232412 292528 232464 292534
rect 232412 292470 232464 292476
rect 232412 282940 232464 282946
rect 232412 282882 232464 282888
rect 232424 273358 232452 282882
rect 232136 273352 232188 273358
rect 232136 273294 232188 273300
rect 232412 273352 232464 273358
rect 232412 273294 232464 273300
rect 232148 271862 232176 273294
rect 232136 271856 232188 271862
rect 232136 271798 232188 271804
rect 232320 262268 232372 262274
rect 232320 262210 232372 262216
rect 232332 253978 232360 262210
rect 232136 253972 232188 253978
rect 232136 253914 232188 253920
rect 232320 253972 232372 253978
rect 232320 253914 232372 253920
rect 232148 244254 232176 253914
rect 231952 244248 232004 244254
rect 231952 244190 232004 244196
rect 232136 244248 232188 244254
rect 232136 244190 232188 244196
rect 231964 226386 231992 244190
rect 231872 226358 231992 226386
rect 231872 225026 231900 226358
rect 231872 224998 232176 225026
rect 232148 224890 232176 224998
rect 232056 224862 232176 224890
rect 232056 216646 232084 224862
rect 231860 216640 231912 216646
rect 231860 216582 231912 216588
rect 232044 216640 232096 216646
rect 232044 216582 232096 216588
rect 231872 205578 231900 216582
rect 231872 205550 231992 205578
rect 231964 196058 231992 205550
rect 231964 196030 232084 196058
rect 232056 191826 232084 196030
rect 231952 191820 232004 191826
rect 231952 191762 232004 191768
rect 232044 191820 232096 191826
rect 232044 191762 232096 191768
rect 231964 186266 231992 191762
rect 231964 186238 232084 186266
rect 232056 182186 232084 186238
rect 232056 182170 232176 182186
rect 231952 182164 232004 182170
rect 232056 182164 232188 182170
rect 232056 182158 232136 182164
rect 231952 182106 232004 182112
rect 232136 182106 232188 182112
rect 231964 164286 231992 182106
rect 231952 164280 232004 164286
rect 231952 164222 232004 164228
rect 232044 164280 232096 164286
rect 232044 164222 232096 164228
rect 232056 157418 232084 164222
rect 232044 157412 232096 157418
rect 232044 157354 232096 157360
rect 232136 157344 232188 157350
rect 232136 157286 232188 157292
rect 232148 147642 232176 157286
rect 231964 147614 232176 147642
rect 231964 137986 231992 147614
rect 231872 137958 231992 137986
rect 231872 128330 231900 137958
rect 231872 128302 232084 128330
rect 232056 118726 232084 128302
rect 231860 118720 231912 118726
rect 231860 118662 231912 118668
rect 232044 118720 232096 118726
rect 232044 118662 232096 118668
rect 231872 109018 231900 118662
rect 231872 108990 232084 109018
rect 232056 101454 232084 108990
rect 231860 101448 231912 101454
rect 231860 101390 231912 101396
rect 232044 101448 232096 101454
rect 232044 101390 232096 101396
rect 231872 89706 231900 101390
rect 231872 89678 232084 89706
rect 232056 77314 232084 89678
rect 232044 77308 232096 77314
rect 232044 77250 232096 77256
rect 232044 77172 232096 77178
rect 232044 77114 232096 77120
rect 232056 67590 232084 77114
rect 231860 67584 231912 67590
rect 231860 67526 231912 67532
rect 232044 67584 232096 67590
rect 232044 67526 232096 67532
rect 231872 61418 231900 67526
rect 231872 61390 232176 61418
rect 232148 57882 232176 61390
rect 232056 57854 232176 57882
rect 232056 52986 232084 57854
rect 231964 52958 232084 52986
rect 231964 46918 231992 52958
rect 231952 46912 232004 46918
rect 231952 46854 232004 46860
rect 232044 37324 232096 37330
rect 232044 37266 232096 37272
rect 232056 35902 232084 37266
rect 232044 35896 232096 35902
rect 232044 35838 232096 35844
rect 231860 26308 231912 26314
rect 231860 26250 231912 26256
rect 231872 26178 231900 26250
rect 231768 26172 231820 26178
rect 231768 26114 231820 26120
rect 231860 26172 231912 26178
rect 231860 26114 231912 26120
rect 231780 21434 231808 26114
rect 231780 21406 231900 21434
rect 231308 7608 231360 7614
rect 231308 7550 231360 7556
rect 230756 4956 230808 4962
rect 230756 4898 230808 4904
rect 230480 4888 230532 4894
rect 230480 4830 230532 4836
rect 229100 4820 229152 4826
rect 229100 4762 229152 4768
rect 230112 4820 230164 4826
rect 230112 4762 230164 4768
rect 230124 480 230152 4762
rect 231320 480 231348 7550
rect 231872 3369 231900 21406
rect 232504 8424 232556 8430
rect 232504 8366 232556 8372
rect 231858 3360 231914 3369
rect 231858 3295 231914 3304
rect 232516 480 232544 8366
rect 233252 5030 233280 340054
rect 233804 335594 233832 340054
rect 234908 337550 234936 340068
rect 234896 337544 234948 337550
rect 234896 337486 234948 337492
rect 235460 337414 235488 340068
rect 235448 337408 235500 337414
rect 235448 337350 235500 337356
rect 234342 336560 234398 336569
rect 234342 336495 234398 336504
rect 233528 335566 233832 335594
rect 233528 318850 233556 335566
rect 234356 327185 234384 336495
rect 234342 327176 234398 327185
rect 234342 327111 234398 327120
rect 233424 318844 233476 318850
rect 233424 318786 233476 318792
rect 233516 318844 233568 318850
rect 233516 318786 233568 318792
rect 233436 318730 233464 318786
rect 233436 318702 233556 318730
rect 233528 302258 233556 318702
rect 234250 303104 234306 303113
rect 234250 303039 234306 303048
rect 233332 302252 233384 302258
rect 233332 302194 233384 302200
rect 233516 302252 233568 302258
rect 233516 302194 233568 302200
rect 233344 302138 233372 302194
rect 233344 302110 233464 302138
rect 233436 292618 233464 302110
rect 234264 299713 234292 303039
rect 234250 299704 234306 299713
rect 234250 299639 234306 299648
rect 233436 292590 233556 292618
rect 233528 282946 233556 292590
rect 233332 282940 233384 282946
rect 233332 282882 233384 282888
rect 233516 282940 233568 282946
rect 233516 282882 233568 282888
rect 233344 282826 233372 282882
rect 233344 282798 233464 282826
rect 233436 273306 233464 282798
rect 233436 273278 233556 273306
rect 233528 263634 233556 273278
rect 233332 263628 233384 263634
rect 233332 263570 233384 263576
rect 233516 263628 233568 263634
rect 233516 263570 233568 263576
rect 233344 263514 233372 263570
rect 236000 263560 236052 263566
rect 233344 263486 233464 263514
rect 236000 263502 236052 263508
rect 233436 253994 233464 263486
rect 233974 262032 234030 262041
rect 233974 261967 234030 261976
rect 233436 253966 233556 253994
rect 233528 244322 233556 253966
rect 233988 252657 234016 261967
rect 236012 254017 236040 263502
rect 235998 254008 236054 254017
rect 235998 253943 236054 253952
rect 233974 252648 234030 252657
rect 233974 252583 234030 252592
rect 233332 244316 233384 244322
rect 233332 244258 233384 244264
rect 233516 244316 233568 244322
rect 233516 244258 233568 244264
rect 233344 244202 233372 244258
rect 233344 244174 233464 244202
rect 233436 234682 233464 244174
rect 233436 234654 233556 234682
rect 233528 225010 233556 234654
rect 233332 225004 233384 225010
rect 233332 224946 233384 224952
rect 233516 225004 233568 225010
rect 233516 224946 233568 224952
rect 233344 224890 233372 224946
rect 233344 224862 233464 224890
rect 233436 215370 233464 224862
rect 233436 215342 233556 215370
rect 233528 205698 233556 215342
rect 234342 206952 234398 206961
rect 234342 206887 234398 206896
rect 233332 205692 233384 205698
rect 233332 205634 233384 205640
rect 233516 205692 233568 205698
rect 233516 205634 233568 205640
rect 233344 205578 233372 205634
rect 233344 205550 233464 205578
rect 233436 196058 233464 205550
rect 234356 197577 234384 206887
rect 234342 197568 234398 197577
rect 234342 197503 234398 197512
rect 233436 196030 233556 196058
rect 233528 186386 233556 196030
rect 234526 187504 234582 187513
rect 234526 187439 234582 187448
rect 233332 186380 233384 186386
rect 233332 186322 233384 186328
rect 233516 186380 233568 186386
rect 233516 186322 233568 186328
rect 233344 176610 233372 186322
rect 234540 178129 234568 187439
rect 234526 178120 234582 178129
rect 234526 178055 234582 178064
rect 233344 176582 233556 176610
rect 233528 167074 233556 176582
rect 233332 167068 233384 167074
rect 233332 167010 233384 167016
rect 233516 167068 233568 167074
rect 233516 167010 233568 167016
rect 233344 157298 233372 167010
rect 233344 157270 233556 157298
rect 233528 147694 233556 157270
rect 233332 147688 233384 147694
rect 233332 147630 233384 147636
rect 233516 147688 233568 147694
rect 233516 147630 233568 147636
rect 233344 137986 233372 147630
rect 234342 138680 234398 138689
rect 234342 138615 234398 138624
rect 233344 137958 233556 137986
rect 233528 128382 233556 137958
rect 233332 128376 233384 128382
rect 233332 128318 233384 128324
rect 233516 128376 233568 128382
rect 233516 128318 233568 128324
rect 233344 118674 233372 128318
rect 234356 121825 234384 138615
rect 234342 121816 234398 121825
rect 234342 121751 234398 121760
rect 234710 121408 234766 121417
rect 234710 121343 234766 121352
rect 233344 118646 233556 118674
rect 233528 109070 233556 118646
rect 234724 112985 234752 121343
rect 234710 112976 234766 112985
rect 234710 112911 234766 112920
rect 233332 109064 233384 109070
rect 233332 109006 233384 109012
rect 233516 109064 233568 109070
rect 233516 109006 233568 109012
rect 233344 99362 233372 109006
rect 233344 99334 233556 99362
rect 233528 89758 233556 99334
rect 233332 89752 233384 89758
rect 233332 89694 233384 89700
rect 233516 89752 233568 89758
rect 233516 89694 233568 89700
rect 233344 80050 233372 89694
rect 233344 80022 233556 80050
rect 233528 48346 233556 80022
rect 233424 48340 233476 48346
rect 233424 48282 233476 48288
rect 233516 48340 233568 48346
rect 233516 48282 233568 48288
rect 233436 41426 233464 48282
rect 233436 41398 233556 41426
rect 233528 31770 233556 41398
rect 233344 31742 233556 31770
rect 233344 31634 233372 31742
rect 233344 31606 233464 31634
rect 233436 8344 233464 31606
rect 233344 8316 233464 8344
rect 236000 8356 236052 8362
rect 233344 7682 233372 8316
rect 236000 8298 236052 8304
rect 233332 7676 233384 7682
rect 233332 7618 233384 7624
rect 234804 7676 234856 7682
rect 234804 7618 234856 7624
rect 233240 5024 233292 5030
rect 233240 4966 233292 4972
rect 233700 4888 233752 4894
rect 233700 4830 233752 4836
rect 233712 480 233740 4830
rect 234816 480 234844 7618
rect 236012 480 236040 8298
rect 236104 5098 236132 340068
rect 236196 340054 236762 340082
rect 236932 340054 237314 340082
rect 237576 340054 237958 340082
rect 238312 340054 238602 340082
rect 238864 340054 239154 340082
rect 236196 11762 236224 340054
rect 236932 328506 236960 340054
rect 237472 335640 237524 335646
rect 237472 335582 237524 335588
rect 236276 328500 236328 328506
rect 236276 328442 236328 328448
rect 236920 328500 236972 328506
rect 236920 328442 236972 328448
rect 236288 318850 236316 328442
rect 236276 318844 236328 318850
rect 236276 318786 236328 318792
rect 236368 318844 236420 318850
rect 236368 318786 236420 318792
rect 236380 304978 236408 318786
rect 236368 304972 236420 304978
rect 236368 304914 236420 304920
rect 236552 304972 236604 304978
rect 236552 304914 236604 304920
rect 236564 295361 236592 304914
rect 236274 295352 236330 295361
rect 236550 295352 236606 295361
rect 236274 295287 236276 295296
rect 236328 295287 236330 295296
rect 236460 295316 236512 295322
rect 236276 295258 236328 295264
rect 236550 295287 236606 295296
rect 236460 295258 236512 295264
rect 236472 292534 236500 295258
rect 236460 292528 236512 292534
rect 236460 292470 236512 292476
rect 236460 284368 236512 284374
rect 236460 284310 236512 284316
rect 236472 276185 236500 284310
rect 236458 276176 236514 276185
rect 236458 276111 236514 276120
rect 236274 276040 236330 276049
rect 236274 275975 236330 275984
rect 236288 273290 236316 275975
rect 236276 273284 236328 273290
rect 236276 273226 236328 273232
rect 236274 254008 236330 254017
rect 236274 253943 236330 253952
rect 236288 253910 236316 253943
rect 236276 253904 236328 253910
rect 236276 253846 236328 253852
rect 236276 234660 236328 234666
rect 236276 234602 236328 234608
rect 236288 225146 236316 234602
rect 236276 225140 236328 225146
rect 236276 225082 236328 225088
rect 236276 225004 236328 225010
rect 236276 224946 236328 224952
rect 236288 224874 236316 224946
rect 236276 224868 236328 224874
rect 236276 224810 236328 224816
rect 236276 215348 236328 215354
rect 236276 215290 236328 215296
rect 236288 215234 236316 215290
rect 236288 215206 236408 215234
rect 236380 207058 236408 215206
rect 236368 207052 236420 207058
rect 236368 206994 236420 207000
rect 236644 206916 236696 206922
rect 236644 206858 236696 206864
rect 236656 198626 236684 206858
rect 236460 198620 236512 198626
rect 236460 198562 236512 198568
rect 236644 198620 236696 198626
rect 236644 198562 236696 198568
rect 236472 187746 236500 198562
rect 236276 187740 236328 187746
rect 236276 187682 236328 187688
rect 236460 187740 236512 187746
rect 236460 187682 236512 187688
rect 236288 187610 236316 187682
rect 236276 187604 236328 187610
rect 236276 187546 236328 187552
rect 236460 178084 236512 178090
rect 236460 178026 236512 178032
rect 236472 163033 236500 178026
rect 236458 163024 236514 163033
rect 236458 162959 236514 162968
rect 236274 162888 236330 162897
rect 236330 162846 236408 162874
rect 236274 162823 236330 162832
rect 236380 151774 236408 162846
rect 236368 151768 236420 151774
rect 236368 151710 236420 151716
rect 236368 143472 236420 143478
rect 236368 143414 236420 143420
rect 236380 134065 236408 143414
rect 236366 134056 236422 134065
rect 236366 133991 236422 134000
rect 236274 133920 236330 133929
rect 236274 133855 236330 133864
rect 236288 125798 236316 133855
rect 236276 125792 236328 125798
rect 236276 125734 236328 125740
rect 236276 125656 236328 125662
rect 236276 125598 236328 125604
rect 236288 118046 236316 125598
rect 236276 118040 236328 118046
rect 236276 117982 236328 117988
rect 236460 118040 236512 118046
rect 236460 117982 236512 117988
rect 236472 113234 236500 117982
rect 236380 113206 236500 113234
rect 236380 113150 236408 113206
rect 236368 113144 236420 113150
rect 236368 113086 236420 113092
rect 236276 103556 236328 103562
rect 236276 103498 236328 103504
rect 236288 103154 236316 103498
rect 236276 103148 236328 103154
rect 236276 103090 236328 103096
rect 236460 103148 236512 103154
rect 236460 103090 236512 103096
rect 236472 96642 236500 103090
rect 236380 96614 236500 96642
rect 236380 95198 236408 96614
rect 236368 95192 236420 95198
rect 236368 95134 236420 95140
rect 236276 85604 236328 85610
rect 236276 85546 236328 85552
rect 236288 85474 236316 85546
rect 236276 85468 236328 85474
rect 236276 85410 236328 85416
rect 236368 75948 236420 75954
rect 236368 75890 236420 75896
rect 236380 67862 236408 75890
rect 236368 67856 236420 67862
rect 236368 67798 236420 67804
rect 236276 67584 236328 67590
rect 236276 67526 236328 67532
rect 236288 66178 236316 67526
rect 236288 66150 236408 66178
rect 236380 48414 236408 66150
rect 236368 48408 236420 48414
rect 236368 48350 236420 48356
rect 236276 48340 236328 48346
rect 236276 48282 236328 48288
rect 236288 46918 236316 48282
rect 236276 46912 236328 46918
rect 236276 46854 236328 46860
rect 236368 37324 236420 37330
rect 236368 37266 236420 37272
rect 236380 26246 236408 37266
rect 236368 26240 236420 26246
rect 236368 26182 236420 26188
rect 236368 16652 236420 16658
rect 236368 16594 236420 16600
rect 236184 11756 236236 11762
rect 236184 11698 236236 11704
rect 236092 5092 236144 5098
rect 236092 5034 236144 5040
rect 236380 3466 236408 16594
rect 237484 5166 237512 335582
rect 237472 5160 237524 5166
rect 237472 5102 237524 5108
rect 237196 4956 237248 4962
rect 237196 4898 237248 4904
rect 236368 3460 236420 3466
rect 236368 3402 236420 3408
rect 237208 480 237236 4898
rect 237576 3534 237604 340054
rect 238312 335646 238340 340054
rect 238300 335640 238352 335646
rect 238300 335582 238352 335588
rect 238864 13122 238892 340054
rect 239784 337414 239812 340068
rect 240428 337754 240456 340068
rect 240416 337748 240468 337754
rect 240416 337690 240468 337696
rect 239772 337408 239824 337414
rect 239772 337350 239824 337356
rect 240520 331242 240548 340190
rect 241638 340054 241744 340082
rect 241520 335640 241572 335646
rect 241520 335582 241572 335588
rect 240152 331214 240548 331242
rect 240152 331106 240180 331214
rect 240152 331078 240272 331106
rect 240244 302274 240272 331078
rect 240152 302246 240272 302274
rect 240152 302138 240180 302246
rect 240152 302110 240272 302138
rect 240244 282962 240272 302110
rect 240152 282934 240272 282962
rect 240152 282826 240180 282934
rect 240152 282798 240272 282826
rect 240244 263650 240272 282798
rect 240152 263622 240272 263650
rect 240152 263514 240180 263622
rect 240152 263486 240272 263514
rect 240244 244338 240272 263486
rect 240152 244310 240272 244338
rect 240152 244202 240180 244310
rect 240152 244174 240272 244202
rect 240244 225026 240272 244174
rect 240152 224998 240272 225026
rect 240152 224890 240180 224998
rect 240152 224862 240272 224890
rect 240244 205714 240272 224862
rect 240152 205686 240272 205714
rect 240152 205578 240180 205686
rect 240152 205550 240272 205578
rect 240244 186402 240272 205550
rect 240152 186374 240272 186402
rect 240152 186266 240180 186374
rect 240152 186238 240272 186266
rect 240244 167090 240272 186238
rect 240152 167062 240272 167090
rect 240152 166954 240180 167062
rect 240152 166926 240272 166954
rect 240244 154737 240272 166926
rect 240230 154728 240286 154737
rect 240230 154663 240286 154672
rect 240230 154592 240286 154601
rect 240230 154527 240286 154536
rect 240244 153202 240272 154527
rect 240232 153196 240284 153202
rect 240232 153138 240284 153144
rect 240508 153196 240560 153202
rect 240508 153138 240560 153144
rect 240520 143585 240548 153138
rect 240322 143576 240378 143585
rect 240322 143511 240378 143520
rect 240506 143576 240562 143585
rect 240506 143511 240562 143520
rect 240336 125662 240364 143511
rect 240140 125656 240192 125662
rect 240140 125598 240192 125604
rect 240324 125656 240376 125662
rect 240324 125598 240376 125604
rect 240152 124166 240180 125598
rect 240140 124160 240192 124166
rect 240140 124102 240192 124108
rect 240232 114572 240284 114578
rect 240232 114514 240284 114520
rect 240244 106282 240272 114514
rect 240232 106276 240284 106282
rect 240232 106218 240284 106224
rect 240140 96688 240192 96694
rect 240140 96630 240192 96636
rect 240152 95198 240180 96630
rect 240140 95192 240192 95198
rect 240140 95134 240192 95140
rect 240232 85672 240284 85678
rect 240232 85614 240284 85620
rect 240244 85524 240272 85614
rect 240244 85496 240456 85524
rect 240428 75954 240456 85496
rect 240232 75948 240284 75954
rect 240232 75890 240284 75896
rect 240416 75948 240468 75954
rect 240416 75890 240468 75896
rect 240244 72570 240272 75890
rect 240244 72542 240364 72570
rect 240336 67658 240364 72542
rect 240140 67652 240192 67658
rect 240140 67594 240192 67600
rect 240324 67652 240376 67658
rect 240324 67594 240376 67600
rect 240046 64968 240102 64977
rect 240046 64903 240102 64912
rect 240060 64530 240088 64903
rect 240048 64524 240100 64530
rect 240048 64466 240100 64472
rect 240152 58002 240180 67594
rect 240140 57996 240192 58002
rect 240140 57938 240192 57944
rect 240232 57996 240284 58002
rect 240232 57938 240284 57944
rect 240244 56574 240272 57938
rect 240232 56568 240284 56574
rect 240232 56510 240284 56516
rect 240232 46980 240284 46986
rect 240232 46922 240284 46928
rect 240046 43888 240102 43897
rect 240046 43823 240102 43832
rect 240060 40225 240088 43823
rect 240046 40216 240102 40225
rect 240046 40151 240102 40160
rect 240244 31890 240272 46922
rect 240232 31884 240284 31890
rect 240232 31826 240284 31832
rect 240232 26376 240284 26382
rect 240232 26318 240284 26324
rect 240244 26246 240272 26318
rect 240232 26240 240284 26246
rect 240232 26182 240284 26188
rect 240324 26172 240376 26178
rect 240324 26114 240376 26120
rect 240138 16824 240194 16833
rect 240138 16759 240194 16768
rect 240152 16674 240180 16759
rect 240230 16688 240286 16697
rect 240152 16646 240230 16674
rect 240230 16623 240286 16632
rect 240048 14068 240100 14074
rect 240048 14010 240100 14016
rect 238852 13116 238904 13122
rect 238852 13058 238904 13064
rect 238392 7064 238444 7070
rect 238392 7006 238444 7012
rect 237564 3528 237616 3534
rect 237564 3470 237616 3476
rect 238404 480 238432 7006
rect 240060 3670 240088 14010
rect 240336 12322 240364 26114
rect 240244 12294 240364 12322
rect 240244 5234 240272 12294
rect 240232 5228 240284 5234
rect 240232 5170 240284 5176
rect 240784 5024 240836 5030
rect 240784 4966 240836 4972
rect 239588 3664 239640 3670
rect 239588 3606 239640 3612
rect 240048 3664 240100 3670
rect 240048 3606 240100 3612
rect 239600 480 239628 3606
rect 240796 480 240824 4966
rect 241532 3602 241560 335582
rect 241716 14482 241744 340054
rect 241992 340054 242282 340082
rect 241992 335646 242020 340054
rect 241980 335640 242032 335646
rect 241980 335582 242032 335588
rect 242360 328506 242388 340190
rect 242912 340054 243478 340082
rect 243832 340054 244122 340082
rect 241796 328500 241848 328506
rect 241796 328442 241848 328448
rect 242348 328500 242400 328506
rect 242348 328442 242400 328448
rect 241808 299470 241836 328442
rect 241796 299464 241848 299470
rect 241796 299406 241848 299412
rect 241796 289876 241848 289882
rect 241796 289818 241848 289824
rect 241808 280158 241836 289818
rect 241796 280152 241848 280158
rect 241796 280094 241848 280100
rect 241796 270564 241848 270570
rect 241796 270506 241848 270512
rect 241808 260846 241836 270506
rect 241796 260840 241848 260846
rect 241796 260782 241848 260788
rect 241796 251252 241848 251258
rect 241796 251194 241848 251200
rect 241808 183569 241836 251194
rect 242714 240136 242770 240145
rect 242714 240071 242770 240080
rect 242728 230518 242756 240071
rect 242716 230512 242768 230518
rect 242716 230454 242768 230460
rect 242808 230512 242860 230518
rect 242808 230454 242860 230460
rect 242820 222222 242848 230454
rect 242808 222216 242860 222222
rect 242808 222158 242860 222164
rect 241794 183560 241850 183569
rect 241794 183495 241850 183504
rect 241978 183560 242034 183569
rect 241978 183495 242034 183504
rect 241992 173942 242020 183495
rect 241796 173936 241848 173942
rect 241796 173878 241848 173884
rect 241980 173936 242032 173942
rect 241980 173878 242032 173884
rect 241808 106282 241836 173878
rect 241796 106276 241848 106282
rect 241796 106218 241848 106224
rect 241980 106276 242032 106282
rect 241980 106218 242032 106224
rect 241992 96665 242020 106218
rect 241794 96656 241850 96665
rect 241794 96591 241850 96600
rect 241978 96656 242034 96665
rect 241978 96591 242034 96600
rect 241808 86970 241836 96591
rect 241796 86964 241848 86970
rect 241796 86906 241848 86912
rect 241796 77308 241848 77314
rect 241796 77250 241848 77256
rect 241704 14476 241756 14482
rect 241704 14418 241756 14424
rect 241520 3596 241572 3602
rect 241520 3538 241572 3544
rect 241808 3534 241836 77250
rect 242912 7750 242940 340054
rect 243832 335646 243860 340054
rect 244660 337550 244688 340068
rect 244844 340054 245318 340082
rect 245764 340054 245962 340082
rect 246224 340054 246514 340082
rect 247158 340054 247264 340082
rect 244648 337544 244700 337550
rect 244648 337486 244700 337492
rect 244844 335730 244872 340054
rect 244476 335702 244872 335730
rect 243084 335640 243136 335646
rect 243084 335582 243136 335588
rect 243820 335640 243872 335646
rect 243820 335582 243872 335588
rect 243096 307766 243124 335582
rect 244476 311930 244504 335702
rect 245660 335640 245712 335646
rect 245660 335582 245712 335588
rect 244384 311902 244504 311930
rect 244384 311794 244412 311902
rect 244384 311766 244504 311794
rect 243084 307760 243136 307766
rect 243084 307702 243136 307708
rect 242992 298240 243044 298246
rect 242992 298182 243044 298188
rect 243004 298110 243032 298182
rect 242992 298104 243044 298110
rect 242992 298046 243044 298052
rect 244476 292534 244504 311766
rect 244464 292528 244516 292534
rect 244464 292470 244516 292476
rect 244464 292392 244516 292398
rect 244464 292334 244516 292340
rect 243176 280220 243228 280226
rect 243176 280162 243228 280168
rect 243188 280129 243216 280162
rect 243174 280120 243230 280129
rect 243174 280055 243230 280064
rect 243358 280120 243414 280129
rect 243358 280055 243414 280064
rect 243372 270745 243400 280055
rect 244476 273222 244504 292334
rect 244464 273216 244516 273222
rect 244464 273158 244516 273164
rect 244464 273080 244516 273086
rect 244464 273022 244516 273028
rect 243358 270736 243414 270745
rect 243358 270671 243414 270680
rect 243082 270600 243138 270609
rect 243082 270535 243138 270544
rect 243096 270502 243124 270535
rect 243084 270496 243136 270502
rect 243084 270438 243136 270444
rect 243176 260908 243228 260914
rect 243176 260850 243228 260856
rect 243188 260817 243216 260850
rect 243174 260808 243230 260817
rect 243174 260743 243230 260752
rect 243358 260808 243414 260817
rect 243358 260743 243414 260752
rect 243372 251433 243400 260743
rect 244476 253910 244504 273022
rect 244464 253904 244516 253910
rect 244464 253846 244516 253852
rect 244464 253768 244516 253774
rect 244464 253710 244516 253716
rect 243358 251424 243414 251433
rect 243358 251359 243414 251368
rect 243082 251288 243138 251297
rect 243082 251223 243138 251232
rect 243096 244322 243124 251223
rect 243084 244316 243136 244322
rect 243084 244258 243136 244264
rect 243176 244180 243228 244186
rect 243176 244122 243228 244128
rect 243188 241482 243216 244122
rect 243004 241454 243216 241482
rect 243004 240145 243032 241454
rect 242990 240136 243046 240145
rect 242990 240071 243046 240080
rect 243188 222222 243216 222253
rect 243176 222216 243228 222222
rect 243096 222164 243176 222170
rect 243096 222158 243228 222164
rect 243096 222142 243216 222158
rect 243096 222086 243124 222142
rect 243084 222080 243136 222086
rect 243084 222022 243136 222028
rect 243176 212560 243228 212566
rect 243176 212502 243228 212508
rect 243188 205698 243216 212502
rect 243176 205692 243228 205698
rect 243176 205634 243228 205640
rect 243188 202910 243216 202941
rect 243176 202904 243228 202910
rect 243096 202852 243176 202858
rect 243096 202846 243228 202852
rect 243096 202830 243216 202846
rect 243096 202774 243124 202830
rect 243084 202768 243136 202774
rect 243084 202710 243136 202716
rect 243176 193248 243228 193254
rect 243176 193190 243228 193196
rect 243188 186386 243216 193190
rect 243176 186380 243228 186386
rect 243176 186322 243228 186328
rect 243084 186312 243136 186318
rect 243084 186254 243136 186260
rect 243096 183705 243124 186254
rect 243082 183696 243138 183705
rect 243082 183631 243138 183640
rect 243266 183560 243322 183569
rect 243266 183495 243322 183504
rect 243280 173942 243308 183495
rect 244476 176662 244504 253710
rect 244464 176656 244516 176662
rect 244464 176598 244516 176604
rect 244464 176520 244516 176526
rect 244464 176462 244516 176468
rect 243176 173936 243228 173942
rect 243176 173878 243228 173884
rect 243268 173936 243320 173942
rect 243268 173878 243320 173884
rect 243188 167142 243216 173878
rect 243176 167136 243228 167142
rect 243176 167078 243228 167084
rect 242992 162920 243044 162926
rect 242992 162862 243044 162868
rect 243004 154562 243032 162862
rect 242992 154556 243044 154562
rect 242992 154498 243044 154504
rect 243084 147620 243136 147626
rect 243084 147562 243136 147568
rect 243096 144922 243124 147562
rect 243096 144906 243216 144922
rect 243096 144900 243228 144906
rect 243096 144894 243176 144900
rect 243176 144842 243228 144848
rect 243268 144900 243320 144906
rect 243268 144842 243320 144848
rect 243280 135289 243308 144842
rect 244476 135425 244504 176462
rect 244462 135416 244518 135425
rect 244462 135351 244518 135360
rect 243082 135280 243138 135289
rect 243082 135215 243084 135224
rect 243136 135215 243138 135224
rect 243266 135280 243322 135289
rect 243266 135215 243268 135224
rect 243084 135186 243136 135192
rect 243320 135215 243322 135224
rect 243268 135186 243320 135192
rect 243280 133890 243308 135186
rect 244462 135144 244518 135153
rect 244462 135079 244518 135088
rect 243268 133884 243320 133890
rect 243268 133826 243320 133832
rect 243360 124228 243412 124234
rect 243360 124170 243412 124176
rect 243372 114578 243400 124170
rect 244476 124148 244504 135079
rect 244384 124120 244504 124148
rect 244384 118726 244412 124120
rect 244372 118720 244424 118726
rect 244372 118662 244424 118668
rect 244464 118652 244516 118658
rect 244464 118594 244516 118600
rect 243176 114572 243228 114578
rect 243096 114532 243176 114560
rect 243096 109750 243124 114532
rect 243176 114514 243228 114520
rect 243360 114572 243412 114578
rect 243360 114514 243412 114520
rect 243084 109744 243136 109750
rect 243084 109686 243136 109692
rect 243268 106208 243320 106214
rect 243268 106150 243320 106156
rect 243280 99362 243308 106150
rect 244476 99482 244504 118594
rect 244464 99476 244516 99482
rect 244464 99418 244516 99424
rect 243004 99334 243308 99362
rect 244464 99340 244516 99346
rect 243004 91798 243032 99334
rect 244464 99282 244516 99288
rect 242992 91792 243044 91798
rect 242992 91734 243044 91740
rect 243452 91792 243504 91798
rect 243452 91734 243504 91740
rect 243464 86986 243492 91734
rect 243372 86958 243492 86986
rect 243372 80782 243400 86958
rect 243360 80776 243412 80782
rect 243360 80718 243412 80724
rect 244476 70514 244504 99282
rect 244464 70508 244516 70514
rect 244464 70450 244516 70456
rect 243176 67652 243228 67658
rect 243176 67594 243228 67600
rect 244464 67652 244516 67658
rect 244464 67594 244516 67600
rect 243188 41426 243216 67594
rect 244476 62914 244504 67594
rect 244476 62886 244596 62914
rect 244568 58002 244596 62886
rect 244372 57996 244424 58002
rect 244372 57938 244424 57944
rect 244556 57996 244608 58002
rect 244556 57938 244608 57944
rect 244384 50946 244412 57938
rect 244384 50918 244504 50946
rect 244476 46918 244504 50918
rect 244464 46912 244516 46918
rect 244464 46854 244516 46860
rect 243096 41398 243216 41426
rect 243096 33810 243124 41398
rect 244556 37324 244608 37330
rect 244556 37266 244608 37272
rect 243004 33782 243124 33810
rect 243004 31634 243032 33782
rect 243004 31606 243216 31634
rect 243188 28966 243216 31606
rect 244568 29034 244596 37266
rect 244372 29028 244424 29034
rect 244372 28970 244424 28976
rect 244556 29028 244608 29034
rect 244556 28970 244608 28976
rect 243084 28960 243136 28966
rect 243084 28902 243136 28908
rect 243176 28960 243228 28966
rect 243176 28902 243228 28908
rect 243096 15910 243124 28902
rect 244384 19446 244412 28970
rect 244372 19440 244424 19446
rect 244372 19382 244424 19388
rect 244280 16652 244332 16658
rect 244280 16594 244332 16600
rect 243084 15904 243136 15910
rect 243084 15846 243136 15852
rect 244188 14476 244240 14482
rect 244188 14418 244240 14424
rect 242900 7744 242952 7750
rect 242900 7686 242952 7692
rect 241980 6996 242032 7002
rect 241980 6938 242032 6944
rect 241796 3528 241848 3534
rect 241796 3470 241848 3476
rect 241992 480 242020 6938
rect 244200 3670 244228 14418
rect 244292 7818 244320 16594
rect 244280 7812 244332 7818
rect 244280 7754 244332 7760
rect 245568 7744 245620 7750
rect 245568 7686 245620 7692
rect 244372 5092 244424 5098
rect 244372 5034 244424 5040
rect 243176 3664 243228 3670
rect 243176 3606 243228 3612
rect 244188 3664 244240 3670
rect 244188 3606 244240 3612
rect 243188 480 243216 3606
rect 244384 480 244412 5034
rect 245580 480 245608 7686
rect 245672 3738 245700 335582
rect 245764 15978 245792 340054
rect 246224 335646 246252 340054
rect 246304 337544 246356 337550
rect 246304 337486 246356 337492
rect 246212 335640 246264 335646
rect 246212 335582 246264 335588
rect 245752 15972 245804 15978
rect 245752 15914 245804 15920
rect 246316 14142 246344 337486
rect 246304 14136 246356 14142
rect 246304 14078 246356 14084
rect 246764 9920 246816 9926
rect 246764 9862 246816 9868
rect 245660 3732 245712 3738
rect 245660 3674 245712 3680
rect 246776 480 246804 9862
rect 247236 7886 247264 340054
rect 247696 337822 247724 340068
rect 247684 337816 247736 337822
rect 247684 337758 247736 337764
rect 248340 337618 248368 340068
rect 248524 340054 248998 340082
rect 249168 340054 249550 340082
rect 249812 340054 250194 340082
rect 250364 340054 250838 340082
rect 248328 337612 248380 337618
rect 248328 337554 248380 337560
rect 248420 335640 248472 335646
rect 248420 335582 248472 335588
rect 248328 64524 248380 64530
rect 248328 64466 248380 64472
rect 248340 63617 248368 64466
rect 248326 63608 248382 63617
rect 248326 63543 248382 63552
rect 247224 7880 247276 7886
rect 247224 7822 247276 7828
rect 247960 5160 248012 5166
rect 247960 5102 248012 5108
rect 247972 480 248000 5102
rect 248432 3874 248460 335582
rect 248524 7954 248552 340054
rect 249168 335646 249196 340054
rect 249156 335640 249208 335646
rect 249156 335582 249208 335588
rect 248512 7948 248564 7954
rect 248512 7890 248564 7896
rect 249156 7812 249208 7818
rect 249156 7754 249208 7760
rect 248420 3868 248472 3874
rect 248420 3810 248472 3816
rect 249168 480 249196 7754
rect 249812 3806 249840 340054
rect 250364 335730 250392 340054
rect 251376 337890 251404 340068
rect 251744 340054 252034 340082
rect 251364 337884 251416 337890
rect 251364 337826 251416 337832
rect 251744 337346 251772 340054
rect 251732 337340 251784 337346
rect 251732 337282 251784 337288
rect 251824 337340 251876 337346
rect 251824 337282 251876 337288
rect 249996 335702 250392 335730
rect 249996 321706 250024 335702
rect 249984 321700 250036 321706
rect 249984 321642 250036 321648
rect 249984 317484 250036 317490
rect 249984 317426 250036 317432
rect 249996 317370 250024 317426
rect 249996 317342 250116 317370
rect 250088 312594 250116 317342
rect 249892 312588 249944 312594
rect 249892 312530 249944 312536
rect 250076 312588 250128 312594
rect 250076 312530 250128 312536
rect 249904 304314 249932 312530
rect 249904 304286 250024 304314
rect 249996 299470 250024 304286
rect 249984 299464 250036 299470
rect 249984 299406 250036 299412
rect 249984 289876 250036 289882
rect 249984 289818 250036 289824
rect 249996 273086 250024 289818
rect 249984 273080 250036 273086
rect 249984 273022 250036 273028
rect 249984 272944 250036 272950
rect 249984 272886 250036 272892
rect 249996 253774 250024 272886
rect 249984 253768 250036 253774
rect 249984 253710 250036 253716
rect 249984 253632 250036 253638
rect 249984 253574 250036 253580
rect 249996 176526 250024 253574
rect 249984 176520 250036 176526
rect 249984 176462 250036 176468
rect 249984 176384 250036 176390
rect 249984 176326 250036 176332
rect 249996 157298 250024 176326
rect 249904 157270 250024 157298
rect 249904 157026 249932 157270
rect 249904 156998 250024 157026
rect 249996 135402 250024 156998
rect 249904 135374 250024 135402
rect 249904 135266 249932 135374
rect 249904 135238 250024 135266
rect 249996 125905 250024 135238
rect 249982 125896 250038 125905
rect 249982 125831 250038 125840
rect 249982 125624 250038 125633
rect 249982 125559 250038 125568
rect 249996 124166 250024 125559
rect 249984 124160 250036 124166
rect 249984 124102 250036 124108
rect 249984 114572 250036 114578
rect 249984 114514 250036 114520
rect 249996 85542 250024 114514
rect 249984 85536 250036 85542
rect 249984 85478 250036 85484
rect 249984 79348 250036 79354
rect 249984 79290 250036 79296
rect 249996 66230 250024 79290
rect 249892 66224 249944 66230
rect 249892 66166 249944 66172
rect 249984 66224 250036 66230
rect 249984 66166 250036 66172
rect 249904 64870 249932 66166
rect 249892 64864 249944 64870
rect 249892 64806 249944 64812
rect 249892 56568 249944 56574
rect 249892 56510 249944 56516
rect 249904 51202 249932 56510
rect 249892 51196 249944 51202
rect 249892 51138 249944 51144
rect 249892 47048 249944 47054
rect 249892 46990 249944 46996
rect 249904 46918 249932 46990
rect 249892 46912 249944 46918
rect 249892 46854 249944 46860
rect 249892 37324 249944 37330
rect 249892 37266 249944 37272
rect 249904 29034 249932 37266
rect 249892 29028 249944 29034
rect 249892 28970 249944 28976
rect 249984 29028 250036 29034
rect 249984 28970 250036 28976
rect 249996 28914 250024 28970
rect 249996 28886 250116 28914
rect 250088 19360 250116 28886
rect 250088 19332 250208 19360
rect 250180 19122 250208 19332
rect 250088 19094 250208 19122
rect 250088 9722 250116 19094
rect 251086 17096 251142 17105
rect 251086 17031 251142 17040
rect 251100 16697 251128 17031
rect 251086 16688 251142 16697
rect 251086 16623 251142 16632
rect 250352 9852 250404 9858
rect 250352 9794 250404 9800
rect 249984 9716 250036 9722
rect 249984 9658 250036 9664
rect 250076 9716 250128 9722
rect 250076 9658 250128 9664
rect 249996 8022 250024 9658
rect 249984 8016 250036 8022
rect 249984 7958 250036 7964
rect 249800 3800 249852 3806
rect 249800 3742 249852 3748
rect 250364 480 250392 9794
rect 251456 5228 251508 5234
rect 251456 5170 251508 5176
rect 251468 480 251496 5170
rect 251836 3942 251864 337282
rect 252560 318844 252612 318850
rect 252560 318786 252612 318792
rect 252572 309194 252600 318786
rect 252560 309188 252612 309194
rect 252560 309130 252612 309136
rect 252560 158024 252612 158030
rect 252560 157966 252612 157972
rect 252572 153241 252600 157966
rect 252558 153232 252614 153241
rect 252558 153167 252614 153176
rect 252558 125352 252614 125361
rect 252558 125287 252614 125296
rect 252572 119406 252600 125287
rect 252560 119400 252612 119406
rect 252560 119342 252612 119348
rect 252664 8090 252692 340068
rect 253216 337346 253244 340068
rect 253308 340054 253874 340082
rect 253952 340054 254518 340082
rect 254780 340054 255070 340082
rect 253204 337340 253256 337346
rect 253204 337282 253256 337288
rect 253308 334626 253336 340054
rect 253388 337680 253440 337686
rect 253388 337622 253440 337628
rect 252744 334620 252796 334626
rect 252744 334562 252796 334568
rect 253296 334620 253348 334626
rect 253296 334562 253348 334568
rect 252756 318918 252784 334562
rect 253400 334506 253428 337622
rect 253216 334478 253428 334506
rect 252744 318912 252796 318918
rect 252744 318854 252796 318860
rect 252744 309188 252796 309194
rect 252744 309130 252796 309136
rect 252756 289814 252784 309130
rect 252744 289808 252796 289814
rect 252744 289750 252796 289756
rect 252744 280220 252796 280226
rect 252744 280162 252796 280168
rect 252756 270502 252784 280162
rect 252744 270496 252796 270502
rect 252744 270438 252796 270444
rect 252744 260908 252796 260914
rect 252744 260850 252796 260856
rect 252756 241482 252784 260850
rect 252756 241454 252876 241482
rect 252848 231962 252876 241454
rect 252756 231934 252876 231962
rect 252756 231849 252784 231934
rect 252742 231840 252798 231849
rect 252742 231775 252798 231784
rect 252926 231840 252982 231849
rect 252926 231775 252982 231784
rect 252756 222222 252784 222253
rect 252940 222222 252968 231775
rect 252744 222216 252796 222222
rect 252928 222216 252980 222222
rect 252796 222164 252876 222170
rect 252744 222158 252876 222164
rect 252928 222158 252980 222164
rect 252756 222142 252876 222158
rect 252848 212566 252876 222142
rect 252744 212560 252796 212566
rect 252742 212528 252744 212537
rect 252836 212560 252888 212566
rect 252796 212528 252798 212537
rect 252836 212502 252888 212508
rect 252926 212528 252982 212537
rect 252742 212463 252798 212472
rect 252926 212463 252982 212472
rect 252940 205578 252968 212463
rect 252848 205550 252968 205578
rect 252848 202881 252876 205550
rect 252834 202872 252890 202881
rect 252834 202807 252890 202816
rect 253018 202872 253074 202881
rect 253018 202807 253074 202816
rect 253032 193254 253060 202807
rect 252836 193248 252888 193254
rect 252834 193216 252836 193225
rect 253020 193248 253072 193254
rect 252888 193216 252890 193225
rect 252834 193151 252890 193160
rect 253018 193216 253020 193225
rect 253072 193216 253074 193225
rect 253018 193151 253074 193160
rect 253032 183598 253060 193151
rect 252836 183592 252888 183598
rect 252836 183534 252888 183540
rect 253020 183592 253072 183598
rect 253020 183534 253072 183540
rect 252848 178838 252876 183534
rect 252836 178832 252888 178838
rect 252836 178774 252888 178780
rect 252744 173936 252796 173942
rect 252744 173878 252796 173884
rect 252756 158030 252784 173878
rect 252744 158024 252796 158030
rect 252744 157966 252796 157972
rect 252834 153232 252890 153241
rect 252834 153167 252890 153176
rect 252848 144974 252876 153167
rect 252744 144968 252796 144974
rect 252744 144910 252796 144916
rect 252836 144968 252888 144974
rect 252836 144910 252888 144916
rect 252756 143546 252784 144910
rect 252744 143540 252796 143546
rect 252744 143482 252796 143488
rect 252928 143540 252980 143546
rect 252928 143482 252980 143488
rect 252940 125633 252968 143482
rect 252926 125624 252982 125633
rect 252926 125559 252982 125568
rect 252744 106344 252796 106350
rect 252744 106286 252796 106292
rect 252756 40186 252784 106286
rect 253110 76528 253166 76537
rect 253110 76463 253166 76472
rect 253124 75993 253152 76463
rect 253110 75984 253166 75993
rect 253110 75919 253166 75928
rect 253110 64288 253166 64297
rect 253110 64223 253166 64232
rect 253124 63345 253152 64223
rect 253110 63336 253166 63345
rect 253110 63271 253166 63280
rect 252744 40180 252796 40186
rect 252744 40122 252796 40128
rect 252836 31680 252888 31686
rect 252836 31622 252888 31628
rect 252848 28966 252876 31622
rect 252836 28960 252888 28966
rect 252836 28902 252888 28908
rect 252836 19372 252888 19378
rect 252836 19314 252888 19320
rect 252848 12578 252876 19314
rect 252836 12572 252888 12578
rect 252836 12514 252888 12520
rect 252744 11756 252796 11762
rect 252744 11698 252796 11704
rect 252652 8084 252704 8090
rect 252652 8026 252704 8032
rect 252652 7880 252704 7886
rect 252652 7822 252704 7828
rect 251824 3936 251876 3942
rect 251824 3878 251876 3884
rect 252664 480 252692 7822
rect 252756 4010 252784 11698
rect 253216 4078 253244 334478
rect 253848 9784 253900 9790
rect 253848 9726 253900 9732
rect 253204 4072 253256 4078
rect 253204 4014 253256 4020
rect 252744 4004 252796 4010
rect 252744 3946 252796 3952
rect 253860 480 253888 9726
rect 253952 6225 253980 340054
rect 254780 330478 254808 340054
rect 255700 337686 255728 340068
rect 255884 340054 256358 340082
rect 256804 340054 256910 340082
rect 255688 337680 255740 337686
rect 255688 337622 255740 337628
rect 255884 331242 255912 340054
rect 255964 337340 256016 337346
rect 255964 337282 256016 337288
rect 255516 331214 255912 331242
rect 254216 330472 254268 330478
rect 254216 330414 254268 330420
rect 254768 330472 254820 330478
rect 254768 330414 254820 330420
rect 254228 321722 254256 330414
rect 254228 321694 254348 321722
rect 254320 321450 254348 321694
rect 254136 321422 254348 321450
rect 254136 318730 254164 321422
rect 254136 318702 254256 318730
rect 254228 292618 254256 318702
rect 255516 317506 255544 331214
rect 255424 317478 255544 317506
rect 255424 317422 255452 317478
rect 255412 317416 255464 317422
rect 255412 317358 255464 317364
rect 255688 317348 255740 317354
rect 255688 317290 255740 317296
rect 255700 315994 255728 317290
rect 255688 315988 255740 315994
rect 255688 315930 255740 315936
rect 255504 298172 255556 298178
rect 255504 298114 255556 298120
rect 255516 292670 255544 298114
rect 254136 292590 254256 292618
rect 255504 292664 255556 292670
rect 255504 292606 255556 292612
rect 254136 289814 254164 292590
rect 255504 292528 255556 292534
rect 255504 292470 255556 292476
rect 254124 289808 254176 289814
rect 254124 289750 254176 289756
rect 254216 277432 254268 277438
rect 254216 277374 254268 277380
rect 254228 267753 254256 277374
rect 255516 273306 255544 292470
rect 255424 273278 255544 273306
rect 255424 273170 255452 273278
rect 255424 273142 255544 273170
rect 254030 267744 254086 267753
rect 254030 267679 254086 267688
rect 254214 267744 254270 267753
rect 254214 267679 254270 267688
rect 254044 258097 254072 267679
rect 254030 258088 254086 258097
rect 254030 258023 254086 258032
rect 254214 258088 254270 258097
rect 254214 258023 254270 258032
rect 254228 254046 254256 258023
rect 254216 254040 254268 254046
rect 255516 253994 255544 273142
rect 254216 253982 254268 253988
rect 255424 253966 255544 253994
rect 255424 253858 255452 253966
rect 255424 253830 255544 253858
rect 254124 248532 254176 248538
rect 254124 248474 254176 248480
rect 254136 248402 254164 248474
rect 254124 248396 254176 248402
rect 254124 248338 254176 248344
rect 254124 244248 254176 244254
rect 254124 244190 254176 244196
rect 254136 238762 254164 244190
rect 255516 241482 255544 253830
rect 255516 241454 255636 241482
rect 254136 238734 254256 238762
rect 254228 212634 254256 238734
rect 255608 234666 255636 241454
rect 255596 234660 255648 234666
rect 255596 234602 255648 234608
rect 255504 234592 255556 234598
rect 255504 234534 255556 234540
rect 255516 222170 255544 234534
rect 255516 222142 255636 222170
rect 255608 215354 255636 222142
rect 255596 215348 255648 215354
rect 255596 215290 255648 215296
rect 255504 215280 255556 215286
rect 255504 215222 255556 215228
rect 254216 212628 254268 212634
rect 254216 212570 254268 212576
rect 254124 212560 254176 212566
rect 254124 212502 254176 212508
rect 254136 207754 254164 212502
rect 255516 211138 255544 215222
rect 255320 211132 255372 211138
rect 255320 211074 255372 211080
rect 255504 211132 255556 211138
rect 255504 211074 255556 211080
rect 254136 207726 254256 207754
rect 254228 198098 254256 207726
rect 255332 201521 255360 211074
rect 255318 201512 255374 201521
rect 255594 201512 255650 201521
rect 255318 201447 255374 201456
rect 255504 201476 255556 201482
rect 255594 201447 255596 201456
rect 255504 201418 255556 201424
rect 255648 201447 255650 201456
rect 255596 201418 255648 201424
rect 255516 200122 255544 201418
rect 255504 200116 255556 200122
rect 255504 200058 255556 200064
rect 254136 198070 254256 198098
rect 254136 193225 254164 198070
rect 254122 193216 254178 193225
rect 254122 193151 254178 193160
rect 254306 193216 254362 193225
rect 254306 193151 254362 193160
rect 254320 173942 254348 193151
rect 255504 190528 255556 190534
rect 255504 190470 255556 190476
rect 255516 180810 255544 190470
rect 255504 180804 255556 180810
rect 255504 180746 255556 180752
rect 254124 173936 254176 173942
rect 254124 173878 254176 173884
rect 254308 173936 254360 173942
rect 254308 173878 254360 173884
rect 254136 172514 254164 173878
rect 254124 172508 254176 172514
rect 254124 172450 254176 172456
rect 254124 167000 254176 167006
rect 254124 166942 254176 166948
rect 255504 167000 255556 167006
rect 255504 166942 255556 166948
rect 254136 153270 254164 166942
rect 254124 153264 254176 153270
rect 254124 153206 254176 153212
rect 254400 153264 254452 153270
rect 254400 153206 254452 153212
rect 254412 153134 254440 153206
rect 254400 153128 254452 153134
rect 254400 153070 254452 153076
rect 254124 143608 254176 143614
rect 254176 143556 254256 143562
rect 254124 143550 254256 143556
rect 254136 143546 254256 143550
rect 254136 143540 254268 143546
rect 254136 143534 254216 143540
rect 254216 143482 254268 143488
rect 255516 138122 255544 166942
rect 255424 138094 255544 138122
rect 255424 137986 255452 138094
rect 255424 137958 255544 137986
rect 254216 124228 254268 124234
rect 254216 124170 254268 124176
rect 254228 115954 254256 124170
rect 254136 115938 254256 115954
rect 254124 115932 254268 115938
rect 254176 115926 254216 115932
rect 254124 115874 254176 115880
rect 254216 115874 254268 115880
rect 254136 115843 254164 115874
rect 254228 114510 254256 115874
rect 254124 114504 254176 114510
rect 254124 114446 254176 114452
rect 254216 114504 254268 114510
rect 254216 114446 254268 114452
rect 254136 104938 254164 114446
rect 254136 104910 254256 104938
rect 254228 103494 254256 104910
rect 254216 103488 254268 103494
rect 254216 103430 254268 103436
rect 255516 99498 255544 137958
rect 255424 99470 255544 99498
rect 255424 99362 255452 99470
rect 255424 99334 255544 99362
rect 254216 93900 254268 93906
rect 254216 93842 254268 93848
rect 254228 85542 254256 93842
rect 254216 85536 254268 85542
rect 254216 85478 254268 85484
rect 255516 80034 255544 99334
rect 255504 80028 255556 80034
rect 255504 79970 255556 79976
rect 255504 74588 255556 74594
rect 255504 74530 255556 74536
rect 254124 67652 254176 67658
rect 254124 67594 254176 67600
rect 254136 60874 254164 67594
rect 255516 64870 255544 74530
rect 255504 64864 255556 64870
rect 255504 64806 255556 64812
rect 254136 60846 254256 60874
rect 254228 60704 254256 60846
rect 254136 60676 254256 60704
rect 254136 53122 254164 60676
rect 255504 55276 255556 55282
rect 255504 55218 255556 55224
rect 255516 55185 255544 55218
rect 255502 55176 255558 55185
rect 255502 55111 255558 55120
rect 255778 55176 255834 55185
rect 255778 55111 255834 55120
rect 254136 53094 254256 53122
rect 254228 28966 254256 53094
rect 255792 45626 255820 55111
rect 255596 45620 255648 45626
rect 255596 45562 255648 45568
rect 255780 45620 255832 45626
rect 255780 45562 255832 45568
rect 254216 28960 254268 28966
rect 254216 28902 254268 28908
rect 254308 28960 254360 28966
rect 254308 28902 254360 28908
rect 254320 19310 254348 28902
rect 255608 19310 255636 45562
rect 254308 19304 254360 19310
rect 254308 19246 254360 19252
rect 255596 19304 255648 19310
rect 255596 19246 255648 19252
rect 254308 19168 254360 19174
rect 254308 19110 254360 19116
rect 255596 19168 255648 19174
rect 255596 19110 255648 19116
rect 254320 9722 254348 19110
rect 255608 9722 255636 19110
rect 254032 9716 254084 9722
rect 254032 9658 254084 9664
rect 254308 9716 254360 9722
rect 254308 9658 254360 9664
rect 255320 9716 255372 9722
rect 255320 9658 255372 9664
rect 255596 9716 255648 9722
rect 255596 9658 255648 9664
rect 254044 8158 254072 9658
rect 254032 8152 254084 8158
rect 254032 8094 254084 8100
rect 253938 6216 253994 6225
rect 255332 6186 255360 9658
rect 253938 6151 253994 6160
rect 255320 6180 255372 6186
rect 255320 6122 255372 6128
rect 255976 4146 256004 337282
rect 256804 8226 256832 340054
rect 257540 337958 257568 340068
rect 258198 340054 258304 340082
rect 257528 337952 257580 337958
rect 257528 337894 257580 337900
rect 257344 337408 257396 337414
rect 257344 337350 257396 337356
rect 256792 8220 256844 8226
rect 256792 8162 256844 8168
rect 256240 7948 256292 7954
rect 256240 7890 256292 7896
rect 255964 4140 256016 4146
rect 255964 4082 256016 4088
rect 255044 3868 255096 3874
rect 255044 3810 255096 3816
rect 255056 480 255084 3810
rect 256252 480 256280 7890
rect 257356 3398 257384 337350
rect 257986 87000 258042 87009
rect 257986 86935 258042 86944
rect 258000 86873 258028 86935
rect 257986 86864 258042 86873
rect 257986 86799 258042 86808
rect 257436 9716 257488 9722
rect 257436 9658 257488 9664
rect 257344 3392 257396 3398
rect 257344 3334 257396 3340
rect 257448 480 257476 9658
rect 258276 6254 258304 340054
rect 258368 340054 258750 340082
rect 258368 8294 258396 340054
rect 258724 337748 258776 337754
rect 258724 337690 258776 337696
rect 258356 8288 258408 8294
rect 258356 8230 258408 8236
rect 258264 6248 258316 6254
rect 258264 6190 258316 6196
rect 258632 3936 258684 3942
rect 258632 3878 258684 3884
rect 258644 480 258672 3878
rect 258736 3330 258764 337690
rect 259380 337346 259408 340068
rect 259472 340054 260038 340082
rect 260300 340054 260590 340082
rect 259368 337340 259420 337346
rect 259368 337282 259420 337288
rect 259368 248396 259420 248402
rect 259368 248338 259420 248344
rect 259380 238785 259408 248338
rect 259366 238776 259422 238785
rect 259366 238711 259422 238720
rect 259366 87136 259422 87145
rect 259366 87071 259422 87080
rect 259380 86873 259408 87071
rect 259366 86864 259422 86873
rect 259366 86799 259422 86808
rect 259472 6322 259500 340054
rect 260300 333334 260328 340054
rect 261220 338026 261248 340068
rect 261208 338020 261260 338026
rect 261208 337962 261260 337968
rect 261312 335594 261340 340190
rect 262324 340054 262430 340082
rect 261484 337476 261536 337482
rect 261484 337418 261536 337424
rect 261036 335566 261340 335594
rect 259644 333328 259696 333334
rect 259644 333270 259696 333276
rect 260288 333328 260340 333334
rect 260288 333270 260340 333276
rect 259656 321638 259684 333270
rect 261036 321706 261064 335566
rect 261024 321700 261076 321706
rect 261024 321642 261076 321648
rect 259644 321632 259696 321638
rect 259644 321574 259696 321580
rect 261024 321564 261076 321570
rect 261024 321506 261076 321512
rect 261036 319025 261064 321506
rect 261022 319016 261078 319025
rect 261022 318951 261078 318960
rect 261022 318880 261078 318889
rect 259644 318844 259696 318850
rect 261022 318815 261078 318824
rect 259644 318786 259696 318792
rect 259656 318730 259684 318786
rect 259656 318702 259776 318730
rect 259748 292618 259776 318702
rect 261036 311930 261064 318815
rect 261036 311902 261156 311930
rect 261128 307834 261156 311902
rect 261024 307828 261076 307834
rect 261024 307770 261076 307776
rect 261116 307828 261168 307834
rect 261116 307770 261168 307776
rect 261036 307737 261064 307770
rect 261022 307728 261078 307737
rect 261022 307663 261078 307672
rect 261206 307728 261262 307737
rect 261206 307663 261262 307672
rect 261220 298178 261248 307663
rect 261024 298172 261076 298178
rect 261024 298114 261076 298120
rect 261208 298172 261260 298178
rect 261208 298114 261260 298120
rect 261036 298058 261064 298114
rect 261036 298030 261156 298058
rect 259656 292590 259776 292618
rect 259656 289814 259684 292590
rect 261128 292346 261156 298030
rect 261036 292318 261156 292346
rect 259644 289808 259696 289814
rect 259644 289750 259696 289756
rect 261036 280140 261064 292318
rect 260852 280112 261064 280140
rect 259736 277432 259788 277438
rect 259736 277374 259788 277380
rect 259748 267753 259776 277374
rect 260852 272898 260880 280112
rect 260852 272870 261064 272898
rect 259550 267744 259606 267753
rect 259550 267679 259606 267688
rect 259734 267744 259790 267753
rect 259734 267679 259790 267688
rect 259564 258097 259592 267679
rect 259550 258088 259606 258097
rect 259550 258023 259606 258032
rect 259734 258088 259790 258097
rect 259734 258023 259790 258032
rect 259748 254046 259776 258023
rect 261036 254046 261064 272870
rect 259736 254040 259788 254046
rect 259736 253982 259788 253988
rect 261024 254040 261076 254046
rect 261024 253982 261076 253988
rect 261024 253904 261076 253910
rect 261024 253846 261076 253852
rect 259644 248532 259696 248538
rect 259644 248474 259696 248480
rect 259656 248402 259684 248474
rect 259644 248396 259696 248402
rect 259644 248338 259696 248344
rect 261036 241482 261064 253846
rect 261036 241454 261156 241482
rect 259550 238776 259606 238785
rect 259550 238711 259606 238720
rect 259564 236586 259592 238711
rect 259564 236558 259684 236586
rect 259656 231810 259684 236558
rect 261128 234666 261156 241454
rect 261116 234660 261168 234666
rect 261116 234602 261168 234608
rect 261024 234592 261076 234598
rect 261024 234534 261076 234540
rect 259644 231804 259696 231810
rect 259644 231746 259696 231752
rect 259736 222216 259788 222222
rect 259736 222158 259788 222164
rect 261036 222170 261064 234534
rect 259748 217462 259776 222158
rect 261036 222142 261156 222170
rect 259736 217456 259788 217462
rect 259736 217398 259788 217404
rect 259644 217388 259696 217394
rect 259644 217330 259696 217336
rect 259656 212498 259684 217330
rect 261128 215354 261156 222142
rect 261116 215348 261168 215354
rect 261116 215290 261168 215296
rect 261024 215280 261076 215286
rect 261024 215222 261076 215228
rect 259644 212492 259696 212498
rect 259644 212434 259696 212440
rect 259736 202904 259788 202910
rect 259736 202846 259788 202852
rect 259748 198150 259776 202846
rect 259736 198144 259788 198150
rect 259736 198086 259788 198092
rect 259644 198076 259696 198082
rect 259644 198018 259696 198024
rect 259656 193225 259684 198018
rect 259642 193216 259698 193225
rect 259642 193151 259698 193160
rect 259826 193216 259882 193225
rect 259826 193151 259882 193160
rect 259840 173942 259868 193151
rect 261036 178786 261064 215222
rect 260944 178758 261064 178786
rect 259736 173936 259788 173942
rect 259736 173878 259788 173884
rect 259828 173936 259880 173942
rect 259828 173878 259880 173884
rect 259748 172514 259776 173878
rect 259736 172508 259788 172514
rect 259736 172450 259788 172456
rect 260944 166954 260972 178758
rect 260944 166926 261064 166954
rect 259644 162920 259696 162926
rect 259644 162862 259696 162868
rect 259656 149682 259684 162862
rect 259656 149654 259776 149682
rect 259748 143546 259776 149654
rect 259736 143540 259788 143546
rect 259736 143482 259788 143488
rect 259736 133816 259788 133822
rect 259736 133758 259788 133764
rect 259748 124370 259776 133758
rect 259736 124364 259788 124370
rect 259736 124306 259788 124312
rect 259736 124228 259788 124234
rect 259736 124170 259788 124176
rect 259748 122806 259776 124170
rect 259736 122800 259788 122806
rect 259736 122742 259788 122748
rect 259828 122800 259880 122806
rect 259828 122742 259880 122748
rect 259840 95266 259868 122742
rect 261036 99498 261064 166926
rect 260944 99470 261064 99498
rect 260944 99362 260972 99470
rect 260944 99334 261064 99362
rect 259644 95260 259696 95266
rect 259644 95202 259696 95208
rect 259828 95260 259880 95266
rect 259828 95202 259880 95208
rect 259656 89758 259684 95202
rect 259644 89752 259696 89758
rect 259644 89694 259696 89700
rect 259736 89616 259788 89622
rect 259736 89558 259788 89564
rect 259748 84182 259776 89558
rect 259736 84176 259788 84182
rect 259736 84118 259788 84124
rect 261036 80186 261064 99334
rect 261036 80158 261156 80186
rect 261128 79914 261156 80158
rect 261036 79886 261156 79914
rect 259644 71120 259696 71126
rect 259644 71062 259696 71068
rect 259656 60858 259684 71062
rect 259644 60852 259696 60858
rect 259644 60794 259696 60800
rect 261036 60738 261064 79886
rect 259644 60716 259696 60722
rect 259644 60658 259696 60664
rect 260944 60710 261064 60738
rect 259656 53122 259684 60658
rect 260944 60602 260972 60710
rect 260944 60574 261064 60602
rect 259656 53094 259776 53122
rect 259748 28966 259776 53094
rect 261036 51134 261064 60574
rect 261024 51128 261076 51134
rect 261024 51070 261076 51076
rect 261024 50992 261076 50998
rect 261024 50934 261076 50940
rect 261036 29102 261064 50934
rect 261024 29096 261076 29102
rect 261024 29038 261076 29044
rect 260932 29028 260984 29034
rect 260932 28970 260984 28976
rect 259552 28960 259604 28966
rect 259552 28902 259604 28908
rect 259736 28960 259788 28966
rect 259736 28902 259788 28908
rect 259564 19394 259592 28902
rect 259564 19366 259684 19394
rect 260944 19378 260972 28970
rect 259656 12594 259684 19366
rect 260932 19372 260984 19378
rect 260932 19314 260984 19320
rect 261024 19372 261076 19378
rect 261024 19314 261076 19320
rect 259656 12566 259776 12594
rect 259748 10305 259776 12566
rect 261036 12186 261064 19314
rect 260944 12158 261064 12186
rect 259734 10296 259790 10305
rect 259734 10231 259790 10240
rect 259828 8016 259880 8022
rect 259828 7958 259880 7964
rect 259460 6316 259512 6322
rect 259460 6258 259512 6264
rect 258724 3324 258776 3330
rect 258724 3266 258776 3272
rect 259840 480 259868 7958
rect 260944 6458 260972 12158
rect 260932 6452 260984 6458
rect 260932 6394 260984 6400
rect 261024 3460 261076 3466
rect 261024 3402 261076 3408
rect 261036 480 261064 3402
rect 261496 3262 261524 337418
rect 262324 10334 262352 340054
rect 262864 337544 262916 337550
rect 262864 337486 262916 337492
rect 262312 10328 262364 10334
rect 262312 10270 262364 10276
rect 262220 4072 262272 4078
rect 262220 4014 262272 4020
rect 261484 3256 261536 3262
rect 261484 3198 261536 3204
rect 262232 480 262260 4014
rect 262876 3194 262904 337486
rect 263060 337414 263088 340068
rect 263048 337408 263100 337414
rect 263048 337350 263100 337356
rect 263416 8084 263468 8090
rect 263416 8026 263468 8032
rect 262864 3188 262916 3194
rect 262864 3130 262916 3136
rect 263428 480 263456 8026
rect 263704 6390 263732 340068
rect 263796 340054 264270 340082
rect 263692 6384 263744 6390
rect 263692 6326 263744 6332
rect 263796 5302 263824 340054
rect 264900 338094 264928 340068
rect 264992 340054 265466 340082
rect 265636 340054 266110 340082
rect 264888 338088 264940 338094
rect 264888 338030 264940 338036
rect 264336 337680 264388 337686
rect 264336 337622 264388 337628
rect 264244 337476 264296 337482
rect 264244 337418 264296 337424
rect 263784 5296 263836 5302
rect 263784 5238 263836 5244
rect 264256 3126 264284 337418
rect 264244 3120 264296 3126
rect 264244 3062 264296 3068
rect 264348 3058 264376 337622
rect 264992 6526 265020 340054
rect 265636 328506 265664 340054
rect 266740 337754 266768 340068
rect 266728 337748 266780 337754
rect 266728 337690 266780 337696
rect 266832 335594 266860 340190
rect 266556 335566 266860 335594
rect 267844 340054 267950 340082
rect 265256 328500 265308 328506
rect 265256 328442 265308 328448
rect 265624 328500 265676 328506
rect 265624 328442 265676 328448
rect 265268 311930 265296 328442
rect 266556 321586 266584 335566
rect 267096 328500 267148 328506
rect 267096 328442 267148 328448
rect 266464 321558 266584 321586
rect 266464 321450 266492 321558
rect 266464 321422 266584 321450
rect 265176 311902 265296 311930
rect 265176 299538 265204 311902
rect 265164 299532 265216 299538
rect 265164 299474 265216 299480
rect 265256 299532 265308 299538
rect 265256 299474 265308 299480
rect 265268 298110 265296 299474
rect 265256 298104 265308 298110
rect 265256 298046 265308 298052
rect 266556 292618 266584 321422
rect 267108 309194 267136 328442
rect 267096 309188 267148 309194
rect 267096 309130 267148 309136
rect 267096 307828 267148 307834
rect 267096 307770 267148 307776
rect 267108 298110 267136 307770
rect 267096 298104 267148 298110
rect 267096 298046 267148 298052
rect 266464 292590 266584 292618
rect 266464 292482 266492 292590
rect 266464 292454 266584 292482
rect 265164 288448 265216 288454
rect 265164 288390 265216 288396
rect 265176 280514 265204 288390
rect 265176 280486 265296 280514
rect 265268 280226 265296 280486
rect 265072 280220 265124 280226
rect 265072 280162 265124 280168
rect 265256 280220 265308 280226
rect 265256 280162 265308 280168
rect 265084 278769 265112 280162
rect 265070 278760 265126 278769
rect 265070 278695 265126 278704
rect 265346 278760 265402 278769
rect 265346 278695 265402 278704
rect 265360 263514 265388 278695
rect 265268 263486 265388 263514
rect 265268 260846 265296 263486
rect 265256 260840 265308 260846
rect 265256 260782 265308 260788
rect 265256 251252 265308 251258
rect 265176 251212 265256 251240
rect 265176 244390 265204 251212
rect 265256 251194 265308 251200
rect 265164 244384 265216 244390
rect 265164 244326 265216 244332
rect 265164 244180 265216 244186
rect 265164 244122 265216 244128
rect 265176 232014 265204 244122
rect 265164 232008 265216 232014
rect 265164 231950 265216 231956
rect 265256 231872 265308 231878
rect 265256 231814 265308 231820
rect 265268 226930 265296 231814
rect 265176 226902 265296 226930
rect 265176 212702 265204 226902
rect 265164 212696 265216 212702
rect 265164 212638 265216 212644
rect 265256 212560 265308 212566
rect 265256 212502 265308 212508
rect 265268 205698 265296 212502
rect 265256 205692 265308 205698
rect 265256 205634 265308 205640
rect 265256 202904 265308 202910
rect 265256 202846 265308 202852
rect 265268 193322 265296 202846
rect 265256 193316 265308 193322
rect 265256 193258 265308 193264
rect 265164 193248 265216 193254
rect 265084 193196 265164 193202
rect 265084 193190 265216 193196
rect 265084 193174 265204 193190
rect 265084 186266 265112 193174
rect 265084 186238 265204 186266
rect 265176 182170 265204 186238
rect 265164 182164 265216 182170
rect 265164 182106 265216 182112
rect 265256 182164 265308 182170
rect 265256 182106 265308 182112
rect 265268 177313 265296 182106
rect 265254 177304 265310 177313
rect 265254 177239 265310 177248
rect 266556 173942 266584 292454
rect 267004 280220 267056 280226
rect 267004 280162 267056 280168
rect 267016 275210 267044 280162
rect 267016 275182 267136 275210
rect 267108 270502 267136 275182
rect 267096 270496 267148 270502
rect 267096 270438 267148 270444
rect 267096 260908 267148 260914
rect 267096 260850 267148 260856
rect 267108 253774 267136 260850
rect 267096 253768 267148 253774
rect 267096 253710 267148 253716
rect 267188 253700 267240 253706
rect 267188 253642 267240 253648
rect 267200 251240 267228 253642
rect 267108 251212 267228 251240
rect 267108 251138 267136 251212
rect 266924 251110 267136 251138
rect 266924 241534 266952 251110
rect 266820 241528 266872 241534
rect 266820 241470 266872 241476
rect 266912 241528 266964 241534
rect 266912 241470 266964 241476
rect 266832 240145 266860 241470
rect 266818 240136 266874 240145
rect 266818 240071 266874 240080
rect 267094 240136 267150 240145
rect 267094 240071 267150 240080
rect 267108 230489 267136 240071
rect 266726 230480 266782 230489
rect 266726 230415 266782 230424
rect 267094 230480 267150 230489
rect 267094 230415 267150 230424
rect 266740 220862 266768 230415
rect 266728 220856 266780 220862
rect 266728 220798 266780 220804
rect 266912 220856 266964 220862
rect 266912 220798 266964 220804
rect 266924 211154 266952 220798
rect 266924 211126 267044 211154
rect 267016 193254 267044 211126
rect 267004 193248 267056 193254
rect 267004 193190 267056 193196
rect 267096 193248 267148 193254
rect 267096 193190 267148 193196
rect 267108 188442 267136 193190
rect 267016 188414 267136 188442
rect 267016 183569 267044 188414
rect 267002 183560 267058 183569
rect 267002 183495 267058 183504
rect 267186 183560 267242 183569
rect 267186 183495 267242 183504
rect 267200 182170 267228 183495
rect 267188 182164 267240 182170
rect 267188 182106 267240 182112
rect 266452 173936 266504 173942
rect 266450 173904 266452 173913
rect 266544 173936 266596 173942
rect 266504 173904 266506 173913
rect 266544 173878 266596 173884
rect 266634 173904 266690 173913
rect 266450 173839 266506 173848
rect 266634 173839 266690 173848
rect 265254 164248 265310 164257
rect 265254 164183 265256 164192
rect 265308 164183 265310 164192
rect 265256 164154 265308 164160
rect 265164 154692 265216 154698
rect 265164 154634 265216 154640
rect 265176 147762 265204 154634
rect 266648 154630 266676 173839
rect 267188 173324 267240 173330
rect 267188 173266 267240 173272
rect 267200 164257 267228 173266
rect 267002 164248 267058 164257
rect 266912 164212 266964 164218
rect 267002 164183 267004 164192
rect 266912 164154 266964 164160
rect 267056 164183 267058 164192
rect 267186 164248 267242 164257
rect 267186 164183 267242 164192
rect 267004 164154 267056 164160
rect 266544 154624 266596 154630
rect 266544 154566 266596 154572
rect 266636 154624 266688 154630
rect 266924 154601 266952 164154
rect 266636 154566 266688 154572
rect 266910 154592 266966 154601
rect 265164 147756 265216 147762
rect 265164 147698 265216 147704
rect 265164 147620 265216 147626
rect 265164 147562 265216 147568
rect 265176 135425 265204 147562
rect 266556 145081 266584 154566
rect 266910 154527 266966 154536
rect 267094 154592 267150 154601
rect 267094 154527 267150 154536
rect 266542 145072 266598 145081
rect 266542 145007 266598 145016
rect 266450 144936 266506 144945
rect 266450 144871 266506 144880
rect 266464 143546 266492 144871
rect 266452 143540 266504 143546
rect 266452 143482 266504 143488
rect 266728 143540 266780 143546
rect 266728 143482 266780 143488
rect 265162 135416 265218 135425
rect 265162 135351 265218 135360
rect 265162 135280 265218 135289
rect 265162 135215 265218 135224
rect 265176 125610 265204 135215
rect 265176 125582 265296 125610
rect 265268 120766 265296 125582
rect 266740 122874 266768 143482
rect 267108 133090 267136 154527
rect 267738 134192 267794 134201
rect 267738 134127 267794 134136
rect 267752 134065 267780 134127
rect 267738 134056 267794 134065
rect 267738 133991 267794 134000
rect 267108 133062 267320 133090
rect 267292 132462 267320 133062
rect 267280 132456 267332 132462
rect 267280 132398 267332 132404
rect 266636 122868 266688 122874
rect 266636 122810 266688 122816
rect 266728 122868 266780 122874
rect 266728 122810 266780 122816
rect 267188 122868 267240 122874
rect 267188 122810 267240 122816
rect 265072 120760 265124 120766
rect 265072 120702 265124 120708
rect 265256 120760 265308 120766
rect 265256 120702 265308 120708
rect 265084 115977 265112 120702
rect 265070 115968 265126 115977
rect 265070 115903 265126 115912
rect 265254 115968 265310 115977
rect 265254 115903 265310 115912
rect 265268 100042 265296 115903
rect 266648 113234 266676 122810
rect 267200 117842 267228 122810
rect 266912 117836 266964 117842
rect 266912 117778 266964 117784
rect 267188 117836 267240 117842
rect 267188 117778 267240 117784
rect 266464 113206 266676 113234
rect 266464 109154 266492 113206
rect 266464 109126 266676 109154
rect 266648 103578 266676 109126
rect 266556 103550 266676 103578
rect 266556 102134 266584 103550
rect 266544 102128 266596 102134
rect 266544 102070 266596 102076
rect 265176 100014 265296 100042
rect 265176 77466 265204 100014
rect 266924 95266 266952 117778
rect 266912 95260 266964 95266
rect 266912 95202 266964 95208
rect 267096 95260 267148 95266
rect 267096 95202 267148 95208
rect 266452 92540 266504 92546
rect 266452 92482 266504 92488
rect 266464 82793 266492 92482
rect 267108 87038 267136 95202
rect 267740 87168 267792 87174
rect 267738 87136 267740 87145
rect 267792 87136 267794 87145
rect 267738 87071 267794 87080
rect 267096 87032 267148 87038
rect 267096 86974 267148 86980
rect 267004 86964 267056 86970
rect 267004 86906 267056 86912
rect 266450 82784 266506 82793
rect 266450 82719 266506 82728
rect 266634 82648 266690 82657
rect 266634 82583 266690 82592
rect 266648 77994 266676 82583
rect 266636 77988 266688 77994
rect 266636 77930 266688 77936
rect 265176 77438 265296 77466
rect 265268 77296 265296 77438
rect 265176 77268 265296 77296
rect 265176 66298 265204 77268
rect 267016 74662 267044 86906
rect 267004 74656 267056 74662
rect 267004 74598 267056 74604
rect 266820 74520 266872 74526
rect 266820 74462 266872 74468
rect 265164 66292 265216 66298
rect 265164 66234 265216 66240
rect 265256 66292 265308 66298
rect 265256 66234 265308 66240
rect 265268 28966 265296 66234
rect 266452 64932 266504 64938
rect 266452 64874 266504 64880
rect 266464 51762 266492 64874
rect 266832 55282 266860 74462
rect 267648 63912 267700 63918
rect 267646 63880 267648 63889
rect 267700 63880 267702 63889
rect 267646 63815 267702 63824
rect 266820 55276 266872 55282
rect 266820 55218 266872 55224
rect 267004 55276 267056 55282
rect 267004 55218 267056 55224
rect 267016 55146 267044 55218
rect 267004 55140 267056 55146
rect 267004 55082 267056 55088
rect 266464 51734 266584 51762
rect 266556 28966 266584 51734
rect 267096 45620 267148 45626
rect 267096 45562 267148 45568
rect 267108 42090 267136 45562
rect 267096 42084 267148 42090
rect 267096 42026 267148 42032
rect 267740 40384 267792 40390
rect 267738 40352 267740 40361
rect 267792 40352 267794 40361
rect 267738 40287 267794 40296
rect 267096 29028 267148 29034
rect 267096 28970 267148 28976
rect 265164 28960 265216 28966
rect 265164 28902 265216 28908
rect 265256 28960 265308 28966
rect 265256 28902 265308 28908
rect 266544 28960 266596 28966
rect 266544 28902 266596 28908
rect 266636 28960 266688 28966
rect 266636 28902 266688 28908
rect 265176 14550 265204 28902
rect 266648 27606 266676 28902
rect 266636 27600 266688 27606
rect 266636 27542 266688 27548
rect 266636 19236 266688 19242
rect 266636 19178 266688 19184
rect 265164 14544 265216 14550
rect 266648 14498 266676 19178
rect 265164 14486 265216 14492
rect 266372 14470 266676 14498
rect 266372 6594 266400 14470
rect 267108 9602 267136 28970
rect 267844 14618 267872 340054
rect 268384 337884 268436 337890
rect 268384 337826 268436 337832
rect 267832 14612 267884 14618
rect 267832 14554 267884 14560
rect 266924 9574 267136 9602
rect 266360 6588 266412 6594
rect 266360 6530 266412 6536
rect 264980 6520 265032 6526
rect 264980 6462 265032 6468
rect 264612 3732 264664 3738
rect 264612 3674 264664 3680
rect 264336 3052 264388 3058
rect 264336 2994 264388 3000
rect 264624 480 264652 3674
rect 265808 3528 265860 3534
rect 265808 3470 265860 3476
rect 265820 480 265848 3470
rect 266924 2990 266952 9574
rect 267004 8152 267056 8158
rect 267004 8094 267056 8100
rect 266912 2984 266964 2990
rect 266912 2926 266964 2932
rect 267016 480 267044 8094
rect 268108 3392 268160 3398
rect 268108 3334 268160 3340
rect 268120 480 268148 3334
rect 268396 2922 268424 337826
rect 268580 336802 268608 340068
rect 268568 336796 268620 336802
rect 268568 336738 268620 336744
rect 268934 171320 268990 171329
rect 268934 171255 268990 171264
rect 268948 170105 268976 171255
rect 268934 170096 268990 170105
rect 268934 170031 268990 170040
rect 269132 6662 269160 340068
rect 269224 340054 269790 340082
rect 269224 14686 269252 340054
rect 269764 337816 269816 337822
rect 269764 337758 269816 337764
rect 269212 14680 269264 14686
rect 269212 14622 269264 14628
rect 269120 6656 269172 6662
rect 269120 6598 269172 6604
rect 269304 3664 269356 3670
rect 269304 3606 269356 3612
rect 268384 2916 268436 2922
rect 268384 2858 268436 2864
rect 269316 480 269344 3606
rect 269776 2854 269804 337758
rect 270420 337346 270448 340068
rect 270512 340054 270986 340082
rect 271156 340054 271630 340082
rect 270408 337340 270460 337346
rect 270408 337282 270460 337288
rect 270512 9602 270540 340054
rect 271156 328506 271184 340054
rect 272260 337278 272288 340068
rect 272444 340054 272826 340082
rect 273364 340054 273470 340082
rect 272248 337272 272300 337278
rect 272248 337214 272300 337220
rect 272444 335730 272472 340054
rect 272076 335702 272472 335730
rect 270776 328500 270828 328506
rect 270776 328442 270828 328448
rect 271144 328500 271196 328506
rect 271144 328442 271196 328448
rect 270788 311930 270816 328442
rect 272076 321586 272104 335702
rect 271984 321558 272104 321586
rect 271984 321450 272012 321558
rect 271984 321422 272104 321450
rect 270696 311902 270816 311930
rect 270696 309126 270724 311902
rect 270684 309120 270736 309126
rect 270684 309062 270736 309068
rect 270776 299532 270828 299538
rect 270776 299474 270828 299480
rect 270788 298110 270816 299474
rect 270776 298104 270828 298110
rect 270776 298046 270828 298052
rect 270868 298104 270920 298110
rect 270868 298046 270920 298052
rect 270880 280158 270908 298046
rect 272076 292618 272104 321422
rect 271984 292590 272104 292618
rect 271984 292482 272012 292590
rect 271984 292454 272104 292482
rect 270592 280152 270644 280158
rect 270592 280094 270644 280100
rect 270868 280152 270920 280158
rect 270868 280094 270920 280100
rect 270604 278730 270632 280094
rect 270592 278724 270644 278730
rect 270592 278666 270644 278672
rect 272076 273222 272104 292454
rect 272064 273216 272116 273222
rect 272064 273158 272116 273164
rect 272064 273080 272116 273086
rect 272064 273022 272116 273028
rect 270776 260908 270828 260914
rect 270776 260850 270828 260856
rect 270788 260817 270816 260850
rect 272076 260846 272104 273022
rect 272064 260840 272116 260846
rect 270774 260808 270830 260817
rect 270774 260743 270830 260752
rect 270958 260808 271014 260817
rect 272064 260782 272116 260788
rect 270958 260743 271014 260752
rect 270972 251258 271000 260743
rect 270684 251252 270736 251258
rect 270684 251194 270736 251200
rect 270960 251252 271012 251258
rect 270960 251194 271012 251200
rect 272064 251252 272116 251258
rect 272064 251194 272116 251200
rect 270696 244322 270724 251194
rect 270684 244316 270736 244322
rect 270684 244258 270736 244264
rect 270776 244180 270828 244186
rect 270776 244122 270828 244128
rect 270788 241482 270816 244122
rect 272076 241505 272104 251194
rect 270696 241454 270816 241482
rect 271878 241496 271934 241505
rect 270696 234818 270724 241454
rect 271878 241431 271934 241440
rect 272062 241496 272118 241505
rect 272062 241431 272118 241440
rect 270604 234790 270724 234818
rect 270604 230518 270632 234790
rect 271892 231878 271920 241431
rect 271880 231872 271932 231878
rect 271880 231814 271932 231820
rect 272064 231872 272116 231878
rect 272064 231814 272116 231820
rect 270592 230512 270644 230518
rect 270592 230454 270644 230460
rect 270684 230512 270736 230518
rect 270736 230460 270816 230466
rect 270684 230454 270816 230460
rect 270696 230438 270816 230454
rect 270788 225010 270816 230438
rect 270776 225004 270828 225010
rect 270776 224946 270828 224952
rect 270684 224936 270736 224942
rect 270684 224878 270736 224884
rect 270696 215422 270724 224878
rect 272076 222193 272104 231814
rect 271878 222184 271934 222193
rect 271878 222119 271934 222128
rect 272062 222184 272118 222193
rect 272062 222119 272118 222128
rect 270684 215416 270736 215422
rect 270684 215358 270736 215364
rect 271892 212566 271920 222119
rect 271880 212560 271932 212566
rect 271880 212502 271932 212508
rect 272064 212560 272116 212566
rect 272064 212502 272116 212508
rect 270684 212492 270736 212498
rect 270684 212434 270736 212440
rect 270696 211138 270724 212434
rect 270684 211132 270736 211138
rect 270684 211074 270736 211080
rect 270684 205624 270736 205630
rect 270684 205566 270736 205572
rect 270696 201498 270724 205566
rect 270696 201470 270816 201498
rect 270788 196110 270816 201470
rect 270776 196104 270828 196110
rect 272076 196058 272104 212502
rect 270776 196046 270828 196052
rect 271984 196030 272104 196058
rect 271984 195922 272012 196030
rect 271984 195894 272104 195922
rect 270592 193180 270644 193186
rect 270592 193122 270644 193128
rect 270604 191826 270632 193122
rect 270592 191820 270644 191826
rect 270592 191762 270644 191768
rect 272076 186454 272104 195894
rect 272064 186448 272116 186454
rect 272064 186390 272116 186396
rect 271972 183592 272024 183598
rect 271972 183534 272024 183540
rect 270684 183524 270736 183530
rect 270684 183466 270736 183472
rect 270696 182186 270724 183466
rect 270696 182158 270816 182186
rect 270788 178786 270816 182158
rect 270788 178758 270908 178786
rect 270880 173942 270908 178758
rect 271984 173942 272012 183534
rect 270684 173936 270736 173942
rect 270684 173878 270736 173884
rect 270868 173936 270920 173942
rect 270868 173878 270920 173884
rect 271972 173936 272024 173942
rect 271972 173878 272024 173884
rect 272064 173936 272116 173942
rect 272064 173878 272116 173884
rect 270696 167074 270724 173878
rect 272076 172514 272104 173878
rect 272064 172508 272116 172514
rect 272064 172450 272116 172456
rect 270684 167068 270736 167074
rect 270684 167010 270736 167016
rect 270776 166932 270828 166938
rect 270776 166874 270828 166880
rect 270788 138258 270816 166874
rect 271972 162920 272024 162926
rect 271972 162862 272024 162868
rect 271984 158030 272012 162862
rect 271972 158024 272024 158030
rect 271972 157966 272024 157972
rect 271972 148640 272024 148646
rect 271972 148582 272024 148588
rect 271984 144906 272012 148582
rect 271972 144900 272024 144906
rect 271972 144842 272024 144848
rect 272064 144900 272116 144906
rect 272064 144842 272116 144848
rect 272076 139890 272104 144842
rect 271984 139862 272104 139890
rect 270788 138230 270908 138258
rect 270880 135289 270908 138230
rect 270682 135280 270738 135289
rect 270682 135215 270738 135224
rect 270866 135280 270922 135289
rect 271984 135250 272012 139862
rect 270866 135215 270922 135224
rect 271880 135244 271932 135250
rect 270696 130370 270724 135215
rect 271880 135186 271932 135192
rect 271972 135244 272024 135250
rect 271972 135186 272024 135192
rect 270696 130342 270816 130370
rect 270788 125594 270816 130342
rect 271892 125633 271920 135186
rect 271878 125624 271934 125633
rect 270592 125588 270644 125594
rect 270592 125530 270644 125536
rect 270776 125588 270828 125594
rect 272062 125624 272118 125633
rect 271878 125559 271934 125568
rect 271972 125588 272024 125594
rect 270776 125530 270828 125536
rect 272062 125559 272064 125568
rect 271972 125530 272024 125536
rect 272116 125559 272118 125568
rect 272064 125530 272116 125536
rect 270604 118674 270632 125530
rect 271984 124166 272012 125530
rect 271972 124160 272024 124166
rect 271972 124102 272024 124108
rect 270604 118646 270724 118674
rect 270696 106298 270724 118646
rect 271972 115388 272024 115394
rect 271972 115330 272024 115336
rect 270696 106270 270816 106298
rect 270788 95441 270816 106270
rect 271984 104922 272012 115330
rect 271880 104916 271932 104922
rect 271880 104858 271932 104864
rect 271972 104916 272024 104922
rect 271972 104858 272024 104864
rect 271892 99346 271920 104858
rect 271880 99340 271932 99346
rect 271880 99282 271932 99288
rect 272064 99340 272116 99346
rect 272064 99282 272116 99288
rect 270774 95432 270830 95441
rect 270774 95367 270830 95376
rect 270682 95296 270738 95305
rect 270682 95231 270738 95240
rect 270696 90386 270724 95231
rect 270604 90358 270724 90386
rect 270604 86902 270632 90358
rect 270592 86896 270644 86902
rect 270592 86838 270644 86844
rect 270868 86896 270920 86902
rect 270868 86838 270920 86844
rect 270880 77314 270908 86838
rect 272076 84318 272104 99282
rect 272064 84312 272116 84318
rect 272064 84254 272116 84260
rect 271972 84244 272024 84250
rect 271972 84186 272024 84192
rect 271984 82822 272012 84186
rect 271972 82816 272024 82822
rect 271972 82758 272024 82764
rect 270684 77308 270736 77314
rect 270684 77250 270736 77256
rect 270868 77308 270920 77314
rect 270868 77250 270920 77256
rect 270696 75886 270724 77250
rect 270684 75880 270736 75886
rect 270684 75822 270736 75828
rect 271972 73228 272024 73234
rect 271972 73170 272024 73176
rect 270776 66292 270828 66298
rect 270776 66234 270828 66240
rect 270788 60858 270816 66234
rect 271984 64870 272012 73170
rect 271972 64864 272024 64870
rect 271972 64806 272024 64812
rect 272064 64864 272116 64870
rect 272064 64806 272116 64812
rect 270776 60852 270828 60858
rect 270776 60794 270828 60800
rect 270684 60716 270736 60722
rect 270684 60658 270736 60664
rect 270696 47054 270724 60658
rect 272076 51814 272104 64806
rect 272064 51808 272116 51814
rect 272064 51750 272116 51756
rect 270684 47048 270736 47054
rect 270684 46990 270736 46996
rect 270592 46980 270644 46986
rect 270592 46922 270644 46928
rect 271972 46980 272024 46986
rect 271972 46922 272024 46928
rect 270604 38706 270632 46922
rect 271984 42974 272012 46922
rect 271972 42968 272024 42974
rect 271972 42910 272024 42916
rect 270604 38678 270724 38706
rect 270696 29034 270724 38678
rect 270684 29028 270736 29034
rect 270684 28970 270736 28976
rect 270776 29028 270828 29034
rect 270776 28970 270828 28976
rect 272064 29028 272116 29034
rect 272064 28970 272116 28976
rect 270788 27606 270816 28970
rect 270776 27600 270828 27606
rect 270776 27542 270828 27548
rect 272076 18086 272104 28970
rect 272064 18080 272116 18086
rect 272064 18022 272116 18028
rect 270684 18012 270736 18018
rect 270684 17954 270736 17960
rect 271972 18012 272024 18018
rect 271972 17954 272024 17960
rect 270696 14754 270724 17954
rect 270684 14748 270736 14754
rect 270684 14690 270736 14696
rect 271984 13138 272012 17954
rect 273364 14822 273392 340054
rect 274100 336870 274128 340068
rect 274088 336864 274140 336870
rect 274088 336806 274140 336812
rect 273720 87168 273772 87174
rect 273718 87136 273720 87145
rect 273772 87136 273774 87145
rect 273718 87071 273774 87080
rect 274086 29200 274142 29209
rect 274270 29200 274326 29209
rect 274142 29158 274270 29186
rect 274086 29135 274142 29144
rect 274270 29135 274326 29144
rect 273352 14816 273404 14822
rect 273352 14758 273404 14764
rect 271800 13110 272012 13138
rect 271800 12322 271828 13110
rect 271800 12294 271920 12322
rect 270512 9574 270632 9602
rect 270500 8220 270552 8226
rect 270500 8162 270552 8168
rect 269764 2848 269816 2854
rect 269764 2790 269816 2796
rect 270512 480 270540 8162
rect 270604 6730 270632 9574
rect 271892 6798 271920 12294
rect 274088 8288 274140 8294
rect 274088 8230 274140 8236
rect 271880 6792 271932 6798
rect 271880 6734 271932 6740
rect 270592 6724 270644 6730
rect 270592 6666 270644 6672
rect 271696 4004 271748 4010
rect 271696 3946 271748 3952
rect 271708 480 271736 3946
rect 272892 3800 272944 3806
rect 272892 3742 272944 3748
rect 272904 480 272932 3742
rect 274100 480 274128 8230
rect 274652 7546 274680 340068
rect 274744 340054 275310 340082
rect 274744 14890 274772 340054
rect 275940 337414 275968 340068
rect 276032 340054 276506 340082
rect 276584 340054 277150 340082
rect 275928 337408 275980 337414
rect 275928 337350 275980 337356
rect 275928 63912 275980 63918
rect 275926 63880 275928 63889
rect 275980 63880 275982 63889
rect 275926 63815 275982 63824
rect 274732 14884 274784 14890
rect 274732 14826 274784 14832
rect 274640 7540 274692 7546
rect 274640 7482 274692 7488
rect 276032 7478 276060 340054
rect 276584 335730 276612 340054
rect 276664 337408 276716 337414
rect 276664 337350 276716 337356
rect 276124 335702 276612 335730
rect 276124 14958 276152 335702
rect 276112 14952 276164 14958
rect 276112 14894 276164 14900
rect 276020 7472 276072 7478
rect 276020 7414 276072 7420
rect 276480 4140 276532 4146
rect 276480 4082 276532 4088
rect 275284 3596 275336 3602
rect 275284 3538 275336 3544
rect 275296 480 275324 3538
rect 276492 480 276520 4082
rect 276676 3602 276704 337350
rect 277780 337210 277808 340068
rect 277964 340054 278346 340082
rect 278884 340054 278990 340082
rect 277768 337204 277820 337210
rect 277768 337146 277820 337152
rect 277964 335730 277992 340054
rect 277596 335702 277992 335730
rect 277596 323610 277624 335702
rect 277308 323604 277360 323610
rect 277308 323546 277360 323552
rect 277584 323604 277636 323610
rect 277584 323546 277636 323552
rect 277320 318889 277348 323546
rect 277306 318880 277362 318889
rect 277306 318815 277362 318824
rect 277582 318880 277638 318889
rect 277582 318815 277638 318824
rect 277596 311982 277624 318815
rect 277584 311976 277636 311982
rect 277584 311918 277636 311924
rect 277492 309052 277544 309058
rect 277492 308994 277544 309000
rect 277504 307850 277532 308994
rect 277504 307822 277624 307850
rect 277596 307766 277624 307822
rect 277584 307760 277636 307766
rect 277584 307702 277636 307708
rect 277584 298240 277636 298246
rect 277584 298182 277636 298188
rect 277596 298110 277624 298182
rect 277584 298104 277636 298110
rect 277584 298046 277636 298052
rect 277676 280220 277728 280226
rect 277676 280162 277728 280168
rect 277688 270473 277716 280162
rect 277674 270464 277730 270473
rect 277674 270399 277730 270408
rect 277766 270328 277822 270337
rect 277766 270263 277822 270272
rect 277780 260930 277808 270263
rect 277596 260902 277808 260930
rect 277596 260846 277624 260902
rect 277584 260840 277636 260846
rect 277584 260782 277636 260788
rect 277676 260840 277728 260846
rect 277676 260782 277728 260788
rect 277688 244202 277716 260782
rect 277596 244174 277716 244202
rect 277596 231878 277624 244174
rect 277584 231872 277636 231878
rect 277584 231814 277636 231820
rect 277676 231872 277728 231878
rect 277676 231814 277728 231820
rect 277688 224890 277716 231814
rect 277596 224862 277716 224890
rect 277596 212566 277624 224862
rect 277584 212560 277636 212566
rect 277584 212502 277636 212508
rect 277676 212560 277728 212566
rect 277676 212502 277728 212508
rect 277688 205578 277716 212502
rect 278686 208584 278742 208593
rect 278686 208519 278742 208528
rect 277596 205550 277716 205578
rect 277596 196058 277624 205550
rect 278700 204649 278728 208519
rect 278686 204640 278742 204649
rect 278686 204575 278742 204584
rect 277504 196030 277624 196058
rect 277504 195974 277532 196030
rect 277492 195968 277544 195974
rect 277492 195910 277544 195916
rect 277676 195968 277728 195974
rect 277676 195910 277728 195916
rect 277688 186454 277716 195910
rect 277676 186448 277728 186454
rect 277676 186390 277728 186396
rect 277676 186244 277728 186250
rect 277676 186186 277728 186192
rect 277688 183546 277716 186186
rect 277596 183518 277716 183546
rect 277596 167090 277624 183518
rect 277504 167062 277624 167090
rect 277504 166954 277532 167062
rect 277504 166926 277624 166954
rect 277596 147778 277624 166926
rect 278686 157584 278742 157593
rect 278686 157519 278742 157528
rect 278700 157457 278728 157519
rect 278686 157448 278742 157457
rect 278686 157383 278742 157392
rect 277504 147750 277624 147778
rect 277504 147642 277532 147750
rect 277504 147614 277716 147642
rect 277688 138106 277716 147614
rect 277676 138100 277728 138106
rect 277676 138042 277728 138048
rect 277584 137964 277636 137970
rect 277584 137906 277636 137912
rect 277596 116113 277624 137906
rect 278686 134192 278742 134201
rect 278686 134127 278742 134136
rect 278700 133929 278728 134127
rect 278686 133920 278742 133929
rect 278686 133855 278742 133864
rect 277582 116104 277638 116113
rect 277582 116039 277638 116048
rect 277490 115968 277546 115977
rect 277490 115903 277492 115912
rect 277544 115903 277546 115912
rect 277676 115932 277728 115938
rect 277492 115874 277544 115880
rect 277676 115874 277728 115880
rect 277688 110922 277716 115874
rect 277596 110894 277716 110922
rect 278778 110936 278834 110945
rect 277596 99482 277624 110894
rect 278778 110871 278834 110880
rect 278792 110537 278820 110871
rect 278778 110528 278834 110537
rect 278778 110463 278834 110472
rect 277584 99476 277636 99482
rect 277584 99418 277636 99424
rect 277584 99340 277636 99346
rect 277584 99282 277636 99288
rect 277596 70514 277624 99282
rect 277584 70508 277636 70514
rect 277584 70450 277636 70456
rect 277584 70372 277636 70378
rect 277584 70314 277636 70320
rect 277306 63880 277362 63889
rect 277306 63815 277362 63824
rect 277320 63617 277348 63815
rect 277306 63608 277362 63617
rect 277306 63543 277362 63552
rect 277596 51762 277624 70314
rect 277596 51734 277716 51762
rect 277308 40384 277360 40390
rect 277306 40352 277308 40361
rect 277360 40352 277362 40361
rect 277306 40287 277362 40296
rect 277688 29050 277716 51734
rect 278686 40352 278742 40361
rect 278686 40287 278742 40296
rect 278700 40089 278728 40287
rect 278686 40080 278742 40089
rect 278686 40015 278742 40024
rect 278780 29232 278832 29238
rect 278778 29200 278780 29209
rect 278832 29200 278834 29209
rect 278778 29135 278834 29144
rect 277596 29022 277716 29050
rect 277596 22166 277624 29022
rect 277584 22160 277636 22166
rect 277584 22102 277636 22108
rect 277492 22092 277544 22098
rect 277492 22034 277544 22040
rect 277504 7410 277532 22034
rect 278884 15026 278912 340054
rect 279620 337482 279648 340068
rect 279608 337476 279660 337482
rect 279608 337418 279660 337424
rect 280068 337476 280120 337482
rect 280068 337418 280120 337424
rect 278872 15020 278924 15026
rect 278872 14962 278924 14968
rect 277676 7540 277728 7546
rect 277676 7482 277728 7488
rect 277492 7404 277544 7410
rect 277492 7346 277544 7352
rect 276664 3596 276716 3602
rect 276664 3538 276716 3544
rect 277688 480 277716 7482
rect 279976 6180 280028 6186
rect 279976 6122 280028 6128
rect 278872 3392 278924 3398
rect 278872 3334 278924 3340
rect 278884 480 278912 3334
rect 279988 3074 280016 6122
rect 280080 3398 280108 337418
rect 280172 10402 280200 340068
rect 280264 340054 280830 340082
rect 280264 15094 280292 340054
rect 281460 337686 281488 340068
rect 281552 340054 282026 340082
rect 282104 340054 282670 340082
rect 281448 337680 281500 337686
rect 281448 337622 281500 337628
rect 280252 15088 280304 15094
rect 280252 15030 280304 15036
rect 281552 10470 281580 340054
rect 282104 331922 282132 340054
rect 283208 337142 283236 340068
rect 283196 337136 283248 337142
rect 283196 337078 283248 337084
rect 283300 335594 283328 340190
rect 284404 340054 284510 340082
rect 283564 337680 283616 337686
rect 283564 337622 283616 337628
rect 281920 331894 282132 331922
rect 283116 335566 283328 335594
rect 281920 330290 281948 331894
rect 281920 330262 282040 330290
rect 282012 327078 282040 330262
rect 281632 327072 281684 327078
rect 281632 327014 281684 327020
rect 282000 327072 282052 327078
rect 282000 327014 282052 327020
rect 281644 317422 281672 327014
rect 283116 318782 283144 335566
rect 283012 318776 283064 318782
rect 283012 318718 283064 318724
rect 283104 318776 283156 318782
rect 283104 318718 283156 318724
rect 283024 317422 283052 318718
rect 281632 317416 281684 317422
rect 281632 317358 281684 317364
rect 283012 317416 283064 317422
rect 283012 317358 283064 317364
rect 281632 307828 281684 307834
rect 281632 307770 281684 307776
rect 283012 307828 283064 307834
rect 283012 307770 283064 307776
rect 281644 302326 281672 307770
rect 283024 302326 283052 307770
rect 281632 302320 281684 302326
rect 281632 302262 281684 302268
rect 283012 302320 283064 302326
rect 283012 302262 283064 302268
rect 281816 302116 281868 302122
rect 281816 302058 281868 302064
rect 283104 302116 283156 302122
rect 283104 302058 283156 302064
rect 281828 299470 281856 302058
rect 283116 299470 283144 302058
rect 281816 299464 281868 299470
rect 281816 299406 281868 299412
rect 283104 299464 283156 299470
rect 283104 299406 283156 299412
rect 281632 289876 281684 289882
rect 281632 289818 281684 289824
rect 283104 289876 283156 289882
rect 283104 289818 283156 289824
rect 281644 289785 281672 289818
rect 281630 289776 281686 289785
rect 281630 289711 281686 289720
rect 281906 289776 281962 289785
rect 281906 289711 281962 289720
rect 281920 280226 281948 289711
rect 281724 280220 281776 280226
rect 281724 280162 281776 280168
rect 281908 280220 281960 280226
rect 281908 280162 281960 280168
rect 281736 280106 281764 280162
rect 281736 280078 281856 280106
rect 281828 269074 281856 280078
rect 283116 273222 283144 289818
rect 283104 273216 283156 273222
rect 283104 273158 283156 273164
rect 283104 273080 283156 273086
rect 283104 273022 283156 273028
rect 281816 269068 281868 269074
rect 281816 269010 281868 269016
rect 282000 259480 282052 259486
rect 282000 259422 282052 259428
rect 282012 248402 282040 259422
rect 283116 253910 283144 273022
rect 283104 253904 283156 253910
rect 283104 253846 283156 253852
rect 283104 253768 283156 253774
rect 283104 253710 283156 253716
rect 282000 248396 282052 248402
rect 282000 248338 282052 248344
rect 282184 248396 282236 248402
rect 282184 248338 282236 248344
rect 282196 238785 282224 248338
rect 281906 238776 281962 238785
rect 281906 238711 281962 238720
rect 282182 238776 282238 238785
rect 282182 238711 282238 238720
rect 281920 234734 281948 238711
rect 281908 234728 281960 234734
rect 283116 234682 283144 253710
rect 281908 234670 281960 234676
rect 283024 234654 283144 234682
rect 281816 234592 281868 234598
rect 281816 234534 281868 234540
rect 283024 234546 283052 234654
rect 281828 229090 281856 234534
rect 283024 234518 283144 234546
rect 281816 229084 281868 229090
rect 281816 229026 281868 229032
rect 283116 215286 283144 234518
rect 283104 215280 283156 215286
rect 283104 215222 283156 215228
rect 283104 215144 283156 215150
rect 283104 215086 283156 215092
rect 281816 212492 281868 212498
rect 281816 212434 281868 212440
rect 281828 211154 281856 212434
rect 281828 211126 281948 211154
rect 281920 202910 281948 211126
rect 281724 202904 281776 202910
rect 281722 202872 281724 202881
rect 281908 202904 281960 202910
rect 281776 202872 281778 202881
rect 281722 202807 281778 202816
rect 281906 202872 281908 202881
rect 281960 202872 281962 202881
rect 281906 202807 281962 202816
rect 281920 201482 281948 202807
rect 281908 201476 281960 201482
rect 281908 201418 281960 201424
rect 281908 193180 281960 193186
rect 281908 193122 281960 193128
rect 281920 191842 281948 193122
rect 281920 191814 282040 191842
rect 282012 183705 282040 191814
rect 281998 183696 282054 183705
rect 281998 183631 282054 183640
rect 281998 183424 282054 183433
rect 281998 183359 282054 183368
rect 282012 176338 282040 183359
rect 281828 176310 282040 176338
rect 281828 159066 281856 176310
rect 283116 167090 283144 215086
rect 283024 167062 283144 167090
rect 283024 166954 283052 167062
rect 283024 166926 283144 166954
rect 281736 159038 281856 159066
rect 281736 153202 281764 159038
rect 283116 154737 283144 166926
rect 283102 154728 283158 154737
rect 283102 154663 283158 154672
rect 283102 154592 283158 154601
rect 283102 154527 283158 154536
rect 281724 153196 281776 153202
rect 281724 153138 281776 153144
rect 281816 153196 281868 153202
rect 281816 153138 281868 153144
rect 281828 118810 281856 153138
rect 283116 144974 283144 154527
rect 283104 144968 283156 144974
rect 283104 144910 283156 144916
rect 283012 144900 283064 144906
rect 283012 144842 283064 144848
rect 283024 142118 283052 144842
rect 283012 142112 283064 142118
rect 283012 142054 283064 142060
rect 283104 132524 283156 132530
rect 283104 132466 283156 132472
rect 283116 125769 283144 132466
rect 283102 125760 283158 125769
rect 283102 125695 283158 125704
rect 283102 125624 283158 125633
rect 283102 125559 283158 125568
rect 281736 118782 281856 118810
rect 283116 118810 283144 125559
rect 283116 118782 283236 118810
rect 281736 109154 281764 118782
rect 283208 114578 283236 118782
rect 283104 114572 283156 114578
rect 283104 114514 283156 114520
rect 283196 114572 283248 114578
rect 283196 114514 283248 114520
rect 283116 109750 283144 114514
rect 282920 109744 282972 109750
rect 282920 109686 282972 109692
rect 283104 109744 283156 109750
rect 283104 109686 283156 109692
rect 281736 109126 281856 109154
rect 281828 106321 281856 109126
rect 281630 106312 281686 106321
rect 281630 106247 281632 106256
rect 281684 106247 281686 106256
rect 281814 106312 281870 106321
rect 281814 106247 281870 106256
rect 281632 106218 281684 106224
rect 282932 104854 282960 109686
rect 282920 104848 282972 104854
rect 282920 104790 282972 104796
rect 281632 101380 281684 101386
rect 281632 101322 281684 101328
rect 281644 96642 281672 101322
rect 281644 96614 281764 96642
rect 281736 91746 281764 96614
rect 282920 95260 282972 95266
rect 282920 95202 282972 95208
rect 282932 91746 282960 95202
rect 281736 91718 281856 91746
rect 282932 91718 283144 91746
rect 281828 89706 281856 91718
rect 281736 89678 281856 89706
rect 281736 77314 281764 89678
rect 281724 77308 281776 77314
rect 281724 77250 281776 77256
rect 281724 75948 281776 75954
rect 281724 75890 281776 75896
rect 281736 67590 281764 75890
rect 283116 70666 283144 91718
rect 283472 76016 283524 76022
rect 283470 75984 283472 75993
rect 283524 75984 283526 75993
rect 283470 75919 283526 75928
rect 283116 70638 283236 70666
rect 281724 67584 281776 67590
rect 281724 67526 281776 67532
rect 283208 66366 283236 70638
rect 283196 66360 283248 66366
rect 283196 66302 283248 66308
rect 281724 61464 281776 61470
rect 281724 61406 281776 61412
rect 281736 56574 281764 61406
rect 283104 56636 283156 56642
rect 283104 56578 283156 56584
rect 281724 56568 281776 56574
rect 281724 56510 281776 56516
rect 281632 46980 281684 46986
rect 281632 46922 281684 46928
rect 281644 46866 281672 46922
rect 283116 46900 283144 56578
rect 283116 46872 283236 46900
rect 281644 46838 281764 46866
rect 281736 28966 281764 46838
rect 283208 45558 283236 46872
rect 283196 45552 283248 45558
rect 283196 45494 283248 45500
rect 282920 35964 282972 35970
rect 282920 35906 282972 35912
rect 282932 31634 282960 35906
rect 282932 31606 283052 31634
rect 281724 28960 281776 28966
rect 281724 28902 281776 28908
rect 281724 19372 281776 19378
rect 281724 19314 281776 19320
rect 281736 16046 281764 19314
rect 281724 16040 281776 16046
rect 281724 15982 281776 15988
rect 283024 10606 283052 31606
rect 283104 29232 283156 29238
rect 283102 29200 283104 29209
rect 283156 29200 283158 29209
rect 283102 29135 283158 29144
rect 283012 10600 283064 10606
rect 283012 10542 283064 10548
rect 281540 10464 281592 10470
rect 281540 10406 281592 10412
rect 280160 10396 280212 10402
rect 280160 10338 280212 10344
rect 283576 8106 283604 337622
rect 283656 337272 283708 337278
rect 283656 337214 283708 337220
rect 283484 8078 283604 8106
rect 281264 7472 281316 7478
rect 281264 7414 281316 7420
rect 280068 3392 280120 3398
rect 280068 3334 280120 3340
rect 279988 3046 280108 3074
rect 280080 480 280108 3046
rect 281276 480 281304 7414
rect 283484 4010 283512 8078
rect 283668 7970 283696 337214
rect 284404 16114 284432 340054
rect 285048 337550 285076 340068
rect 285036 337544 285088 337550
rect 285036 337486 285088 337492
rect 284944 337340 284996 337346
rect 284944 337282 284996 337288
rect 284392 16108 284444 16114
rect 284392 16050 284444 16056
rect 283576 7942 283696 7970
rect 283576 4554 283604 7942
rect 284760 7404 284812 7410
rect 284760 7346 284812 7352
rect 283656 6248 283708 6254
rect 283656 6190 283708 6196
rect 283564 4548 283616 4554
rect 283564 4490 283616 4496
rect 283472 4004 283524 4010
rect 283472 3946 283524 3952
rect 282460 3392 282512 3398
rect 282460 3334 282512 3340
rect 282472 480 282500 3334
rect 283668 480 283696 6190
rect 284772 480 284800 7346
rect 284956 4486 284984 337282
rect 285692 10538 285720 340068
rect 285784 340054 286350 340082
rect 285784 16182 285812 340054
rect 286888 337074 286916 340068
rect 287072 340054 287546 340082
rect 287716 340054 288190 340082
rect 286968 337544 287020 337550
rect 286968 337486 287020 337492
rect 286876 337068 286928 337074
rect 286876 337010 286928 337016
rect 285772 16176 285824 16182
rect 285772 16118 285824 16124
rect 285680 10532 285732 10538
rect 285680 10474 285732 10480
rect 284944 4480 284996 4486
rect 284944 4422 284996 4428
rect 286980 3194 287008 337486
rect 287072 10674 287100 340054
rect 287716 337906 287744 340054
rect 287256 337878 287744 337906
rect 288728 337890 288756 340068
rect 288716 337884 288768 337890
rect 287256 323626 287284 337878
rect 288716 337826 288768 337832
rect 287704 337748 287756 337754
rect 287704 337690 287756 337696
rect 287164 323598 287284 323626
rect 287164 307902 287192 323598
rect 287152 307896 287204 307902
rect 287152 307838 287204 307844
rect 287336 307896 287388 307902
rect 287336 307838 287388 307844
rect 287348 307766 287376 307838
rect 287336 307760 287388 307766
rect 287336 307702 287388 307708
rect 287244 298172 287296 298178
rect 287244 298114 287296 298120
rect 287256 278769 287284 298114
rect 287242 278760 287298 278769
rect 287242 278695 287298 278704
rect 287426 278760 287482 278769
rect 287426 278695 287482 278704
rect 287440 269142 287468 278695
rect 287244 269136 287296 269142
rect 287244 269078 287296 269084
rect 287428 269136 287480 269142
rect 287428 269078 287480 269084
rect 287256 259457 287284 269078
rect 287242 259448 287298 259457
rect 287242 259383 287298 259392
rect 287334 259312 287390 259321
rect 287334 259247 287390 259256
rect 287348 249898 287376 259247
rect 287152 249892 287204 249898
rect 287152 249834 287204 249840
rect 287336 249892 287388 249898
rect 287336 249834 287388 249840
rect 287164 249801 287192 249834
rect 287150 249792 287206 249801
rect 287150 249727 287206 249736
rect 287426 249792 287482 249801
rect 287426 249727 287482 249736
rect 287440 240174 287468 249727
rect 287244 240168 287296 240174
rect 287244 240110 287296 240116
rect 287428 240168 287480 240174
rect 287428 240110 287480 240116
rect 287256 220726 287284 240110
rect 287244 220720 287296 220726
rect 287244 220662 287296 220668
rect 287336 220720 287388 220726
rect 287336 220662 287388 220668
rect 287348 211313 287376 220662
rect 287334 211304 287390 211313
rect 287334 211239 287390 211248
rect 287242 211168 287298 211177
rect 287242 211103 287298 211112
rect 287256 206258 287284 211103
rect 287164 206230 287284 206258
rect 287164 201521 287192 206230
rect 287150 201512 287206 201521
rect 287150 201447 287206 201456
rect 287334 201512 287390 201521
rect 287334 201447 287336 201456
rect 287388 201447 287390 201456
rect 287336 201418 287388 201424
rect 287428 201408 287480 201414
rect 287428 201350 287480 201356
rect 287440 183598 287468 201350
rect 287244 183592 287296 183598
rect 287244 183534 287296 183540
rect 287428 183592 287480 183598
rect 287428 183534 287480 183540
rect 287256 182170 287284 183534
rect 287244 182164 287296 182170
rect 287244 182106 287296 182112
rect 287428 182164 287480 182170
rect 287428 182106 287480 182112
rect 287440 172553 287468 182106
rect 287242 172544 287298 172553
rect 287242 172479 287298 172488
rect 287426 172544 287482 172553
rect 287426 172479 287482 172488
rect 287256 145081 287284 172479
rect 287242 145072 287298 145081
rect 287242 145007 287298 145016
rect 287242 144936 287298 144945
rect 287242 144871 287298 144880
rect 287256 143546 287284 144871
rect 287244 143540 287296 143546
rect 287244 143482 287296 143488
rect 287244 133952 287296 133958
rect 287244 133894 287296 133900
rect 287256 125769 287284 133894
rect 287242 125760 287298 125769
rect 287242 125695 287298 125704
rect 287242 125624 287298 125633
rect 287242 125559 287298 125568
rect 287256 124166 287284 125559
rect 287244 124160 287296 124166
rect 287244 124102 287296 124108
rect 287152 114572 287204 114578
rect 287152 114514 287204 114520
rect 287164 106162 287192 114514
rect 287164 106134 287284 106162
rect 287256 104802 287284 106134
rect 287256 104774 287376 104802
rect 287348 95282 287376 104774
rect 287256 95254 287376 95282
rect 287256 95198 287284 95254
rect 287244 95192 287296 95198
rect 287244 95134 287296 95140
rect 287152 85672 287204 85678
rect 287152 85614 287204 85620
rect 287164 85542 287192 85614
rect 287152 85536 287204 85542
rect 287152 85478 287204 85484
rect 287244 75948 287296 75954
rect 287244 75890 287296 75896
rect 287256 66366 287284 75890
rect 287244 66360 287296 66366
rect 287244 66302 287296 66308
rect 287244 56704 287296 56710
rect 287244 56646 287296 56652
rect 287256 56574 287284 56646
rect 287244 56568 287296 56574
rect 287244 56510 287296 56516
rect 287244 47048 287296 47054
rect 287244 46990 287296 46996
rect 287256 46900 287284 46990
rect 287256 46872 287376 46900
rect 287348 37330 287376 46872
rect 287244 37324 287296 37330
rect 287244 37266 287296 37272
rect 287336 37324 287388 37330
rect 287336 37266 287388 37272
rect 287256 37210 287284 37266
rect 287164 37182 287284 37210
rect 287164 31634 287192 37182
rect 287164 31606 287284 31634
rect 287256 16250 287284 31606
rect 287244 16244 287296 16250
rect 287244 16186 287296 16192
rect 287060 10668 287112 10674
rect 287060 10610 287112 10616
rect 287612 10532 287664 10538
rect 287612 10474 287664 10480
rect 287152 6316 287204 6322
rect 287152 6258 287204 6264
rect 285956 3188 286008 3194
rect 285956 3130 286008 3136
rect 286968 3188 287020 3194
rect 286968 3130 287020 3136
rect 285968 480 285996 3130
rect 287164 480 287192 6258
rect 287624 3534 287652 10474
rect 287716 3738 287744 337690
rect 288820 335594 288848 340190
rect 290016 337618 290044 340068
rect 290004 337612 290056 337618
rect 290004 337554 290056 337560
rect 290568 337006 290596 340068
rect 290556 337000 290608 337006
rect 290556 336942 290608 336948
rect 288544 335566 288848 335594
rect 288544 321314 288572 335566
rect 288544 321286 288664 321314
rect 288636 318782 288664 321286
rect 288624 318776 288676 318782
rect 288624 318718 288676 318724
rect 288624 309188 288676 309194
rect 288624 309130 288676 309136
rect 288636 299470 288664 309130
rect 288624 299464 288676 299470
rect 288624 299406 288676 299412
rect 288624 289876 288676 289882
rect 288624 289818 288676 289824
rect 288636 280158 288664 289818
rect 288624 280152 288676 280158
rect 288624 280094 288676 280100
rect 288624 270564 288676 270570
rect 288624 270506 288676 270512
rect 288636 260846 288664 270506
rect 288624 260840 288676 260846
rect 288624 260782 288676 260788
rect 288624 251252 288676 251258
rect 288624 251194 288676 251200
rect 288636 234682 288664 251194
rect 288544 234654 288664 234682
rect 288544 234546 288572 234654
rect 288544 234518 288664 234546
rect 288636 222193 288664 234518
rect 288438 222184 288494 222193
rect 288438 222119 288494 222128
rect 288622 222184 288678 222193
rect 288622 222119 288678 222128
rect 288452 212566 288480 222119
rect 288440 212560 288492 212566
rect 288440 212502 288492 212508
rect 288624 212560 288676 212566
rect 288624 212502 288676 212508
rect 288636 202881 288664 212502
rect 289818 204776 289874 204785
rect 289818 204711 289874 204720
rect 289832 204513 289860 204711
rect 289818 204504 289874 204513
rect 289818 204439 289874 204448
rect 288438 202872 288494 202881
rect 288438 202807 288494 202816
rect 288622 202872 288678 202881
rect 288622 202807 288678 202816
rect 288452 193254 288480 202807
rect 288440 193248 288492 193254
rect 288440 193190 288492 193196
rect 288624 193248 288676 193254
rect 288624 193190 288676 193196
rect 288636 183569 288664 193190
rect 288438 183560 288494 183569
rect 288438 183495 288494 183504
rect 288622 183560 288678 183569
rect 288622 183495 288678 183504
rect 288452 173942 288480 183495
rect 288440 173936 288492 173942
rect 288440 173878 288492 173884
rect 288624 173936 288676 173942
rect 288624 173878 288676 173884
rect 288348 170128 288400 170134
rect 288346 170096 288348 170105
rect 288400 170096 288402 170105
rect 288346 170031 288402 170040
rect 288636 157434 288664 173878
rect 288544 157406 288664 157434
rect 288544 157162 288572 157406
rect 288544 157134 288664 157162
rect 288636 138122 288664 157134
rect 288544 138094 288664 138122
rect 288544 137986 288572 138094
rect 288544 137958 288664 137986
rect 288636 125769 288664 137958
rect 288622 125760 288678 125769
rect 288622 125695 288678 125704
rect 288622 125624 288678 125633
rect 288622 125559 288678 125568
rect 288636 118810 288664 125559
rect 288636 118782 288756 118810
rect 288728 118538 288756 118782
rect 288636 118510 288756 118538
rect 288636 99414 288664 118510
rect 288624 99408 288676 99414
rect 288624 99350 288676 99356
rect 288624 96688 288676 96694
rect 288624 96630 288676 96636
rect 288636 86970 288664 96630
rect 288624 86964 288676 86970
rect 288624 86906 288676 86912
rect 288624 77308 288676 77314
rect 288624 77250 288676 77256
rect 288636 47002 288664 77250
rect 290556 76016 290608 76022
rect 290556 75958 290608 75964
rect 290568 75857 290596 75958
rect 290554 75848 290610 75857
rect 290554 75783 290610 75792
rect 288544 46974 288664 47002
rect 288544 46918 288572 46974
rect 288532 46912 288584 46918
rect 288532 46854 288584 46860
rect 288624 46912 288676 46918
rect 288624 46854 288676 46860
rect 288636 28966 288664 46854
rect 288440 28960 288492 28966
rect 288440 28902 288492 28908
rect 288624 28960 288676 28966
rect 288624 28902 288676 28908
rect 288452 19394 288480 28902
rect 288452 19366 288572 19394
rect 288544 19310 288572 19366
rect 288532 19304 288584 19310
rect 288532 19246 288584 19252
rect 291212 10810 291240 340068
rect 291304 340054 291870 340082
rect 291304 16318 291332 340054
rect 292408 337822 292436 340068
rect 292592 340054 293066 340082
rect 293236 340054 293710 340082
rect 292396 337816 292448 337822
rect 292396 337758 292448 337764
rect 291292 16312 291344 16318
rect 291292 16254 291344 16260
rect 292592 10878 292620 340054
rect 293236 327321 293264 340054
rect 293868 337612 293920 337618
rect 293868 337554 293920 337560
rect 293222 327312 293278 327321
rect 293222 327247 293278 327256
rect 292762 327176 292818 327185
rect 292762 327111 292818 327120
rect 292776 327078 292804 327111
rect 292764 327072 292816 327078
rect 292764 327014 292816 327020
rect 292764 317484 292816 317490
rect 292764 317426 292816 317432
rect 292776 298110 292804 317426
rect 292764 298104 292816 298110
rect 292764 298046 292816 298052
rect 292672 288448 292724 288454
rect 292672 288390 292724 288396
rect 292684 280226 292712 288390
rect 292672 280220 292724 280226
rect 292672 280162 292724 280168
rect 292764 280220 292816 280226
rect 292764 280162 292816 280168
rect 292776 274258 292804 280162
rect 292776 274230 292988 274258
rect 292960 269249 292988 274230
rect 292670 269240 292726 269249
rect 292670 269175 292726 269184
rect 292946 269240 293002 269249
rect 292946 269175 293002 269184
rect 292684 269074 292712 269175
rect 292672 269068 292724 269074
rect 292672 269010 292724 269016
rect 292764 260772 292816 260778
rect 292764 260714 292816 260720
rect 292776 251190 292804 260714
rect 292764 251184 292816 251190
rect 292764 251126 292816 251132
rect 292764 240168 292816 240174
rect 292764 240110 292816 240116
rect 292776 240038 292804 240110
rect 292764 240032 292816 240038
rect 292764 239974 292816 239980
rect 292764 230512 292816 230518
rect 292764 230454 292816 230460
rect 292776 220930 292804 230454
rect 292764 220924 292816 220930
rect 292764 220866 292816 220872
rect 292672 220856 292724 220862
rect 292672 220798 292724 220804
rect 292684 211206 292712 220798
rect 292672 211200 292724 211206
rect 292672 211142 292724 211148
rect 292764 211200 292816 211206
rect 292764 211142 292816 211148
rect 292776 205698 292804 211142
rect 292764 205692 292816 205698
rect 292764 205634 292816 205640
rect 292856 205556 292908 205562
rect 292856 205498 292908 205504
rect 292868 198098 292896 205498
rect 292868 198070 292988 198098
rect 292960 193254 292988 198070
rect 292764 193248 292816 193254
rect 292762 193216 292764 193225
rect 292948 193248 293000 193254
rect 292816 193216 292818 193225
rect 292762 193151 292818 193160
rect 292946 193216 292948 193225
rect 293000 193216 293002 193225
rect 292946 193151 293002 193160
rect 292960 182170 292988 193151
rect 292856 182164 292908 182170
rect 292856 182106 292908 182112
rect 292948 182164 293000 182170
rect 292948 182106 293000 182112
rect 292868 172530 292896 182106
rect 292776 172514 292896 172530
rect 292764 172508 292896 172514
rect 292816 172502 292896 172508
rect 292764 172450 292816 172456
rect 292776 172419 292804 172450
rect 292764 164212 292816 164218
rect 292764 164154 292816 164160
rect 292776 162874 292804 164154
rect 292776 162846 292896 162874
rect 292868 155922 292896 162846
rect 292856 155916 292908 155922
rect 292856 155858 292908 155864
rect 292764 147620 292816 147626
rect 292764 147562 292816 147568
rect 292776 144906 292804 147562
rect 292764 144900 292816 144906
rect 292764 144842 292816 144848
rect 292764 135312 292816 135318
rect 292764 135254 292816 135260
rect 292776 133890 292804 135254
rect 292764 133884 292816 133890
rect 292764 133826 292816 133832
rect 292764 125588 292816 125594
rect 292764 125530 292816 125536
rect 292776 124250 292804 125530
rect 292776 124222 292896 124250
rect 292868 124166 292896 124222
rect 292856 124160 292908 124166
rect 292856 124102 292908 124108
rect 292948 113212 293000 113218
rect 292948 113154 293000 113160
rect 292960 104922 292988 113154
rect 292764 104916 292816 104922
rect 292764 104858 292816 104864
rect 292948 104916 293000 104922
rect 292948 104858 293000 104864
rect 292776 98818 292804 104858
rect 292776 98790 292896 98818
rect 292868 77466 292896 98790
rect 292776 77438 292896 77466
rect 292776 77194 292804 77438
rect 292776 77166 292896 77194
rect 292868 67658 292896 77166
rect 292764 67652 292816 67658
rect 292764 67594 292816 67600
rect 292856 67652 292908 67658
rect 292856 67594 292908 67600
rect 292776 66230 292804 67594
rect 292764 66224 292816 66230
rect 292764 66166 292816 66172
rect 292856 47048 292908 47054
rect 292856 46990 292908 46996
rect 292868 45558 292896 46990
rect 292856 45552 292908 45558
rect 292856 45494 292908 45500
rect 292856 35964 292908 35970
rect 292856 35906 292908 35912
rect 292868 30546 292896 35906
rect 292776 30518 292896 30546
rect 292776 16386 292804 30518
rect 293222 29336 293278 29345
rect 293222 29271 293278 29280
rect 293236 28937 293264 29271
rect 293222 28928 293278 28937
rect 293222 28863 293278 28872
rect 292764 16380 292816 16386
rect 292764 16322 292816 16328
rect 292580 10872 292632 10878
rect 292580 10814 292632 10820
rect 291200 10804 291252 10810
rect 291200 10746 291252 10752
rect 289912 10668 289964 10674
rect 289912 10610 289964 10616
rect 289820 10600 289872 10606
rect 289820 10542 289872 10548
rect 287704 3732 287756 3738
rect 287704 3674 287756 3680
rect 289832 3670 289860 10542
rect 289820 3664 289872 3670
rect 289820 3606 289872 3612
rect 289544 3596 289596 3602
rect 289544 3538 289596 3544
rect 287612 3528 287664 3534
rect 287612 3470 287664 3476
rect 288348 3256 288400 3262
rect 288348 3198 288400 3204
rect 288360 480 288388 3198
rect 289556 480 289584 3538
rect 289924 3534 289952 10610
rect 292948 10328 293000 10334
rect 292948 10270 293000 10276
rect 290740 6384 290792 6390
rect 290740 6326 290792 6332
rect 289912 3528 289964 3534
rect 289912 3470 289964 3476
rect 290752 480 290780 6326
rect 291936 3664 291988 3670
rect 291936 3606 291988 3612
rect 291948 480 291976 3606
rect 292960 3262 292988 10270
rect 292948 3256 293000 3262
rect 292948 3198 293000 3204
rect 293880 3194 293908 337554
rect 294248 336938 294276 340068
rect 294236 336932 294288 336938
rect 294236 336874 294288 336880
rect 294524 335306 294552 340190
rect 295352 340054 295550 340082
rect 295812 340054 296102 340082
rect 294604 337816 294656 337822
rect 294604 337758 294656 337764
rect 294512 335300 294564 335306
rect 294512 335242 294564 335248
rect 294052 325712 294104 325718
rect 294142 325680 294198 325689
rect 294104 325660 294142 325666
rect 294052 325654 294142 325660
rect 294064 325638 294142 325654
rect 294142 325615 294198 325624
rect 294326 325680 294382 325689
rect 294326 325615 294382 325624
rect 294340 316062 294368 325615
rect 294144 316056 294196 316062
rect 294144 315998 294196 316004
rect 294328 316056 294380 316062
rect 294328 315998 294380 316004
rect 294156 311982 294184 315998
rect 294144 311976 294196 311982
rect 294144 311918 294196 311924
rect 294144 311840 294196 311846
rect 294144 311782 294196 311788
rect 294156 273222 294184 311782
rect 294144 273216 294196 273222
rect 294144 273158 294196 273164
rect 294144 273080 294196 273086
rect 294144 273022 294196 273028
rect 294156 260846 294184 273022
rect 294144 260840 294196 260846
rect 294144 260782 294196 260788
rect 294144 251252 294196 251258
rect 294144 251194 294196 251200
rect 294156 241505 294184 251194
rect 293958 241496 294014 241505
rect 293958 241431 294014 241440
rect 294142 241496 294198 241505
rect 294142 241431 294198 241440
rect 293972 231878 294000 241431
rect 293960 231872 294012 231878
rect 293960 231814 294012 231820
rect 294144 231872 294196 231878
rect 294144 231814 294196 231820
rect 294156 222193 294184 231814
rect 293958 222184 294014 222193
rect 293958 222119 294014 222128
rect 294142 222184 294198 222193
rect 294142 222119 294198 222128
rect 293972 218362 294000 222119
rect 293972 218334 294276 218362
rect 294248 211154 294276 218334
rect 294156 211126 294276 211154
rect 294156 200122 294184 211126
rect 294144 200116 294196 200122
rect 294144 200058 294196 200064
rect 294236 200116 294288 200122
rect 294236 200058 294288 200064
rect 294248 174010 294276 200058
rect 294236 174004 294288 174010
rect 294236 173946 294288 173952
rect 294144 173868 294196 173874
rect 294144 173810 294196 173816
rect 294156 168994 294184 173810
rect 294064 168966 294184 168994
rect 294064 157434 294092 168966
rect 293972 157406 294092 157434
rect 293972 157298 294000 157406
rect 293972 157270 294092 157298
rect 294064 144906 294092 157270
rect 294052 144900 294104 144906
rect 294052 144842 294104 144848
rect 294236 144900 294288 144906
rect 294236 144842 294288 144848
rect 294248 139890 294276 144842
rect 294156 139862 294276 139890
rect 294156 125769 294184 139862
rect 294142 125760 294198 125769
rect 294142 125695 294198 125704
rect 294050 125624 294106 125633
rect 294050 125559 294106 125568
rect 294064 114646 294092 125559
rect 294052 114640 294104 114646
rect 294052 114582 294104 114588
rect 294144 114572 294196 114578
rect 294144 114514 294196 114520
rect 294156 109750 294184 114514
rect 294144 109744 294196 109750
rect 294144 109686 294196 109692
rect 294144 109608 294196 109614
rect 294144 109550 294196 109556
rect 294156 98818 294184 109550
rect 294064 98790 294184 98818
rect 294064 93922 294092 98790
rect 294064 93894 294184 93922
rect 294156 93838 294184 93894
rect 294144 93832 294196 93838
rect 294144 93774 294196 93780
rect 294144 84244 294196 84250
rect 294144 84186 294196 84192
rect 294156 77364 294184 84186
rect 294156 77336 294276 77364
rect 294248 77194 294276 77336
rect 294064 77166 294276 77194
rect 294064 72486 294092 77166
rect 294052 72480 294104 72486
rect 294052 72422 294104 72428
rect 294236 72480 294288 72486
rect 294236 72422 294288 72428
rect 294248 66230 294276 72422
rect 293960 66224 294012 66230
rect 293960 66166 294012 66172
rect 294236 66224 294288 66230
rect 294236 66166 294288 66172
rect 293972 51762 294000 66166
rect 293972 51734 294092 51762
rect 294064 42106 294092 51734
rect 294064 42078 294276 42106
rect 294248 41290 294276 42078
rect 294156 41262 294276 41290
rect 294156 28966 294184 41262
rect 293960 28960 294012 28966
rect 293960 28902 294012 28908
rect 294144 28960 294196 28966
rect 294144 28902 294196 28908
rect 293972 12510 294000 28902
rect 293960 12504 294012 12510
rect 293960 12446 294012 12452
rect 294328 5296 294380 5302
rect 294328 5238 294380 5244
rect 293132 3188 293184 3194
rect 293132 3130 293184 3136
rect 293868 3188 293920 3194
rect 293868 3130 293920 3136
rect 293144 480 293172 3130
rect 294340 480 294368 5238
rect 294616 3398 294644 337758
rect 295246 134192 295302 134201
rect 295246 134127 295302 134136
rect 295260 133657 295288 134127
rect 295246 133648 295302 133657
rect 295246 133583 295302 133592
rect 295352 11830 295380 340054
rect 295812 331294 295840 340054
rect 295800 331288 295852 331294
rect 295800 331230 295852 331236
rect 295616 331220 295668 331226
rect 295616 331162 295668 331168
rect 295628 311930 295656 331162
rect 295536 311902 295656 311930
rect 295536 307766 295564 311902
rect 295524 307760 295576 307766
rect 295524 307702 295576 307708
rect 295708 293276 295760 293282
rect 295708 293218 295760 293224
rect 295720 280158 295748 293218
rect 295432 280152 295484 280158
rect 295432 280094 295484 280100
rect 295708 280152 295760 280158
rect 295708 280094 295760 280100
rect 295444 273970 295472 280094
rect 295432 273964 295484 273970
rect 295432 273906 295484 273912
rect 295616 263492 295668 263498
rect 295616 263434 295668 263440
rect 295628 260846 295656 263434
rect 295616 260840 295668 260846
rect 295616 260782 295668 260788
rect 295524 251252 295576 251258
rect 295524 251194 295576 251200
rect 295536 246378 295564 251194
rect 295536 246350 295748 246378
rect 295720 241534 295748 246350
rect 295708 241528 295760 241534
rect 295708 241470 295760 241476
rect 295800 241528 295852 241534
rect 295800 241470 295852 241476
rect 295812 231878 295840 241470
rect 295524 231872 295576 231878
rect 295524 231814 295576 231820
rect 295800 231872 295852 231878
rect 295800 231814 295852 231820
rect 295536 222222 295564 231814
rect 295524 222216 295576 222222
rect 295524 222158 295576 222164
rect 295800 222216 295852 222222
rect 295800 222158 295852 222164
rect 295812 216050 295840 222158
rect 295536 216022 295840 216050
rect 295536 209778 295564 216022
rect 295524 209772 295576 209778
rect 295524 209714 295576 209720
rect 295524 202836 295576 202842
rect 295524 202778 295576 202784
rect 295536 200122 295564 202778
rect 295524 200116 295576 200122
rect 295524 200058 295576 200064
rect 295708 183524 295760 183530
rect 295708 183466 295760 183472
rect 295720 172582 295748 183466
rect 295616 172576 295668 172582
rect 295616 172518 295668 172524
rect 295708 172576 295760 172582
rect 295708 172518 295760 172524
rect 295628 157434 295656 172518
rect 296628 170128 296680 170134
rect 296626 170096 296628 170105
rect 296680 170096 296682 170105
rect 296626 170031 296682 170040
rect 295628 157406 295748 157434
rect 295720 153218 295748 157406
rect 295628 153190 295748 153218
rect 295628 144906 295656 153190
rect 295616 144900 295668 144906
rect 295616 144842 295668 144848
rect 295708 144900 295760 144906
rect 295708 144842 295760 144848
rect 295720 135289 295748 144842
rect 295522 135280 295578 135289
rect 295522 135215 295578 135224
rect 295706 135280 295762 135289
rect 295706 135215 295762 135224
rect 295536 129010 295564 135215
rect 295444 128982 295564 129010
rect 295444 125338 295472 128982
rect 295444 125310 295656 125338
rect 295628 124166 295656 125310
rect 295524 124160 295576 124166
rect 295524 124102 295576 124108
rect 295616 124160 295668 124166
rect 295616 124102 295668 124108
rect 295536 113506 295564 124102
rect 295536 113478 295656 113506
rect 295628 113234 295656 113478
rect 295536 113206 295656 113234
rect 295536 113150 295564 113206
rect 295524 113144 295576 113150
rect 295524 113086 295576 113092
rect 295524 103556 295576 103562
rect 295524 103498 295576 103504
rect 295536 95266 295564 103498
rect 295524 95260 295576 95266
rect 295524 95202 295576 95208
rect 295616 95124 295668 95130
rect 295616 95066 295668 95072
rect 295628 85610 295656 95066
rect 295524 85604 295576 85610
rect 295524 85546 295576 85552
rect 295616 85604 295668 85610
rect 295616 85546 295668 85552
rect 295536 56522 295564 85546
rect 295536 56494 295748 56522
rect 295720 37330 295748 56494
rect 295524 37324 295576 37330
rect 295524 37266 295576 37272
rect 295708 37324 295760 37330
rect 295708 37266 295760 37272
rect 295536 15162 295564 37266
rect 295524 15156 295576 15162
rect 295524 15098 295576 15104
rect 295340 11824 295392 11830
rect 295340 11766 295392 11772
rect 296732 5370 296760 340068
rect 296916 340054 297390 340082
rect 297560 340054 297942 340082
rect 298112 340054 298586 340082
rect 298756 340054 299230 340082
rect 299584 340054 299782 340082
rect 300136 340054 300426 340082
rect 300872 340054 300978 340082
rect 301056 340054 301622 340082
rect 302266 340054 302464 340082
rect 296812 334484 296864 334490
rect 296812 334426 296864 334432
rect 296824 8974 296852 334426
rect 296916 13190 296944 340054
rect 297560 334490 297588 340054
rect 297548 334484 297600 334490
rect 297548 334426 297600 334432
rect 298006 170096 298062 170105
rect 298006 170031 298062 170040
rect 298020 169833 298048 170031
rect 298006 169824 298062 169833
rect 298006 169759 298062 169768
rect 298006 134192 298062 134201
rect 298006 134127 298008 134136
rect 298060 134127 298062 134136
rect 298008 134098 298060 134104
rect 298006 110800 298062 110809
rect 298006 110735 298062 110744
rect 298020 110537 298048 110735
rect 298006 110528 298062 110537
rect 298006 110463 298062 110472
rect 296904 13184 296956 13190
rect 296904 13126 296956 13132
rect 296812 8968 296864 8974
rect 296812 8910 296864 8916
rect 298112 5438 298140 340054
rect 298756 331242 298784 340054
rect 299480 333940 299532 333946
rect 299480 333882 299532 333888
rect 298388 331214 298784 331242
rect 298388 311930 298416 331214
rect 298296 311902 298416 311930
rect 298296 302326 298324 311902
rect 298284 302320 298336 302326
rect 298284 302262 298336 302268
rect 298376 302116 298428 302122
rect 298376 302058 298428 302064
rect 298388 296682 298416 302058
rect 298376 296676 298428 296682
rect 298376 296618 298428 296624
rect 298468 287088 298520 287094
rect 298468 287030 298520 287036
rect 298480 280158 298508 287030
rect 298468 280152 298520 280158
rect 298468 280094 298520 280100
rect 298284 280084 298336 280090
rect 298284 280026 298336 280032
rect 298296 278769 298324 280026
rect 298282 278760 298338 278769
rect 298282 278695 298338 278704
rect 298558 278760 298614 278769
rect 298558 278695 298614 278704
rect 298572 253858 298600 278695
rect 298296 253830 298600 253858
rect 298296 251190 298324 253830
rect 298284 251184 298336 251190
rect 298284 251126 298336 251132
rect 298560 251184 298612 251190
rect 298560 251126 298612 251132
rect 298572 231878 298600 251126
rect 298284 231872 298336 231878
rect 298284 231814 298336 231820
rect 298560 231872 298612 231878
rect 298560 231814 298612 231820
rect 298296 222222 298324 231814
rect 298284 222216 298336 222222
rect 298284 222158 298336 222164
rect 298560 222216 298612 222222
rect 298560 222158 298612 222164
rect 298572 212566 298600 222158
rect 298284 212560 298336 212566
rect 298284 212502 298336 212508
rect 298560 212560 298612 212566
rect 298560 212502 298612 212508
rect 298296 205698 298324 212502
rect 298284 205692 298336 205698
rect 298284 205634 298336 205640
rect 298376 205624 298428 205630
rect 298376 205566 298428 205572
rect 298388 198098 298416 205566
rect 298388 198070 298508 198098
rect 298480 193254 298508 198070
rect 298284 193248 298336 193254
rect 298284 193190 298336 193196
rect 298468 193248 298520 193254
rect 298468 193190 298520 193196
rect 298296 186454 298324 193190
rect 298284 186448 298336 186454
rect 298284 186390 298336 186396
rect 298284 183592 298336 183598
rect 298284 183534 298336 183540
rect 298296 182170 298324 183534
rect 298284 182164 298336 182170
rect 298284 182106 298336 182112
rect 298468 182164 298520 182170
rect 298468 182106 298520 182112
rect 298480 172553 298508 182106
rect 298190 172544 298246 172553
rect 298190 172479 298246 172488
rect 298466 172544 298522 172553
rect 298466 172479 298522 172488
rect 298204 164286 298232 172479
rect 299388 169720 299440 169726
rect 299386 169688 299388 169697
rect 299440 169688 299442 169697
rect 299386 169623 299442 169632
rect 298192 164280 298244 164286
rect 298192 164222 298244 164228
rect 298284 164280 298336 164286
rect 298284 164222 298336 164228
rect 298296 162858 298324 164222
rect 298284 162852 298336 162858
rect 298284 162794 298336 162800
rect 298284 157344 298336 157350
rect 298284 157286 298336 157292
rect 298296 153218 298324 157286
rect 298296 153190 298416 153218
rect 298388 149818 298416 153190
rect 298388 149790 298508 149818
rect 298480 144945 298508 149790
rect 298282 144936 298338 144945
rect 298282 144871 298284 144880
rect 298336 144871 298338 144880
rect 298466 144936 298522 144945
rect 298466 144871 298468 144880
rect 298284 144842 298336 144848
rect 298520 144871 298522 144880
rect 298468 144842 298520 144848
rect 298480 139890 298508 144842
rect 298388 139862 298508 139890
rect 298388 124250 298416 139862
rect 298296 124222 298416 124250
rect 298296 118794 298324 124222
rect 298284 118788 298336 118794
rect 298284 118730 298336 118736
rect 298376 102196 298428 102202
rect 298376 102138 298428 102144
rect 298388 99482 298416 102138
rect 298376 99476 298428 99482
rect 298376 99418 298428 99424
rect 298376 93832 298428 93838
rect 298376 93774 298428 93780
rect 298388 89010 298416 93774
rect 298376 89004 298428 89010
rect 298376 88946 298428 88952
rect 298560 84244 298612 84250
rect 298560 84186 298612 84192
rect 298572 75993 298600 84186
rect 298282 75984 298338 75993
rect 298282 75919 298338 75928
rect 298558 75984 298614 75993
rect 298558 75919 298614 75928
rect 298296 58002 298324 75919
rect 298284 57996 298336 58002
rect 298284 57938 298336 57944
rect 298376 57860 298428 57866
rect 298376 57802 298428 57808
rect 298388 55214 298416 57802
rect 298376 55208 298428 55214
rect 298376 55150 298428 55156
rect 298468 55208 298520 55214
rect 298468 55150 298520 55156
rect 298480 12186 298508 55150
rect 298204 12158 298508 12186
rect 298204 9602 298232 12158
rect 298204 9574 298324 9602
rect 298296 7585 298324 9574
rect 298282 7576 298338 7585
rect 298282 7511 298338 7520
rect 299492 5506 299520 333882
rect 299584 8945 299612 340054
rect 300136 333946 300164 340054
rect 300124 333940 300176 333946
rect 300124 333882 300176 333888
rect 299664 10464 299716 10470
rect 299664 10406 299716 10412
rect 299570 8936 299626 8945
rect 299570 8871 299626 8880
rect 299480 5500 299532 5506
rect 299480 5442 299532 5448
rect 298100 5432 298152 5438
rect 298100 5374 298152 5380
rect 296720 5364 296772 5370
rect 296720 5306 296772 5312
rect 297916 5364 297968 5370
rect 297916 5306 297968 5312
rect 296720 3596 296772 3602
rect 296720 3538 296772 3544
rect 294604 3392 294656 3398
rect 294604 3334 294656 3340
rect 295524 3392 295576 3398
rect 295524 3334 295576 3340
rect 295536 480 295564 3334
rect 296732 480 296760 3538
rect 297928 480 297956 5306
rect 299112 3732 299164 3738
rect 299112 3674 299164 3680
rect 299124 480 299152 3674
rect 299676 3670 299704 10406
rect 300872 7342 300900 340054
rect 300950 204776 301006 204785
rect 300950 204711 301006 204720
rect 300964 204377 300992 204711
rect 300950 204368 301006 204377
rect 300950 204303 301006 204312
rect 301056 10946 301084 340054
rect 302332 335640 302384 335646
rect 302332 335582 302384 335588
rect 301594 134192 301650 134201
rect 301594 134127 301596 134136
rect 301648 134127 301650 134136
rect 301596 134098 301648 134104
rect 302344 11014 302372 335582
rect 302436 11966 302464 340054
rect 302528 340054 302818 340082
rect 303080 340054 303462 340082
rect 303724 340054 304106 340082
rect 304368 340054 304658 340082
rect 305012 340054 305302 340082
rect 305380 340054 305946 340082
rect 302424 11960 302476 11966
rect 302424 11902 302476 11908
rect 302332 11008 302384 11014
rect 302332 10950 302384 10956
rect 301044 10940 301096 10946
rect 301044 10882 301096 10888
rect 300952 10396 301004 10402
rect 300952 10338 301004 10344
rect 300860 7336 300912 7342
rect 300860 7278 300912 7284
rect 300308 4004 300360 4010
rect 300308 3946 300360 3952
rect 299664 3664 299716 3670
rect 299664 3606 299716 3612
rect 300320 480 300348 3946
rect 300964 3738 300992 10338
rect 302528 7274 302556 340054
rect 303080 335646 303108 340054
rect 303068 335640 303120 335646
rect 303068 335582 303120 335588
rect 303620 335640 303672 335646
rect 303620 335582 303672 335588
rect 302976 169720 303028 169726
rect 302974 169688 302976 169697
rect 303028 169688 303030 169697
rect 302974 169623 303030 169632
rect 303632 13326 303660 335582
rect 303620 13320 303672 13326
rect 303620 13262 303672 13268
rect 303724 13258 303752 340054
rect 304368 335646 304396 340054
rect 304356 335640 304408 335646
rect 304356 335582 304408 335588
rect 304908 124228 304960 124234
rect 304908 124170 304960 124176
rect 304920 115977 304948 124170
rect 304906 115968 304962 115977
rect 304906 115903 304962 115912
rect 304262 64152 304318 64161
rect 304262 64087 304318 64096
rect 304276 63617 304304 64087
rect 304262 63608 304318 63617
rect 304262 63543 304318 63552
rect 303712 13252 303764 13258
rect 303712 13194 303764 13200
rect 305012 10266 305040 340054
rect 305380 335594 305408 340054
rect 305196 335566 305408 335594
rect 305196 331226 305224 335566
rect 306380 331968 306432 331974
rect 306380 331910 306432 331916
rect 305184 331220 305236 331226
rect 305184 331162 305236 331168
rect 305276 331152 305328 331158
rect 305276 331094 305328 331100
rect 305288 309194 305316 331094
rect 305184 309188 305236 309194
rect 305184 309130 305236 309136
rect 305276 309188 305328 309194
rect 305276 309130 305328 309136
rect 305196 299470 305224 309130
rect 305184 299464 305236 299470
rect 305184 299406 305236 299412
rect 305184 289876 305236 289882
rect 305184 289818 305236 289824
rect 305196 280158 305224 289818
rect 305184 280152 305236 280158
rect 305184 280094 305236 280100
rect 305184 270564 305236 270570
rect 305184 270506 305236 270512
rect 305196 260846 305224 270506
rect 305184 260840 305236 260846
rect 305184 260782 305236 260788
rect 305184 251252 305236 251258
rect 305184 251194 305236 251200
rect 305196 241505 305224 251194
rect 305182 241496 305238 241505
rect 305182 241431 305238 241440
rect 305366 241496 305422 241505
rect 305366 241431 305422 241440
rect 305380 231878 305408 241431
rect 305184 231872 305236 231878
rect 305184 231814 305236 231820
rect 305368 231872 305420 231878
rect 305368 231814 305420 231820
rect 305196 222193 305224 231814
rect 305182 222184 305238 222193
rect 305182 222119 305238 222128
rect 305366 222184 305422 222193
rect 305366 222119 305422 222128
rect 305380 212566 305408 222119
rect 305184 212560 305236 212566
rect 305184 212502 305236 212508
rect 305368 212560 305420 212566
rect 305368 212502 305420 212508
rect 305196 202881 305224 212502
rect 305182 202872 305238 202881
rect 305182 202807 305238 202816
rect 305366 202872 305422 202881
rect 305366 202807 305422 202816
rect 305380 193254 305408 202807
rect 305184 193248 305236 193254
rect 305184 193190 305236 193196
rect 305368 193248 305420 193254
rect 305368 193190 305420 193196
rect 305196 167090 305224 193190
rect 305104 167062 305224 167090
rect 305104 166954 305132 167062
rect 305104 166926 305224 166954
rect 305196 154737 305224 166926
rect 305182 154728 305238 154737
rect 305182 154663 305238 154672
rect 305182 154592 305238 154601
rect 305182 154527 305238 154536
rect 305196 147778 305224 154527
rect 305196 147750 305316 147778
rect 305288 145081 305316 147750
rect 305274 145072 305330 145081
rect 305274 145007 305330 145016
rect 305090 144936 305146 144945
rect 305090 144871 305146 144880
rect 305104 143546 305132 144871
rect 305092 143540 305144 143546
rect 305092 143482 305144 143488
rect 305092 133952 305144 133958
rect 305092 133894 305144 133900
rect 305104 125730 305132 133894
rect 305092 125724 305144 125730
rect 305092 125666 305144 125672
rect 305090 115968 305146 115977
rect 305090 115903 305092 115912
rect 305144 115903 305146 115912
rect 305092 115874 305144 115880
rect 305184 106344 305236 106350
rect 305184 106287 305236 106292
rect 305182 106278 305238 106287
rect 305182 106213 305238 106222
rect 305274 106040 305330 106049
rect 305274 105975 305330 105984
rect 305288 99226 305316 105975
rect 305196 99198 305316 99226
rect 305196 86970 305224 99198
rect 305184 86964 305236 86970
rect 305184 86906 305236 86912
rect 305184 77308 305236 77314
rect 305184 77250 305236 77256
rect 305196 70514 305224 77250
rect 305184 70508 305236 70514
rect 305184 70450 305236 70456
rect 305184 67652 305236 67658
rect 305184 67594 305236 67600
rect 305196 51202 305224 67594
rect 305184 51196 305236 51202
rect 305184 51138 305236 51144
rect 305092 51060 305144 51066
rect 305092 51002 305144 51008
rect 305104 19310 305132 51002
rect 305092 19304 305144 19310
rect 305092 19246 305144 19252
rect 305000 10260 305052 10266
rect 305000 10202 305052 10208
rect 306392 10198 306420 331910
rect 306484 13530 306512 340068
rect 306760 340054 307142 340082
rect 307786 340054 307984 340082
rect 306760 331974 306788 340054
rect 307852 335640 307904 335646
rect 307852 335582 307904 335588
rect 306748 331968 306800 331974
rect 306748 331910 306800 331916
rect 307574 134056 307630 134065
rect 307758 134056 307814 134065
rect 307630 134014 307758 134042
rect 307574 133991 307630 134000
rect 307758 133991 307814 134000
rect 307864 13598 307892 335582
rect 307852 13592 307904 13598
rect 307852 13534 307904 13540
rect 306472 13524 306524 13530
rect 306472 13466 306524 13472
rect 307956 13394 307984 340054
rect 308048 340054 308338 340082
rect 308508 340054 308982 340082
rect 309152 340054 309626 340082
rect 309704 340054 310178 340082
rect 310532 340054 310822 340082
rect 311176 340054 311466 340082
rect 308048 335646 308076 340054
rect 308036 335640 308088 335646
rect 308036 335582 308088 335588
rect 308508 331242 308536 340054
rect 308048 331214 308536 331242
rect 308048 222193 308076 331214
rect 308034 222184 308090 222193
rect 308034 222119 308090 222128
rect 308310 222184 308366 222193
rect 308310 222119 308366 222128
rect 308324 212566 308352 222119
rect 308128 212560 308180 212566
rect 308128 212502 308180 212508
rect 308312 212560 308364 212566
rect 308312 212502 308364 212508
rect 308140 202881 308168 212502
rect 308126 202872 308182 202881
rect 308126 202807 308182 202816
rect 308310 202872 308366 202881
rect 308310 202807 308366 202816
rect 308324 193254 308352 202807
rect 308128 193248 308180 193254
rect 308128 193190 308180 193196
rect 308312 193248 308364 193254
rect 308312 193190 308364 193196
rect 308140 176610 308168 193190
rect 309046 181248 309102 181257
rect 309046 181183 309102 181192
rect 309060 180849 309088 181183
rect 309046 180840 309102 180849
rect 309046 180775 309102 180784
rect 308140 176582 308260 176610
rect 308232 173942 308260 176582
rect 308128 173936 308180 173942
rect 308128 173878 308180 173884
rect 308220 173936 308272 173942
rect 308220 173878 308272 173884
rect 308140 169130 308168 173878
rect 309048 169856 309100 169862
rect 309046 169824 309048 169833
rect 309100 169824 309102 169833
rect 309046 169759 309102 169768
rect 308048 169102 308168 169130
rect 308048 164218 308076 169102
rect 308036 164212 308088 164218
rect 308036 164154 308088 164160
rect 308220 164212 308272 164218
rect 308220 164154 308272 164160
rect 308232 162858 308260 164154
rect 308220 162852 308272 162858
rect 308220 162794 308272 162800
rect 308404 162852 308456 162858
rect 308404 162794 308456 162800
rect 308416 153241 308444 162794
rect 308218 153232 308274 153241
rect 308218 153167 308274 153176
rect 308402 153232 308458 153241
rect 308402 153167 308458 153176
rect 308232 144974 308260 153167
rect 308128 144968 308180 144974
rect 308128 144910 308180 144916
rect 308220 144968 308272 144974
rect 308220 144910 308272 144916
rect 308140 138122 308168 144910
rect 308048 138094 308168 138122
rect 308048 137986 308076 138094
rect 308048 137958 308168 137986
rect 308140 118726 308168 137958
rect 308128 118720 308180 118726
rect 308128 118662 308180 118668
rect 308128 118584 308180 118590
rect 308128 118526 308180 118532
rect 308140 99414 308168 118526
rect 308128 99408 308180 99414
rect 308128 99350 308180 99356
rect 308128 96688 308180 96694
rect 308128 96630 308180 96636
rect 308140 86970 308168 96630
rect 308128 86964 308180 86970
rect 308128 86906 308180 86912
rect 308128 77308 308180 77314
rect 308128 77250 308180 77256
rect 308140 58002 308168 77250
rect 309046 76256 309102 76265
rect 309046 76191 309048 76200
rect 309100 76191 309102 76200
rect 309048 76162 309100 76168
rect 308036 57996 308088 58002
rect 308036 57938 308088 57944
rect 308128 57996 308180 58002
rect 308128 57938 308180 57944
rect 308048 50946 308076 57938
rect 308048 50918 308168 50946
rect 308140 21978 308168 50918
rect 308048 21950 308168 21978
rect 308048 19310 308076 21950
rect 308036 19304 308088 19310
rect 308036 19246 308088 19252
rect 309152 13666 309180 340054
rect 309704 328506 309732 340054
rect 309784 337952 309836 337958
rect 309784 337894 309836 337900
rect 309416 328500 309468 328506
rect 309416 328442 309468 328448
rect 309692 328500 309744 328506
rect 309692 328442 309744 328448
rect 309428 311930 309456 328442
rect 309336 311902 309456 311930
rect 309336 309126 309364 311902
rect 309324 309120 309376 309126
rect 309324 309062 309376 309068
rect 309416 299532 309468 299538
rect 309416 299474 309468 299480
rect 309428 299441 309456 299474
rect 309414 299432 309470 299441
rect 309414 299367 309470 299376
rect 309598 299432 309654 299441
rect 309598 299367 309654 299376
rect 309612 289882 309640 299367
rect 309324 289876 309376 289882
rect 309324 289818 309376 289824
rect 309600 289876 309652 289882
rect 309600 289818 309652 289824
rect 309336 289746 309364 289818
rect 309324 289740 309376 289746
rect 309324 289682 309376 289688
rect 309416 280220 309468 280226
rect 309416 280162 309468 280168
rect 309428 280129 309456 280162
rect 309414 280120 309470 280129
rect 309414 280055 309470 280064
rect 309598 280120 309654 280129
rect 309598 280055 309654 280064
rect 309612 270570 309640 280055
rect 309324 270564 309376 270570
rect 309324 270506 309376 270512
rect 309600 270564 309652 270570
rect 309600 270506 309652 270512
rect 309336 270434 309364 270506
rect 309324 270428 309376 270434
rect 309324 270370 309376 270376
rect 309416 260908 309468 260914
rect 309416 260850 309468 260856
rect 309428 260778 309456 260850
rect 309416 260772 309468 260778
rect 309416 260714 309468 260720
rect 309324 251252 309376 251258
rect 309324 251194 309376 251200
rect 309336 251161 309364 251194
rect 309322 251152 309378 251161
rect 309322 251087 309378 251096
rect 309506 251152 309562 251161
rect 309506 251087 309562 251096
rect 309520 241534 309548 251087
rect 309508 241528 309560 241534
rect 309508 241470 309560 241476
rect 309600 241528 309652 241534
rect 309600 241470 309652 241476
rect 309612 234598 309640 241470
rect 309324 234592 309376 234598
rect 309324 234534 309376 234540
rect 309600 234592 309652 234598
rect 309600 234534 309652 234540
rect 309336 231810 309364 234534
rect 309324 231804 309376 231810
rect 309324 231746 309376 231752
rect 309508 222216 309560 222222
rect 309508 222158 309560 222164
rect 309520 211177 309548 222158
rect 309322 211168 309378 211177
rect 309322 211103 309378 211112
rect 309506 211168 309562 211177
rect 309506 211103 309562 211112
rect 309336 202978 309364 211103
rect 309324 202972 309376 202978
rect 309324 202914 309376 202920
rect 309416 202972 309468 202978
rect 309416 202914 309468 202920
rect 309428 201482 309456 202914
rect 309416 201476 309468 201482
rect 309416 201418 309468 201424
rect 309508 183592 309560 183598
rect 309508 183534 309560 183540
rect 309520 174078 309548 183534
rect 309508 174072 309560 174078
rect 309508 174014 309560 174020
rect 309508 173868 309560 173874
rect 309508 173810 309560 173816
rect 309520 154737 309548 173810
rect 309506 154728 309562 154737
rect 309506 154663 309562 154672
rect 309322 154592 309378 154601
rect 309322 154527 309378 154536
rect 309336 147694 309364 154527
rect 309324 147688 309376 147694
rect 309324 147630 309376 147636
rect 309416 147620 309468 147626
rect 309416 147562 309468 147568
rect 309428 143546 309456 147562
rect 309416 143540 309468 143546
rect 309416 143482 309468 143488
rect 309692 143540 309744 143546
rect 309692 143482 309744 143488
rect 309704 133929 309732 143482
rect 309506 133920 309562 133929
rect 309506 133855 309562 133864
rect 309690 133920 309746 133929
rect 309690 133855 309746 133864
rect 309520 124166 309548 133855
rect 309508 124160 309560 124166
rect 309508 124102 309560 124108
rect 309324 124024 309376 124030
rect 309324 123966 309376 123972
rect 309336 106282 309364 123966
rect 309232 106276 309284 106282
rect 309232 106218 309284 106224
rect 309324 106276 309376 106282
rect 309324 106218 309376 106224
rect 309244 104854 309272 106218
rect 309232 104848 309284 104854
rect 309232 104790 309284 104796
rect 309324 89684 309376 89690
rect 309324 89626 309376 89632
rect 309336 80102 309364 89626
rect 309324 80096 309376 80102
rect 309324 80038 309376 80044
rect 309232 77308 309284 77314
rect 309232 77250 309284 77256
rect 309244 67726 309272 77250
rect 309232 67720 309284 67726
rect 309232 67662 309284 67668
rect 309324 67652 309376 67658
rect 309324 67594 309376 67600
rect 309336 51134 309364 67594
rect 309324 51128 309376 51134
rect 309324 51070 309376 51076
rect 309416 50992 309468 50998
rect 309416 50934 309468 50940
rect 309428 46918 309456 50934
rect 309416 46912 309468 46918
rect 309416 46854 309468 46860
rect 309324 37324 309376 37330
rect 309324 37266 309376 37272
rect 309336 27554 309364 37266
rect 309336 27526 309456 27554
rect 309428 18193 309456 27526
rect 309414 18184 309470 18193
rect 309414 18119 309470 18128
rect 309322 18048 309378 18057
rect 309322 17983 309378 17992
rect 309336 14346 309364 17983
rect 309324 14340 309376 14346
rect 309324 14282 309376 14288
rect 309140 13660 309192 13666
rect 309140 13602 309192 13608
rect 307944 13388 307996 13394
rect 307944 13330 307996 13336
rect 306380 10192 306432 10198
rect 306380 10134 306432 10140
rect 302516 7268 302568 7274
rect 302516 7210 302568 7216
rect 308588 6520 308640 6526
rect 308588 6462 308640 6468
rect 305000 6452 305052 6458
rect 305000 6394 305052 6400
rect 301412 5432 301464 5438
rect 301412 5374 301464 5380
rect 300952 3732 301004 3738
rect 300952 3674 301004 3680
rect 301424 480 301452 5374
rect 303804 3664 303856 3670
rect 303804 3606 303856 3612
rect 302608 3256 302660 3262
rect 302608 3198 302660 3204
rect 302620 480 302648 3198
rect 303816 480 303844 3606
rect 305012 480 305040 6394
rect 307392 3732 307444 3738
rect 307392 3674 307444 3680
rect 306196 3324 306248 3330
rect 306196 3266 306248 3272
rect 306208 480 306236 3266
rect 307404 480 307432 3674
rect 308600 480 308628 6462
rect 309796 3738 309824 337894
rect 310532 10062 310560 340054
rect 311176 335646 311204 340054
rect 311900 337884 311952 337890
rect 311900 337826 311952 337832
rect 310704 335640 310756 335646
rect 310704 335582 310756 335588
rect 311164 335640 311216 335646
rect 311164 335582 311216 335588
rect 310716 311930 310744 335582
rect 310624 311902 310744 311930
rect 310624 311794 310652 311902
rect 310624 311766 310744 311794
rect 310716 299470 310744 311766
rect 310704 299464 310756 299470
rect 310704 299406 310756 299412
rect 310704 289876 310756 289882
rect 310704 289818 310756 289824
rect 310716 280158 310744 289818
rect 310704 280152 310756 280158
rect 310704 280094 310756 280100
rect 310704 270564 310756 270570
rect 310704 270506 310756 270512
rect 310716 260846 310744 270506
rect 310704 260840 310756 260846
rect 310704 260782 310756 260788
rect 310704 251252 310756 251258
rect 310704 251194 310756 251200
rect 310716 241505 310744 251194
rect 310702 241496 310758 241505
rect 310702 241431 310758 241440
rect 310886 241496 310942 241505
rect 310886 241431 310942 241440
rect 310900 231878 310928 241431
rect 310704 231872 310756 231878
rect 310704 231814 310756 231820
rect 310888 231872 310940 231878
rect 310888 231814 310940 231820
rect 310716 222193 310744 231814
rect 310702 222184 310758 222193
rect 310702 222119 310758 222128
rect 310886 222184 310942 222193
rect 310886 222119 310942 222128
rect 310900 212566 310928 222119
rect 310704 212560 310756 212566
rect 310704 212502 310756 212508
rect 310888 212560 310940 212566
rect 310888 212502 310940 212508
rect 310716 196058 310744 212502
rect 310624 196030 310744 196058
rect 310624 195922 310652 196030
rect 310624 195894 310744 195922
rect 310716 183569 310744 195894
rect 310702 183560 310758 183569
rect 310702 183495 310758 183504
rect 310886 183560 310942 183569
rect 310886 183495 310942 183504
rect 310900 173942 310928 183495
rect 310704 173936 310756 173942
rect 310704 173878 310756 173884
rect 310888 173936 310940 173942
rect 310888 173878 310940 173884
rect 310716 164218 310744 173878
rect 310704 164212 310756 164218
rect 310704 164154 310756 164160
rect 310888 164212 310940 164218
rect 310888 164154 310940 164160
rect 310900 154601 310928 164154
rect 310702 154592 310758 154601
rect 310702 154527 310758 154536
rect 310886 154592 310942 154601
rect 310886 154527 310942 154536
rect 310716 138122 310744 154527
rect 310624 138094 310744 138122
rect 310624 137986 310652 138094
rect 310624 137958 310744 137986
rect 310716 125594 310744 137958
rect 310704 125588 310756 125594
rect 310704 125530 310756 125536
rect 310704 118652 310756 118658
rect 310704 118594 310756 118600
rect 310716 99414 310744 118594
rect 310704 99408 310756 99414
rect 310704 99350 310756 99356
rect 310704 96688 310756 96694
rect 310704 96630 310756 96636
rect 310716 86970 310744 96630
rect 310704 86964 310756 86970
rect 310704 86906 310756 86912
rect 310704 77308 310756 77314
rect 310704 77250 310756 77256
rect 310716 67658 310744 77250
rect 310612 67652 310664 67658
rect 310612 67594 310664 67600
rect 310704 67652 310756 67658
rect 310704 67594 310756 67600
rect 310624 64870 310652 67594
rect 310612 64864 310664 64870
rect 310612 64806 310664 64812
rect 310888 55276 310940 55282
rect 310888 55218 310940 55224
rect 310900 47025 310928 55218
rect 310886 47016 310942 47025
rect 310886 46951 310942 46960
rect 310794 46744 310850 46753
rect 310794 46679 310850 46688
rect 310808 37330 310836 46679
rect 311808 40112 311860 40118
rect 311806 40080 311808 40089
rect 311860 40080 311862 40089
rect 311806 40015 311862 40024
rect 310612 37324 310664 37330
rect 310612 37266 310664 37272
rect 310796 37324 310848 37330
rect 310796 37266 310848 37272
rect 310624 22794 310652 37266
rect 310624 22766 310744 22794
rect 310716 13734 310744 22766
rect 310704 13728 310756 13734
rect 310704 13670 310756 13676
rect 310520 10056 310572 10062
rect 310520 9998 310572 10004
rect 311912 9994 311940 337826
rect 312004 14414 312032 340068
rect 312280 340054 312662 340082
rect 313306 340054 313412 340082
rect 312280 337890 312308 340054
rect 312268 337884 312320 337890
rect 312268 337826 312320 337832
rect 311992 14408 312044 14414
rect 311992 14350 312044 14356
rect 313384 12034 313412 340054
rect 313568 340054 313858 340082
rect 314120 340054 314502 340082
rect 314764 340054 315146 340082
rect 315408 340054 315698 340082
rect 316144 340054 316342 340082
rect 316696 340054 316986 340082
rect 317432 340054 317538 340082
rect 317708 340054 318182 340082
rect 318352 340054 318734 340082
rect 318812 340054 319378 340082
rect 319640 340054 320022 340082
rect 320284 340054 320574 340082
rect 320928 340054 321218 340082
rect 321572 340054 321862 340082
rect 321940 340054 322414 340082
rect 322952 340054 323058 340082
rect 323228 340054 323702 340082
rect 323872 340054 324254 340082
rect 324332 340054 324898 340082
rect 325068 340054 325542 340082
rect 325804 340054 326094 340082
rect 326448 340054 326738 340082
rect 327092 340054 327382 340082
rect 327460 340054 327934 340082
rect 328472 340054 328578 340082
rect 328748 340054 329222 340082
rect 329392 340054 329774 340082
rect 329852 340054 330418 340082
rect 330588 340054 331062 340082
rect 331232 340054 331614 340082
rect 313464 337884 313516 337890
rect 313464 337826 313516 337832
rect 313476 14278 313504 337826
rect 313464 14272 313516 14278
rect 313464 14214 313516 14220
rect 313372 12028 313424 12034
rect 313372 11970 313424 11976
rect 311900 9988 311952 9994
rect 311900 9930 311952 9936
rect 313568 6866 313596 340054
rect 314120 337890 314148 340054
rect 314108 337884 314160 337890
rect 314108 337826 314160 337832
rect 314660 337884 314712 337890
rect 314660 337826 314712 337832
rect 313556 6860 313608 6866
rect 313556 6802 313608 6808
rect 312176 6588 312228 6594
rect 312176 6530 312228 6536
rect 309784 3732 309836 3738
rect 309784 3674 309836 3680
rect 309784 3188 309836 3194
rect 309784 3130 309836 3136
rect 309796 480 309824 3130
rect 310980 2848 311032 2854
rect 310980 2790 311032 2796
rect 310992 480 311020 2790
rect 312188 480 312216 6530
rect 314672 6202 314700 337826
rect 314764 12102 314792 340054
rect 315408 337890 315436 340054
rect 316040 337952 316092 337958
rect 316040 337894 316092 337900
rect 315396 337884 315448 337890
rect 315396 337826 315448 337832
rect 316052 12170 316080 337894
rect 316144 14210 316172 340054
rect 316696 337958 316724 340054
rect 316684 337952 316736 337958
rect 316684 337894 316736 337900
rect 316684 337204 316736 337210
rect 316684 337146 316736 337152
rect 316132 14204 316184 14210
rect 316132 14146 316184 14152
rect 316040 12164 316092 12170
rect 316040 12106 316092 12112
rect 314752 12096 314804 12102
rect 314752 12038 314804 12044
rect 314580 6174 314700 6202
rect 314580 6118 314608 6174
rect 314568 6112 314620 6118
rect 314568 6054 314620 6060
rect 314660 6112 314712 6118
rect 314660 6054 314712 6060
rect 314672 4214 314700 6054
rect 316592 5976 316644 5982
rect 316592 5918 316644 5924
rect 315764 5500 315816 5506
rect 315764 5442 315816 5448
rect 314660 4208 314712 4214
rect 314660 4150 314712 4156
rect 314568 4140 314620 4146
rect 314568 4082 314620 4088
rect 313372 3120 313424 3126
rect 313372 3062 313424 3068
rect 313384 480 313412 3062
rect 314580 480 314608 4082
rect 315776 480 315804 5442
rect 316604 3806 316632 5918
rect 316696 4146 316724 337146
rect 317326 170096 317382 170105
rect 317326 170031 317382 170040
rect 317340 169862 317368 170031
rect 317328 169856 317380 169862
rect 317328 169798 317380 169804
rect 317326 157856 317382 157865
rect 317326 157791 317382 157800
rect 317340 157593 317368 157791
rect 317326 157584 317382 157593
rect 317326 157519 317382 157528
rect 317326 76256 317382 76265
rect 317326 76191 317328 76200
rect 317380 76191 317382 76200
rect 317328 76162 317380 76168
rect 317326 40216 317382 40225
rect 317326 40151 317382 40160
rect 317340 40118 317368 40151
rect 317328 40112 317380 40118
rect 317328 40054 317380 40060
rect 317326 29472 317382 29481
rect 317326 29407 317382 29416
rect 317340 28937 317368 29407
rect 317326 28928 317382 28937
rect 317326 28863 317382 28872
rect 317432 6050 317460 340054
rect 317604 337952 317656 337958
rect 317604 337894 317656 337900
rect 317616 12238 317644 337894
rect 317604 12232 317656 12238
rect 317604 12174 317656 12180
rect 317708 9042 317736 340054
rect 318352 337958 318380 340054
rect 318340 337952 318392 337958
rect 318340 337894 318392 337900
rect 318706 76256 318762 76265
rect 318706 76191 318762 76200
rect 318720 76129 318748 76191
rect 318706 76120 318762 76129
rect 318706 76055 318762 76064
rect 318706 29472 318762 29481
rect 318706 29407 318762 29416
rect 318720 29345 318748 29407
rect 318706 29336 318762 29345
rect 318706 29271 318762 29280
rect 318708 16720 318760 16726
rect 318706 16688 318708 16697
rect 318760 16688 318762 16697
rect 318706 16623 318762 16632
rect 317696 9036 317748 9042
rect 317696 8978 317748 8984
rect 318812 6882 318840 340054
rect 319640 335374 319668 340054
rect 320180 337952 320232 337958
rect 320180 337894 320232 337900
rect 318984 335368 319036 335374
rect 318984 335310 319036 335316
rect 319628 335368 319680 335374
rect 319628 335310 319680 335316
rect 318996 316146 319024 335310
rect 318904 316118 319024 316146
rect 318904 311846 318932 316118
rect 318892 311840 318944 311846
rect 318892 311782 318944 311788
rect 319076 311840 319128 311846
rect 319076 311782 319128 311788
rect 319088 309126 319116 311782
rect 319076 309120 319128 309126
rect 319076 309062 319128 309068
rect 318984 299532 319036 299538
rect 318984 299474 319036 299480
rect 318996 294658 319024 299474
rect 318996 294630 319116 294658
rect 319088 282826 319116 294630
rect 318996 282798 319116 282826
rect 318996 280158 319024 282798
rect 318984 280152 319036 280158
rect 318984 280094 319036 280100
rect 319076 280152 319128 280158
rect 319076 280094 319128 280100
rect 319088 263514 319116 280094
rect 318996 263486 319116 263514
rect 318996 260846 319024 263486
rect 318984 260840 319036 260846
rect 318984 260782 319036 260788
rect 319076 260840 319128 260846
rect 319076 260782 319128 260788
rect 319088 244202 319116 260782
rect 318996 244174 319116 244202
rect 318996 231878 319024 244174
rect 318984 231872 319036 231878
rect 318984 231814 319036 231820
rect 319076 231872 319128 231878
rect 319076 231814 319128 231820
rect 319088 224890 319116 231814
rect 318996 224862 319116 224890
rect 318996 212566 319024 224862
rect 318984 212560 319036 212566
rect 318984 212502 319036 212508
rect 319076 212560 319128 212566
rect 319076 212502 319128 212508
rect 319088 205578 319116 212502
rect 318996 205550 319116 205578
rect 318996 202842 319024 205550
rect 318984 202836 319036 202842
rect 318984 202778 319036 202784
rect 319076 202836 319128 202842
rect 319076 202778 319128 202784
rect 319088 167074 319116 202778
rect 318892 167068 318944 167074
rect 318892 167010 318944 167016
rect 319076 167068 319128 167074
rect 319076 167010 319128 167016
rect 318904 166954 318932 167010
rect 318904 166926 319024 166954
rect 318996 159338 319024 166926
rect 318996 159310 319116 159338
rect 319088 147694 319116 159310
rect 318892 147688 318944 147694
rect 319076 147688 319128 147694
rect 318944 147636 319024 147642
rect 318892 147630 319024 147636
rect 319076 147630 319128 147636
rect 318904 147614 319024 147630
rect 318996 137850 319024 147614
rect 318996 137822 319116 137850
rect 319088 128382 319116 137822
rect 318892 128376 318944 128382
rect 319076 128376 319128 128382
rect 318944 128324 319076 128330
rect 318892 128318 319128 128324
rect 318904 128302 319116 128318
rect 319088 114617 319116 128302
rect 319074 114608 319130 114617
rect 319074 114543 319130 114552
rect 319074 114472 319130 114481
rect 319074 114407 319130 114416
rect 319088 106350 319116 114407
rect 319076 106344 319128 106350
rect 319076 106286 319128 106292
rect 319076 106208 319128 106214
rect 319076 106150 319128 106156
rect 319088 104854 319116 106150
rect 319076 104848 319128 104854
rect 319076 104790 319128 104796
rect 319076 95260 319128 95266
rect 319076 95202 319128 95208
rect 319088 85490 319116 95202
rect 319088 85462 319208 85490
rect 319180 75954 319208 85462
rect 319076 75948 319128 75954
rect 319076 75890 319128 75896
rect 319168 75948 319220 75954
rect 319168 75890 319220 75896
rect 319088 67658 319116 75890
rect 318984 67652 319036 67658
rect 318984 67594 319036 67600
rect 319076 67652 319128 67658
rect 319076 67594 319128 67600
rect 318996 60738 319024 67594
rect 318996 60710 319116 60738
rect 319088 51082 319116 60710
rect 318904 51054 319116 51082
rect 318904 50946 318932 51054
rect 318904 50918 319024 50946
rect 318996 27606 319024 50918
rect 318984 27600 319036 27606
rect 318984 27542 319036 27548
rect 318984 18012 319036 18018
rect 318984 17954 319036 17960
rect 318996 14498 319024 17954
rect 319626 16824 319682 16833
rect 319626 16759 319682 16768
rect 319640 16726 319668 16759
rect 319628 16720 319680 16726
rect 319628 16662 319680 16668
rect 318996 14470 319116 14498
rect 319088 9110 319116 14470
rect 319076 9104 319128 9110
rect 319076 9046 319128 9052
rect 318812 6854 318932 6882
rect 318800 6724 318852 6730
rect 318800 6666 318852 6672
rect 317420 6044 317472 6050
rect 317420 5986 317472 5992
rect 316684 4140 316736 4146
rect 316684 4082 316736 4088
rect 316960 3868 317012 3874
rect 316960 3810 317012 3816
rect 316592 3800 316644 3806
rect 316592 3742 316644 3748
rect 316972 480 317000 3810
rect 318064 3800 318116 3806
rect 318064 3742 318116 3748
rect 318076 480 318104 3742
rect 318812 3398 318840 6666
rect 318904 5914 318932 6854
rect 320192 6798 320220 337894
rect 320284 12306 320312 340054
rect 320928 337958 320956 340054
rect 320916 337952 320968 337958
rect 320916 337894 320968 337900
rect 321466 325680 321522 325689
rect 321466 325615 321522 325624
rect 321480 316062 321508 325615
rect 321468 316056 321520 316062
rect 321466 316024 321468 316033
rect 321520 316024 321522 316033
rect 321466 315959 321522 315968
rect 321480 311234 321508 315959
rect 321468 311228 321520 311234
rect 321468 311170 321520 311176
rect 321468 168632 321520 168638
rect 321468 168574 321520 168580
rect 321480 159390 321508 168574
rect 321572 164393 321600 340054
rect 321940 335345 321968 340054
rect 322756 338020 322808 338026
rect 322756 337962 322808 337968
rect 321926 335336 321982 335345
rect 321926 335271 321982 335280
rect 322110 335336 322166 335345
rect 322110 335271 322166 335280
rect 322124 325718 322152 335271
rect 321652 325712 321704 325718
rect 321650 325680 321652 325689
rect 322112 325712 322164 325718
rect 321704 325680 321706 325689
rect 322112 325654 322164 325660
rect 321650 325615 321706 325624
rect 321756 316062 321784 316093
rect 321744 316056 321796 316062
rect 321650 316024 321706 316033
rect 321706 316004 321744 316010
rect 321706 315998 321796 316004
rect 321706 315982 321784 315998
rect 321650 315959 321706 315968
rect 321744 311228 321796 311234
rect 321744 311170 321796 311176
rect 321756 292670 321784 311170
rect 321744 292664 321796 292670
rect 321744 292606 321796 292612
rect 321744 292528 321796 292534
rect 321744 292470 321796 292476
rect 321756 280158 321784 292470
rect 321744 280152 321796 280158
rect 321744 280094 321796 280100
rect 321744 272196 321796 272202
rect 321744 272138 321796 272144
rect 321756 260846 321784 272138
rect 321744 260840 321796 260846
rect 321744 260782 321796 260788
rect 321744 251252 321796 251258
rect 321744 251194 321796 251200
rect 321756 241482 321784 251194
rect 321756 241454 321876 241482
rect 321848 234666 321876 241454
rect 321836 234660 321888 234666
rect 321836 234602 321888 234608
rect 321744 234592 321796 234598
rect 321744 234534 321796 234540
rect 321756 216034 321784 234534
rect 321744 216028 321796 216034
rect 321744 215970 321796 215976
rect 321928 216028 321980 216034
rect 321928 215970 321980 215976
rect 321940 211177 321968 215970
rect 321742 211168 321798 211177
rect 321742 211103 321798 211112
rect 321926 211168 321982 211177
rect 321926 211103 321982 211112
rect 321756 201482 321784 211103
rect 321744 201476 321796 201482
rect 321744 201418 321796 201424
rect 321928 201476 321980 201482
rect 321928 201418 321980 201424
rect 321940 191865 321968 201418
rect 321742 191856 321798 191865
rect 321742 191791 321798 191800
rect 321926 191856 321982 191865
rect 321926 191791 321982 191800
rect 321756 186454 321784 191791
rect 321744 186448 321796 186454
rect 321744 186390 321796 186396
rect 321652 183592 321704 183598
rect 321652 183534 321704 183540
rect 321664 173942 321692 183534
rect 321652 173936 321704 173942
rect 321652 173878 321704 173884
rect 321744 173936 321796 173942
rect 321744 173878 321796 173884
rect 321756 168638 321784 173878
rect 321744 168632 321796 168638
rect 321744 168574 321796 168580
rect 321558 164384 321614 164393
rect 321558 164319 321614 164328
rect 321558 164248 321614 164257
rect 321558 164183 321614 164192
rect 321468 159384 321520 159390
rect 321468 159326 321520 159332
rect 321466 87408 321522 87417
rect 321466 87343 321522 87352
rect 321480 87145 321508 87343
rect 321466 87136 321522 87145
rect 321466 87071 321522 87080
rect 320272 12300 320324 12306
rect 320272 12242 320324 12248
rect 321572 9178 321600 164183
rect 321744 159384 321796 159390
rect 321744 159326 321796 159332
rect 321756 149682 321784 159326
rect 321664 149654 321784 149682
rect 321664 143546 321692 149654
rect 321652 143540 321704 143546
rect 321652 143482 321704 143488
rect 321652 135244 321704 135250
rect 321652 135186 321704 135192
rect 321664 130098 321692 135186
rect 321664 130070 321784 130098
rect 321756 118862 321784 130070
rect 321744 118856 321796 118862
rect 321744 118798 321796 118804
rect 321744 114572 321796 114578
rect 321744 114514 321796 114520
rect 321756 51202 321784 114514
rect 321744 51196 321796 51202
rect 321744 51138 321796 51144
rect 321744 47048 321796 47054
rect 321744 46990 321796 46996
rect 321756 46918 321784 46990
rect 321652 46912 321704 46918
rect 321652 46854 321704 46860
rect 321744 46912 321796 46918
rect 321744 46854 321796 46860
rect 321664 29034 321692 46854
rect 321652 29028 321704 29034
rect 321652 28970 321704 28976
rect 321744 29028 321796 29034
rect 321744 28970 321796 28976
rect 321756 12374 321784 28970
rect 321744 12368 321796 12374
rect 321744 12310 321796 12316
rect 321560 9172 321612 9178
rect 321560 9114 321612 9120
rect 322572 9172 322624 9178
rect 322572 9114 322624 9120
rect 320180 6792 320232 6798
rect 320180 6734 320232 6740
rect 320180 6656 320232 6662
rect 320180 6598 320232 6604
rect 318892 5908 318944 5914
rect 318892 5850 318944 5856
rect 319260 4548 319312 4554
rect 319260 4490 319312 4496
rect 318800 3392 318852 3398
rect 318800 3334 318852 3340
rect 319272 480 319300 4490
rect 320192 3262 320220 6598
rect 321652 4140 321704 4146
rect 321652 4082 321704 4088
rect 320180 3256 320232 3262
rect 320180 3198 320232 3204
rect 320456 3052 320508 3058
rect 320456 2994 320508 3000
rect 320468 480 320496 2994
rect 321664 480 321692 4082
rect 322584 3942 322612 9114
rect 322664 5840 322716 5846
rect 322664 5782 322716 5788
rect 322676 4078 322704 5782
rect 322768 4146 322796 337962
rect 322952 6050 322980 340054
rect 323124 335640 323176 335646
rect 323124 335582 323176 335588
rect 323136 12442 323164 335582
rect 323124 12436 323176 12442
rect 323124 12378 323176 12384
rect 323228 9246 323256 340054
rect 323872 335646 323900 340054
rect 323860 335640 323912 335646
rect 323860 335582 323912 335588
rect 323216 9240 323268 9246
rect 323216 9182 323268 9188
rect 323584 9036 323636 9042
rect 323584 8978 323636 8984
rect 322940 6044 322992 6050
rect 322940 5986 322992 5992
rect 322848 4480 322900 4486
rect 322848 4422 322900 4428
rect 322756 4140 322808 4146
rect 322756 4082 322808 4088
rect 322664 4072 322716 4078
rect 322664 4014 322716 4020
rect 322572 3936 322624 3942
rect 322572 3878 322624 3884
rect 322860 480 322888 4422
rect 323596 3194 323624 8978
rect 324332 5778 324360 340054
rect 325068 331906 325096 340054
rect 325700 335640 325752 335646
rect 325700 335582 325752 335588
rect 324412 331900 324464 331906
rect 324412 331842 324464 331848
rect 325056 331900 325108 331906
rect 325056 331842 325108 331848
rect 324424 327162 324452 331842
rect 324424 327134 324544 327162
rect 324516 317665 324544 327134
rect 324502 317656 324558 317665
rect 324502 317591 324558 317600
rect 324410 317520 324466 317529
rect 324410 317455 324466 317464
rect 324424 316033 324452 317455
rect 324410 316024 324466 316033
rect 324410 315959 324466 315968
rect 324686 316024 324742 316033
rect 324686 315959 324742 315968
rect 324700 289882 324728 315959
rect 324504 289876 324556 289882
rect 324504 289818 324556 289824
rect 324688 289876 324740 289882
rect 324688 289818 324740 289824
rect 324516 289785 324544 289818
rect 324502 289776 324558 289785
rect 324502 289711 324558 289720
rect 324686 289776 324742 289785
rect 324686 289711 324742 289720
rect 324700 280226 324728 289711
rect 324412 280220 324464 280226
rect 324412 280162 324464 280168
rect 324688 280220 324740 280226
rect 324688 280162 324740 280168
rect 324424 280106 324452 280162
rect 324424 280078 324544 280106
rect 324516 276706 324544 280078
rect 324424 276678 324544 276706
rect 324424 263634 324452 276678
rect 324412 263628 324464 263634
rect 324412 263570 324464 263576
rect 324412 260908 324464 260914
rect 324412 260850 324464 260856
rect 324424 260794 324452 260850
rect 324424 260766 324544 260794
rect 324516 258754 324544 260766
rect 324424 258726 324544 258754
rect 324424 244322 324452 258726
rect 324412 244316 324464 244322
rect 324412 244258 324464 244264
rect 324412 241596 324464 241602
rect 324412 241538 324464 241544
rect 324424 241466 324452 241538
rect 324412 241460 324464 241466
rect 324412 241402 324464 241408
rect 324504 241460 324556 241466
rect 324504 241402 324556 241408
rect 324516 216034 324544 241402
rect 324504 216028 324556 216034
rect 324504 215970 324556 215976
rect 324688 216028 324740 216034
rect 324688 215970 324740 215976
rect 324700 211177 324728 215970
rect 324502 211168 324558 211177
rect 324502 211103 324558 211112
rect 324686 211168 324742 211177
rect 324686 211103 324742 211112
rect 324516 201482 324544 211103
rect 324504 201476 324556 201482
rect 324504 201418 324556 201424
rect 324688 201476 324740 201482
rect 324688 201418 324740 201424
rect 324700 191865 324728 201418
rect 324502 191856 324558 191865
rect 324502 191791 324558 191800
rect 324686 191856 324742 191865
rect 324686 191791 324742 191800
rect 324516 186454 324544 191791
rect 324504 186448 324556 186454
rect 324504 186390 324556 186396
rect 324412 183592 324464 183598
rect 324412 183534 324464 183540
rect 324424 173942 324452 183534
rect 324412 173936 324464 173942
rect 324412 173878 324464 173884
rect 324504 173936 324556 173942
rect 324504 173878 324556 173884
rect 324516 157418 324544 173878
rect 324504 157412 324556 157418
rect 324504 157354 324556 157360
rect 324412 157276 324464 157282
rect 324412 157218 324464 157224
rect 324424 147642 324452 157218
rect 324424 147614 324544 147642
rect 324516 135425 324544 147614
rect 324502 135416 324558 135425
rect 324502 135351 324558 135360
rect 324502 135280 324558 135289
rect 324502 135215 324558 135224
rect 324516 125769 324544 135215
rect 324502 125760 324558 125769
rect 324502 125695 324558 125704
rect 324502 125624 324558 125633
rect 324502 125559 324558 125568
rect 324516 118862 324544 125559
rect 324504 118856 324556 118862
rect 324504 118798 324556 118804
rect 324504 114572 324556 114578
rect 324504 114514 324556 114520
rect 324516 106282 324544 114514
rect 324504 106276 324556 106282
rect 324504 106218 324556 106224
rect 324504 96688 324556 96694
rect 324504 96630 324556 96636
rect 324516 86970 324544 96630
rect 324504 86964 324556 86970
rect 324504 86906 324556 86912
rect 324596 86964 324648 86970
rect 324596 86906 324648 86912
rect 324608 67674 324636 86906
rect 324516 67646 324636 67674
rect 324516 66230 324544 67646
rect 324504 66224 324556 66230
rect 324504 66166 324556 66172
rect 324504 56636 324556 56642
rect 324504 56578 324556 56584
rect 324516 40186 324544 56578
rect 324504 40180 324556 40186
rect 324504 40122 324556 40128
rect 324504 29028 324556 29034
rect 324504 28970 324556 28976
rect 324516 27606 324544 28970
rect 324504 27600 324556 27606
rect 324504 27542 324556 27548
rect 324412 18012 324464 18018
rect 324412 17954 324464 17960
rect 324424 9314 324452 17954
rect 324412 9308 324464 9314
rect 324412 9250 324464 9256
rect 325516 9172 325568 9178
rect 325516 9114 325568 9120
rect 325332 5908 325384 5914
rect 325332 5850 325384 5856
rect 324320 5772 324372 5778
rect 324320 5714 324372 5720
rect 325240 3936 325292 3942
rect 325240 3878 325292 3884
rect 324044 3392 324096 3398
rect 324044 3334 324096 3340
rect 323584 3188 323636 3194
rect 323584 3130 323636 3136
rect 324056 480 324084 3334
rect 325252 480 325280 3878
rect 325344 3738 325372 5850
rect 325332 3732 325384 3738
rect 325332 3674 325384 3680
rect 325528 3126 325556 9114
rect 325608 6792 325660 6798
rect 325608 6734 325660 6740
rect 325620 3330 325648 6734
rect 325712 5710 325740 335582
rect 325804 11694 325832 340054
rect 326448 335646 326476 340054
rect 326436 335640 326488 335646
rect 326436 335582 326488 335588
rect 326802 40216 326858 40225
rect 326802 40151 326858 40160
rect 326816 40066 326844 40151
rect 326986 40080 327042 40089
rect 326816 40038 326986 40066
rect 326986 40015 327042 40024
rect 325792 11688 325844 11694
rect 325792 11630 325844 11636
rect 327092 9382 327120 340054
rect 327460 331906 327488 340054
rect 327264 331900 327316 331906
rect 327264 331842 327316 331848
rect 327448 331900 327500 331906
rect 327448 331842 327500 331848
rect 327276 321638 327304 331842
rect 327264 321632 327316 321638
rect 327264 321574 327316 321580
rect 327264 321496 327316 321502
rect 327264 321438 327316 321444
rect 327276 317422 327304 321438
rect 327264 317416 327316 317422
rect 327264 317358 327316 317364
rect 327264 317280 327316 317286
rect 327264 317222 327316 317228
rect 327276 292670 327304 317222
rect 327264 292664 327316 292670
rect 327264 292606 327316 292612
rect 327264 292528 327316 292534
rect 327264 292470 327316 292476
rect 327276 280158 327304 292470
rect 327264 280152 327316 280158
rect 327264 280094 327316 280100
rect 327264 272196 327316 272202
rect 327264 272138 327316 272144
rect 327276 260846 327304 272138
rect 327264 260840 327316 260846
rect 327264 260782 327316 260788
rect 327264 251252 327316 251258
rect 327264 251194 327316 251200
rect 327276 230489 327304 251194
rect 327262 230480 327318 230489
rect 327262 230415 327318 230424
rect 327446 230480 327502 230489
rect 327446 230415 327502 230424
rect 327460 220862 327488 230415
rect 327264 220856 327316 220862
rect 327264 220798 327316 220804
rect 327448 220856 327500 220862
rect 327448 220798 327500 220804
rect 327276 202910 327304 220798
rect 327264 202904 327316 202910
rect 327264 202846 327316 202852
rect 327356 202904 327408 202910
rect 327356 202846 327408 202852
rect 327368 193254 327396 202846
rect 327264 193248 327316 193254
rect 327264 193190 327316 193196
rect 327356 193248 327408 193254
rect 327356 193190 327408 193196
rect 327276 186454 327304 193190
rect 327264 186448 327316 186454
rect 327264 186390 327316 186396
rect 327172 186312 327224 186318
rect 327172 186254 327224 186260
rect 327184 173942 327212 186254
rect 327172 173936 327224 173942
rect 327264 173936 327316 173942
rect 327224 173884 327264 173890
rect 327172 173878 327316 173884
rect 327184 173862 327304 173878
rect 327184 164218 327212 173862
rect 328366 170096 328422 170105
rect 328366 170031 328368 170040
rect 328420 170031 328422 170040
rect 328368 170002 328420 170008
rect 327172 164212 327224 164218
rect 327172 164154 327224 164160
rect 327264 164144 327316 164150
rect 327264 164086 327316 164092
rect 327276 162858 327304 164086
rect 327264 162852 327316 162858
rect 327264 162794 327316 162800
rect 327448 162852 327500 162858
rect 327448 162794 327500 162800
rect 327460 153241 327488 162794
rect 327262 153232 327318 153241
rect 327262 153167 327318 153176
rect 327446 153232 327502 153241
rect 327446 153167 327502 153176
rect 327276 149682 327304 153167
rect 327184 149654 327304 149682
rect 327184 124166 327212 149654
rect 327172 124160 327224 124166
rect 327172 124102 327224 124108
rect 327264 124160 327316 124166
rect 327264 124102 327316 124108
rect 327276 122806 327304 124102
rect 327264 122800 327316 122806
rect 327264 122742 327316 122748
rect 327264 113212 327316 113218
rect 327264 113154 327316 113160
rect 327276 104990 327304 113154
rect 327264 104984 327316 104990
rect 327264 104926 327316 104932
rect 327172 104916 327224 104922
rect 327172 104858 327224 104864
rect 327184 95266 327212 104858
rect 327172 95260 327224 95266
rect 327172 95202 327224 95208
rect 327264 95260 327316 95266
rect 327264 95202 327316 95208
rect 327276 85610 327304 95202
rect 327172 85604 327224 85610
rect 327172 85546 327224 85552
rect 327264 85604 327316 85610
rect 327264 85546 327316 85552
rect 327184 75954 327212 85546
rect 327172 75948 327224 75954
rect 327172 75890 327224 75896
rect 327264 75948 327316 75954
rect 327264 75890 327316 75896
rect 327276 60738 327304 75890
rect 327184 60710 327304 60738
rect 327184 60602 327212 60710
rect 327184 60574 327304 60602
rect 327276 51134 327304 60574
rect 327264 51128 327316 51134
rect 327264 51070 327316 51076
rect 327264 50992 327316 50998
rect 327264 50934 327316 50940
rect 327276 32450 327304 50934
rect 327184 32422 327304 32450
rect 327184 27606 327212 32422
rect 327172 27600 327224 27606
rect 327172 27542 327224 27548
rect 327264 27600 327316 27606
rect 327264 27542 327316 27548
rect 327276 11626 327304 27542
rect 327264 11620 327316 11626
rect 327264 11562 327316 11568
rect 327080 9376 327132 9382
rect 327080 9318 327132 9324
rect 327080 9240 327132 9246
rect 327080 9182 327132 9188
rect 325700 5704 325752 5710
rect 325700 5646 325752 5652
rect 326436 4412 326488 4418
rect 326436 4354 326488 4360
rect 325608 3324 325660 3330
rect 325608 3266 325660 3272
rect 325516 3120 325568 3126
rect 325516 3062 325568 3068
rect 326448 480 326476 4354
rect 327092 3874 327120 9182
rect 328472 5642 328500 340054
rect 328644 335640 328696 335646
rect 328644 335582 328696 335588
rect 328552 87168 328604 87174
rect 328550 87136 328552 87145
rect 328604 87136 328606 87145
rect 328550 87071 328606 87080
rect 328656 11558 328684 335582
rect 328644 11552 328696 11558
rect 328644 11494 328696 11500
rect 328748 9450 328776 340054
rect 329392 335646 329420 340054
rect 329380 335640 329432 335646
rect 329380 335582 329432 335588
rect 328736 9444 328788 9450
rect 328736 9386 328788 9392
rect 328552 9104 328604 9110
rect 328552 9046 328604 9052
rect 328460 5636 328512 5642
rect 328460 5578 328512 5584
rect 327080 3868 327132 3874
rect 327080 3810 327132 3816
rect 327632 3188 327684 3194
rect 327632 3130 327684 3136
rect 327644 480 327672 3130
rect 328564 3058 328592 9046
rect 329852 5574 329880 340054
rect 330588 328506 330616 340054
rect 330024 328500 330076 328506
rect 330024 328442 330076 328448
rect 330576 328500 330628 328506
rect 330576 328442 330628 328448
rect 330036 292670 330064 328442
rect 330024 292664 330076 292670
rect 330024 292606 330076 292612
rect 330024 292528 330076 292534
rect 330024 292470 330076 292476
rect 330036 273358 330064 292470
rect 330024 273352 330076 273358
rect 330024 273294 330076 273300
rect 330024 273216 330076 273222
rect 330024 273158 330076 273164
rect 330036 254046 330064 273158
rect 331128 260840 331180 260846
rect 331128 260782 331180 260788
rect 330024 254040 330076 254046
rect 330024 253982 330076 253988
rect 330024 253904 330076 253910
rect 330024 253846 330076 253852
rect 330036 241482 330064 253846
rect 331140 251297 331168 260782
rect 331126 251288 331182 251297
rect 331126 251223 331182 251232
rect 331126 251152 331182 251161
rect 331126 251087 331182 251096
rect 331140 241534 331168 251087
rect 331128 241528 331180 241534
rect 330036 241454 330156 241482
rect 331128 241470 331180 241476
rect 330128 234666 330156 241454
rect 330116 234660 330168 234666
rect 330116 234602 330168 234608
rect 330024 234592 330076 234598
rect 330024 234534 330076 234540
rect 330036 222170 330064 234534
rect 330036 222142 330156 222170
rect 330128 215354 330156 222142
rect 330116 215348 330168 215354
rect 330116 215290 330168 215296
rect 330024 215280 330076 215286
rect 330024 215222 330076 215228
rect 330036 193254 330064 215222
rect 331128 209772 331180 209778
rect 331128 209714 331180 209720
rect 331140 200161 331168 209714
rect 331126 200152 331182 200161
rect 331126 200087 331182 200096
rect 330024 193248 330076 193254
rect 330024 193190 330076 193196
rect 330116 193180 330168 193186
rect 330116 193122 330168 193128
rect 330128 183598 330156 193122
rect 329932 183592 329984 183598
rect 329932 183534 329984 183540
rect 330116 183592 330168 183598
rect 330116 183534 330168 183540
rect 329944 176730 329972 183534
rect 329932 176724 329984 176730
rect 329932 176666 329984 176672
rect 330024 176588 330076 176594
rect 330024 176530 330076 176536
rect 330036 169266 330064 176530
rect 330036 169238 330156 169266
rect 330128 164257 330156 169238
rect 329930 164248 329986 164257
rect 329930 164183 329932 164192
rect 329984 164183 329986 164192
rect 330114 164248 330170 164257
rect 330114 164183 330116 164192
rect 329932 164154 329984 164160
rect 330168 164183 330170 164192
rect 330116 164154 330168 164160
rect 330128 145081 330156 164154
rect 330114 145072 330170 145081
rect 330114 145007 330170 145016
rect 330022 144936 330078 144945
rect 330022 144871 330078 144880
rect 330036 128450 330064 144871
rect 330024 128444 330076 128450
rect 330024 128386 330076 128392
rect 329932 128308 329984 128314
rect 329932 128250 329984 128256
rect 329944 120290 329972 128250
rect 329932 120284 329984 120290
rect 329932 120226 329984 120232
rect 330024 106344 330076 106350
rect 330024 106286 330076 106292
rect 330036 99498 330064 106286
rect 330036 99470 330156 99498
rect 330128 99226 330156 99470
rect 330036 99198 330156 99226
rect 330036 60738 330064 99198
rect 329944 60710 330064 60738
rect 329944 60602 329972 60710
rect 329944 60574 330064 60602
rect 330036 56574 330064 60574
rect 329932 56568 329984 56574
rect 329932 56510 329984 56516
rect 330024 56568 330076 56574
rect 330024 56510 330076 56516
rect 329944 55214 329972 56510
rect 329932 55208 329984 55214
rect 329932 55150 329984 55156
rect 330024 46980 330076 46986
rect 330024 46922 330076 46928
rect 330036 44130 330064 46922
rect 330024 44124 330076 44130
rect 330024 44066 330076 44072
rect 330116 26308 330168 26314
rect 330116 26250 330168 26256
rect 330128 17950 330156 26250
rect 330116 17944 330168 17950
rect 330116 17886 330168 17892
rect 331232 11490 331260 340054
rect 331692 328506 331720 340190
rect 332612 340054 332902 340082
rect 333164 340054 333454 340082
rect 332508 338088 332560 338094
rect 332508 338030 332560 338036
rect 331496 328500 331548 328506
rect 331496 328442 331548 328448
rect 331680 328500 331732 328506
rect 331680 328442 331732 328448
rect 331508 309210 331536 328442
rect 331416 309182 331536 309210
rect 331416 304314 331444 309182
rect 331324 304286 331444 304314
rect 331324 302002 331352 304286
rect 331324 301974 331536 302002
rect 331508 299470 331536 301974
rect 331404 299464 331456 299470
rect 331404 299406 331456 299412
rect 331496 299464 331548 299470
rect 331496 299406 331548 299412
rect 331416 290057 331444 299406
rect 331402 290048 331458 290057
rect 331402 289983 331458 289992
rect 331310 289776 331366 289785
rect 331310 289711 331366 289720
rect 331324 282826 331352 289711
rect 331324 282798 331536 282826
rect 331508 280158 331536 282798
rect 331404 280152 331456 280158
rect 331404 280094 331456 280100
rect 331496 280152 331548 280158
rect 331496 280094 331548 280100
rect 331416 270745 331444 280094
rect 331402 270736 331458 270745
rect 331402 270671 331458 270680
rect 331310 270464 331366 270473
rect 331310 270399 331366 270408
rect 331324 263566 331352 270399
rect 331312 263560 331364 263566
rect 331312 263502 331364 263508
rect 331496 263492 331548 263498
rect 331496 263434 331548 263440
rect 331508 260846 331536 263434
rect 331496 260840 331548 260846
rect 331496 260782 331548 260788
rect 331496 241528 331548 241534
rect 331496 241470 331548 241476
rect 331508 231878 331536 241470
rect 331496 231872 331548 231878
rect 331496 231814 331548 231820
rect 331312 227792 331364 227798
rect 331312 227734 331364 227740
rect 331324 209778 331352 227734
rect 331312 209772 331364 209778
rect 331312 209714 331364 209720
rect 331402 200152 331458 200161
rect 331402 200087 331458 200096
rect 331416 183598 331444 200087
rect 331404 183592 331456 183598
rect 331404 183534 331456 183540
rect 331496 183592 331548 183598
rect 331496 183534 331548 183540
rect 331508 182170 331536 183534
rect 331496 182164 331548 182170
rect 331496 182106 331548 182112
rect 331588 182164 331640 182170
rect 331588 182106 331640 182112
rect 331600 154601 331628 182106
rect 331402 154592 331458 154601
rect 331402 154527 331404 154536
rect 331456 154527 331458 154536
rect 331586 154592 331642 154601
rect 331586 154527 331642 154536
rect 331404 154498 331456 154504
rect 331496 147484 331548 147490
rect 331496 147426 331548 147432
rect 331508 133906 331536 147426
rect 331416 133878 331536 133906
rect 331416 128194 331444 133878
rect 331416 128166 331536 128194
rect 331508 119354 331536 128166
rect 331508 119326 331628 119354
rect 331600 110922 331628 119326
rect 331508 110894 331628 110922
rect 331508 99634 331536 110894
rect 331416 99606 331536 99634
rect 331416 96642 331444 99606
rect 331416 96614 331536 96642
rect 331508 96506 331536 96614
rect 331324 96478 331536 96506
rect 331324 87038 331352 96478
rect 331312 87032 331364 87038
rect 331312 86974 331364 86980
rect 331404 87032 331456 87038
rect 331404 86974 331456 86980
rect 331416 67794 331444 86974
rect 331404 67788 331456 67794
rect 331404 67730 331456 67736
rect 331404 67652 331456 67658
rect 331404 67594 331456 67600
rect 331416 64870 331444 67594
rect 331404 64864 331456 64870
rect 331404 64806 331456 64812
rect 331496 48340 331548 48346
rect 331496 48282 331548 48288
rect 331508 37330 331536 48282
rect 331404 37324 331456 37330
rect 331404 37266 331456 37272
rect 331496 37324 331548 37330
rect 331496 37266 331548 37272
rect 331416 27606 331444 37266
rect 331312 27600 331364 27606
rect 331312 27542 331364 27548
rect 331404 27600 331456 27606
rect 331404 27542 331456 27548
rect 331324 13054 331352 27542
rect 331312 13048 331364 13054
rect 331312 12990 331364 12996
rect 331220 11484 331272 11490
rect 331220 11426 331272 11432
rect 329840 5568 329892 5574
rect 329840 5510 329892 5516
rect 330024 4344 330076 4350
rect 330024 4286 330076 4292
rect 328828 3256 328880 3262
rect 328828 3198 328880 3204
rect 328552 3052 328604 3058
rect 328552 2994 328604 3000
rect 328840 480 328868 3198
rect 330036 480 330064 4286
rect 332520 4146 332548 338030
rect 332612 9586 332640 340054
rect 333164 338076 333192 340054
rect 332796 338048 333192 338076
rect 332796 328522 332824 338048
rect 334084 335442 334112 340068
rect 334268 340054 334742 340082
rect 334072 335436 334124 335442
rect 334072 335378 334124 335384
rect 334164 335232 334216 335238
rect 334164 335174 334216 335180
rect 333980 331628 334032 331634
rect 333980 331570 334032 331576
rect 332704 328494 332824 328522
rect 332704 317422 332732 328494
rect 332692 317416 332744 317422
rect 332692 317358 332744 317364
rect 332876 317416 332928 317422
rect 332876 317358 332928 317364
rect 332888 306474 332916 317358
rect 332692 306468 332744 306474
rect 332692 306410 332744 306416
rect 332876 306468 332928 306474
rect 332876 306410 332928 306416
rect 332704 306377 332732 306410
rect 332690 306368 332746 306377
rect 332690 306303 332746 306312
rect 332966 306368 333022 306377
rect 332966 306303 333022 306312
rect 332980 296750 333008 306303
rect 332784 296744 332836 296750
rect 332784 296686 332836 296692
rect 332968 296744 333020 296750
rect 332968 296686 333020 296692
rect 332796 230466 332824 296686
rect 332796 230438 332916 230466
rect 332888 229090 332916 230438
rect 332876 229084 332928 229090
rect 332876 229026 332928 229032
rect 333060 229084 333112 229090
rect 333060 229026 333112 229032
rect 333072 219473 333100 229026
rect 332782 219464 332838 219473
rect 332782 219399 332838 219408
rect 333058 219464 333114 219473
rect 333058 219399 333114 219408
rect 332796 209930 332824 219399
rect 332796 209902 332916 209930
rect 332888 209778 332916 209902
rect 332692 209772 332744 209778
rect 332692 209714 332744 209720
rect 332876 209772 332928 209778
rect 332876 209714 332928 209720
rect 332704 200297 332732 209714
rect 332690 200288 332746 200297
rect 332690 200223 332746 200232
rect 332782 200152 332838 200161
rect 332782 200087 332838 200096
rect 332796 198694 332824 200087
rect 332784 198688 332836 198694
rect 332784 198630 332836 198636
rect 332784 189100 332836 189106
rect 332784 189042 332836 189048
rect 332796 182238 332824 189042
rect 332784 182232 332836 182238
rect 332784 182174 332836 182180
rect 332692 182164 332744 182170
rect 332692 182106 332744 182112
rect 332704 172514 332732 182106
rect 332692 172508 332744 172514
rect 332692 172450 332744 172456
rect 332784 172508 332836 172514
rect 332784 172450 332836 172456
rect 332796 157298 332824 172450
rect 332704 157270 332824 157298
rect 332704 157026 332732 157270
rect 332704 156998 332824 157026
rect 332796 118726 332824 156998
rect 333886 134464 333942 134473
rect 333886 134399 333942 134408
rect 333900 134065 333928 134399
rect 333886 134056 333942 134065
rect 333886 133991 333942 134000
rect 332784 118720 332836 118726
rect 332784 118662 332836 118668
rect 332784 118584 332836 118590
rect 332784 118526 332836 118532
rect 332796 99498 332824 118526
rect 332704 99470 332824 99498
rect 332704 99362 332732 99470
rect 332704 99334 332824 99362
rect 332796 80102 332824 99334
rect 332784 80096 332836 80102
rect 332784 80038 332836 80044
rect 332784 79960 332836 79966
rect 332784 79902 332836 79908
rect 332796 60738 332824 79902
rect 332704 60710 332824 60738
rect 332704 60602 332732 60710
rect 332704 60574 332824 60602
rect 332796 48414 332824 60574
rect 332784 48408 332836 48414
rect 332784 48350 332836 48356
rect 332692 48272 332744 48278
rect 332692 48214 332744 48220
rect 332704 42090 332732 48214
rect 332692 42084 332744 42090
rect 332692 42026 332744 42032
rect 332876 42084 332928 42090
rect 332876 42026 332928 42032
rect 332888 11422 332916 42026
rect 332876 11416 332928 11422
rect 332876 11358 332928 11364
rect 333992 9654 334020 331570
rect 334072 16720 334124 16726
rect 334070 16688 334072 16697
rect 334124 16688 334126 16697
rect 334070 16623 334126 16632
rect 334176 13802 334204 335174
rect 334268 331634 334296 340054
rect 334256 331628 334308 331634
rect 334256 331570 334308 331576
rect 334820 328506 334848 340190
rect 335464 340054 335938 340082
rect 336200 340054 336490 340082
rect 335360 335640 335412 335646
rect 335360 335582 335412 335588
rect 334440 328500 334492 328506
rect 334440 328442 334492 328448
rect 334808 328500 334860 328506
rect 334808 328442 334860 328448
rect 334452 317490 334480 328442
rect 334440 317484 334492 317490
rect 334440 317426 334492 317432
rect 334532 317484 334584 317490
rect 334532 317426 334584 317432
rect 334544 311250 334572 317426
rect 334268 311222 334572 311250
rect 334268 298178 334296 311222
rect 334256 298172 334308 298178
rect 334256 298114 334308 298120
rect 334256 296744 334308 296750
rect 334256 296686 334308 296692
rect 334268 289814 334296 296686
rect 334256 289808 334308 289814
rect 334256 289750 334308 289756
rect 334440 282804 334492 282810
rect 334440 282746 334492 282752
rect 334452 280158 334480 282746
rect 334440 280152 334492 280158
rect 334440 280094 334492 280100
rect 334348 273216 334400 273222
rect 334348 273158 334400 273164
rect 334360 263634 334388 273158
rect 334348 263628 334400 263634
rect 334348 263570 334400 263576
rect 334440 263492 334492 263498
rect 334440 263434 334492 263440
rect 334452 260846 334480 263434
rect 334440 260840 334492 260846
rect 334440 260782 334492 260788
rect 334348 251320 334400 251326
rect 334348 251262 334400 251268
rect 334360 251190 334388 251262
rect 334348 251184 334400 251190
rect 334348 251126 334400 251132
rect 334348 244180 334400 244186
rect 334348 244122 334400 244128
rect 334360 232014 334388 244122
rect 334348 232008 334400 232014
rect 334348 231950 334400 231956
rect 334440 231872 334492 231878
rect 334440 231814 334492 231820
rect 334452 226930 334480 231814
rect 334360 226902 334480 226930
rect 334360 219434 334388 226902
rect 334348 219428 334400 219434
rect 334348 219370 334400 219376
rect 334440 212492 334492 212498
rect 334440 212434 334492 212440
rect 334452 209794 334480 212434
rect 334452 209766 334572 209794
rect 334544 205578 334572 209766
rect 334452 205550 334572 205578
rect 334452 193254 334480 205550
rect 334348 193248 334400 193254
rect 334348 193190 334400 193196
rect 334440 193248 334492 193254
rect 334440 193190 334492 193196
rect 334360 183598 334388 193190
rect 334348 183592 334400 183598
rect 334348 183534 334400 183540
rect 334440 183592 334492 183598
rect 334440 183534 334492 183540
rect 334452 182170 334480 183534
rect 334440 182164 334492 182170
rect 334440 182106 334492 182112
rect 334532 182164 334584 182170
rect 334532 182106 334584 182112
rect 334544 161430 334572 182106
rect 334532 161424 334584 161430
rect 334532 161366 334584 161372
rect 334624 153196 334676 153202
rect 334624 153138 334676 153144
rect 334636 151774 334664 153138
rect 334624 151768 334676 151774
rect 334624 151710 334676 151716
rect 334440 142180 334492 142186
rect 334440 142122 334492 142128
rect 334452 133890 334480 142122
rect 334440 133884 334492 133890
rect 334440 133826 334492 133832
rect 334440 124228 334492 124234
rect 334440 124170 334492 124176
rect 334452 119354 334480 124170
rect 334452 119326 334572 119354
rect 334544 110922 334572 119326
rect 334452 110894 334572 110922
rect 334452 99498 334480 110894
rect 334452 99470 334572 99498
rect 334544 96506 334572 99470
rect 334452 96478 334572 96506
rect 334452 87038 334480 96478
rect 334256 87032 334308 87038
rect 334256 86974 334308 86980
rect 334440 87032 334492 87038
rect 334440 86974 334492 86980
rect 334268 85542 334296 86974
rect 334256 85536 334308 85542
rect 334256 85478 334308 85484
rect 334440 79348 334492 79354
rect 334440 79290 334492 79296
rect 334452 74526 334480 79290
rect 334440 74520 334492 74526
rect 334440 74462 334492 74468
rect 334348 65000 334400 65006
rect 334348 64942 334400 64948
rect 334360 64870 334388 64942
rect 334348 64864 334400 64870
rect 334348 64806 334400 64812
rect 334440 48340 334492 48346
rect 334440 48282 334492 48288
rect 334452 37330 334480 48282
rect 334348 37324 334400 37330
rect 334348 37266 334400 37272
rect 334440 37324 334492 37330
rect 334440 37266 334492 37272
rect 334360 17950 334388 37266
rect 334348 17944 334400 17950
rect 334348 17886 334400 17892
rect 334164 13796 334216 13802
rect 334164 13738 334216 13744
rect 333980 9648 334032 9654
rect 333980 9590 334032 9596
rect 332600 9580 332652 9586
rect 332600 9522 332652 9528
rect 334716 8968 334768 8974
rect 334716 8910 334768 8916
rect 333612 4276 333664 4282
rect 333612 4218 333664 4224
rect 331220 4140 331272 4146
rect 331220 4082 331272 4088
rect 332508 4140 332560 4146
rect 332508 4082 332560 4088
rect 331232 480 331260 4082
rect 332416 3868 332468 3874
rect 332416 3810 332468 3816
rect 332428 480 332456 3810
rect 333624 480 333652 4218
rect 334728 480 334756 8910
rect 335372 8838 335400 335582
rect 335464 12986 335492 340054
rect 336200 335646 336228 340054
rect 337120 337278 337148 340068
rect 337108 337272 337160 337278
rect 337108 337214 337160 337220
rect 336188 335640 336240 335646
rect 336188 335582 336240 335588
rect 337212 328506 337240 340190
rect 338224 340054 338330 340082
rect 336924 328500 336976 328506
rect 336924 328442 336976 328448
rect 337200 328500 337252 328506
rect 337200 328442 337252 328448
rect 336936 309194 336964 328442
rect 336832 309188 336884 309194
rect 336832 309130 336884 309136
rect 336924 309188 336976 309194
rect 336924 309130 336976 309136
rect 336844 302274 336872 309130
rect 336752 302246 336872 302274
rect 336752 302138 336780 302246
rect 336752 302110 336872 302138
rect 336844 282962 336872 302110
rect 336752 282934 336872 282962
rect 336752 282826 336780 282934
rect 336752 282798 336872 282826
rect 336844 263650 336872 282798
rect 336752 263622 336872 263650
rect 336752 263514 336780 263622
rect 336752 263486 336872 263514
rect 336844 244338 336872 263486
rect 336752 244310 336872 244338
rect 336752 244202 336780 244310
rect 336752 244174 336872 244202
rect 336844 225026 336872 244174
rect 336752 224998 336872 225026
rect 336752 224890 336780 224998
rect 336752 224862 336872 224890
rect 336844 205698 336872 224862
rect 336832 205692 336884 205698
rect 336832 205634 336884 205640
rect 336740 204400 336792 204406
rect 336738 204368 336740 204377
rect 338120 204400 338172 204406
rect 336792 204368 336794 204377
rect 336738 204303 336794 204312
rect 338118 204368 338120 204377
rect 338172 204368 338174 204377
rect 338118 204303 338174 204312
rect 336832 202904 336884 202910
rect 336832 202846 336884 202852
rect 336844 193254 336872 202846
rect 336740 193248 336792 193254
rect 336740 193190 336792 193196
rect 336832 193248 336884 193254
rect 336832 193190 336884 193196
rect 336752 183598 336780 193190
rect 336740 183592 336792 183598
rect 336740 183534 336792 183540
rect 336832 183592 336884 183598
rect 336832 183534 336884 183540
rect 336844 182170 336872 183534
rect 336832 182164 336884 182170
rect 336832 182106 336884 182112
rect 336832 176588 336884 176594
rect 336832 176530 336884 176536
rect 336646 170096 336702 170105
rect 336646 170031 336648 170040
rect 336700 170031 336702 170040
rect 336648 170002 336700 170008
rect 336844 138122 336872 176530
rect 336752 138094 336872 138122
rect 336752 137986 336780 138094
rect 336752 137958 336872 137986
rect 336844 118726 336872 137958
rect 338026 134056 338082 134065
rect 338082 134014 338160 134042
rect 338026 133991 338082 134000
rect 338132 133521 338160 134014
rect 338118 133512 338174 133521
rect 338118 133447 338174 133456
rect 336832 118720 336884 118726
rect 336832 118662 336884 118668
rect 336832 118584 336884 118590
rect 336832 118526 336884 118532
rect 336738 110800 336794 110809
rect 336738 110735 336740 110744
rect 336792 110735 336794 110744
rect 336740 110706 336792 110712
rect 336844 80102 336872 118526
rect 338026 87272 338082 87281
rect 338026 87207 338082 87216
rect 338040 87174 338068 87207
rect 338028 87168 338080 87174
rect 338028 87110 338080 87116
rect 336832 80096 336884 80102
rect 336832 80038 336884 80044
rect 336832 79960 336884 79966
rect 336832 79902 336884 79908
rect 336844 60738 336872 79902
rect 337474 63608 337530 63617
rect 337474 63543 337476 63552
rect 337528 63543 337530 63552
rect 337476 63514 337528 63520
rect 336752 60710 336872 60738
rect 336752 60602 336780 60710
rect 336752 60574 336872 60602
rect 336844 27690 336872 60574
rect 336752 27662 336872 27690
rect 336752 24857 336780 27662
rect 336554 24848 336610 24857
rect 336554 24783 336610 24792
rect 336738 24848 336794 24857
rect 336738 24783 336794 24792
rect 336568 15230 336596 24783
rect 338120 16720 338172 16726
rect 338118 16688 338120 16697
rect 338172 16688 338174 16697
rect 338118 16623 338174 16632
rect 336556 15224 336608 15230
rect 336556 15166 336608 15172
rect 336832 15224 336884 15230
rect 336832 15166 336884 15172
rect 335452 12980 335504 12986
rect 335452 12922 335504 12928
rect 336844 12850 336872 15166
rect 336832 12844 336884 12850
rect 336832 12786 336884 12792
rect 338224 8906 338252 340054
rect 338960 337346 338988 340068
rect 339618 340054 339724 340082
rect 338948 337340 339000 337346
rect 338948 337282 339000 337288
rect 339408 337272 339460 337278
rect 339408 337214 339460 337220
rect 338212 8900 338264 8906
rect 338212 8842 338264 8848
rect 335360 8832 335412 8838
rect 335360 8774 335412 8780
rect 337108 4208 337160 4214
rect 337108 4150 337160 4156
rect 335912 3120 335964 3126
rect 335912 3062 335964 3068
rect 335924 480 335952 3062
rect 337120 480 337148 4150
rect 339420 3058 339448 337214
rect 339500 333260 339552 333266
rect 339500 333202 339552 333208
rect 339512 4758 339540 333202
rect 339696 12918 339724 340054
rect 339788 340054 340170 340082
rect 340432 340054 340814 340082
rect 340984 340054 341458 340082
rect 341720 340054 342010 340082
rect 342272 340054 342654 340082
rect 343008 340054 343298 340082
rect 343744 340054 343850 340082
rect 344112 340054 344494 340082
rect 339684 12912 339736 12918
rect 339684 12854 339736 12860
rect 339788 8770 339816 340054
rect 340432 333266 340460 340054
rect 340880 335640 340932 335646
rect 340880 335582 340932 335588
rect 340420 333260 340472 333266
rect 340420 333202 340472 333208
rect 340786 87272 340842 87281
rect 340786 87207 340842 87216
rect 340800 87174 340828 87207
rect 340788 87168 340840 87174
rect 340788 87110 340840 87116
rect 339776 8764 339828 8770
rect 339776 8706 339828 8712
rect 340892 8634 340920 335582
rect 340984 12782 341012 340054
rect 341720 335646 341748 340054
rect 341708 335640 341760 335646
rect 341708 335582 341760 335588
rect 341062 40216 341118 40225
rect 341062 40151 341118 40160
rect 341076 39817 341104 40151
rect 341062 39808 341118 39817
rect 341062 39743 341118 39752
rect 340972 12776 341024 12782
rect 340972 12718 341024 12724
rect 340880 8628 340932 8634
rect 340880 8570 340932 8576
rect 342272 4865 342300 340054
rect 343008 328506 343036 340054
rect 343640 332240 343692 332246
rect 343640 332182 343692 332188
rect 342628 328500 342680 328506
rect 342628 328442 342680 328448
rect 342996 328500 343048 328506
rect 342996 328442 343048 328448
rect 342640 309262 342668 328442
rect 342628 309256 342680 309262
rect 342628 309198 342680 309204
rect 342444 309188 342496 309194
rect 342444 309130 342496 309136
rect 342456 309058 342484 309130
rect 342444 309052 342496 309058
rect 342444 308994 342496 309000
rect 342536 299600 342588 299606
rect 342536 299542 342588 299548
rect 342548 299452 342576 299542
rect 342548 299424 342760 299452
rect 342732 289898 342760 299424
rect 342548 289870 342760 289898
rect 342548 282946 342576 289870
rect 342536 282940 342588 282946
rect 342536 282882 342588 282888
rect 342536 280288 342588 280294
rect 342536 280230 342588 280236
rect 342548 280140 342576 280230
rect 342548 280112 342760 280140
rect 342732 270586 342760 280112
rect 342548 270558 342760 270586
rect 342548 263634 342576 270558
rect 342536 263628 342588 263634
rect 342536 263570 342588 263576
rect 342536 260908 342588 260914
rect 342536 260850 342588 260856
rect 342548 260778 342576 260850
rect 342536 260772 342588 260778
rect 342536 260714 342588 260720
rect 342444 251252 342496 251258
rect 342444 251194 342496 251200
rect 342456 251161 342484 251194
rect 342442 251152 342498 251161
rect 342442 251087 342498 251096
rect 342626 251152 342682 251161
rect 342626 251087 342682 251096
rect 342640 241516 342668 251087
rect 342640 241488 342760 241516
rect 342732 234546 342760 241488
rect 342456 234518 342760 234546
rect 342456 231849 342484 234518
rect 342442 231840 342498 231849
rect 342442 231775 342498 231784
rect 342718 231840 342774 231849
rect 342718 231775 342774 231784
rect 342732 212809 342760 231775
rect 342718 212800 342774 212809
rect 342718 212735 342774 212744
rect 342442 212562 342498 212571
rect 342442 212497 342498 212506
rect 342456 207890 342484 212497
rect 342456 207862 342760 207890
rect 342732 196654 342760 207862
rect 342720 196648 342772 196654
rect 342720 196590 342772 196596
rect 342904 196648 342956 196654
rect 342904 196590 342956 196596
rect 342916 191865 342944 196590
rect 342718 191856 342774 191865
rect 342718 191791 342774 191800
rect 342902 191856 342958 191865
rect 342902 191791 342958 191800
rect 342732 186946 342760 191791
rect 342732 186918 342944 186946
rect 342916 172553 342944 186918
rect 343546 181384 343602 181393
rect 343546 181319 343602 181328
rect 343560 181257 343588 181319
rect 343546 181248 343602 181257
rect 343546 181183 343602 181192
rect 342534 172544 342590 172553
rect 342534 172479 342536 172488
rect 342588 172479 342590 172488
rect 342902 172544 342958 172553
rect 342902 172479 342958 172488
rect 342536 172450 342588 172456
rect 342352 162920 342404 162926
rect 342352 162862 342404 162868
rect 342364 154601 342392 162862
rect 342350 154592 342406 154601
rect 342350 154527 342406 154536
rect 342534 154592 342590 154601
rect 342534 154527 342590 154536
rect 342548 138122 342576 154527
rect 342456 138094 342576 138122
rect 342456 137986 342484 138094
rect 342456 137958 342576 137986
rect 342548 130370 342576 137958
rect 342456 130342 342576 130370
rect 342456 125594 342484 130342
rect 342444 125588 342496 125594
rect 342444 125530 342496 125536
rect 342628 125588 342680 125594
rect 342628 125530 342680 125536
rect 342640 124166 342668 125530
rect 342628 124160 342680 124166
rect 342628 124102 342680 124108
rect 342628 114572 342680 114578
rect 342628 114514 342680 114520
rect 342640 106350 342668 114514
rect 342536 106344 342588 106350
rect 342536 106286 342588 106292
rect 342628 106344 342680 106350
rect 342628 106286 342680 106292
rect 342548 99498 342576 106286
rect 342456 99470 342576 99498
rect 342456 89826 342484 99470
rect 342444 89820 342496 89826
rect 342444 89762 342496 89768
rect 342444 89684 342496 89690
rect 342444 89626 342496 89632
rect 342456 86986 342484 89626
rect 342456 86970 342576 86986
rect 342456 86964 342588 86970
rect 342456 86958 342536 86964
rect 342536 86906 342588 86912
rect 342536 80028 342588 80034
rect 342536 79970 342588 79976
rect 342548 60738 342576 79970
rect 342456 60710 342576 60738
rect 342456 60602 342484 60710
rect 342456 60574 342576 60602
rect 342548 55214 342576 60574
rect 342536 55208 342588 55214
rect 342536 55150 342588 55156
rect 342444 45620 342496 45626
rect 342444 45562 342496 45568
rect 342456 45506 342484 45562
rect 342364 45478 342484 45506
rect 342364 37210 342392 45478
rect 342364 37182 342484 37210
rect 342456 32434 342484 37182
rect 342444 32428 342496 32434
rect 342444 32370 342496 32376
rect 342352 19372 342404 19378
rect 342352 19314 342404 19320
rect 342364 12714 342392 19314
rect 342352 12708 342404 12714
rect 342352 12650 342404 12656
rect 342258 4856 342314 4865
rect 342258 4791 342314 4800
rect 339500 4752 339552 4758
rect 339500 4694 339552 4700
rect 340696 4752 340748 4758
rect 340696 4694 340748 4700
rect 339500 4072 339552 4078
rect 339500 4014 339552 4020
rect 338304 3052 338356 3058
rect 338304 2994 338356 3000
rect 339408 3052 339460 3058
rect 339408 2994 339460 3000
rect 338316 480 338344 2994
rect 339512 480 339540 4014
rect 340708 480 340736 4694
rect 343652 4690 343680 332182
rect 343744 8702 343772 340054
rect 344112 332246 344140 340054
rect 345020 335640 345072 335646
rect 345020 335582 345072 335588
rect 344100 332240 344152 332246
rect 344100 332182 344152 332188
rect 344926 123312 344982 123321
rect 344926 123247 344982 123256
rect 344940 122913 344968 123247
rect 344926 122904 344982 122913
rect 344926 122839 344982 122848
rect 344926 63608 344982 63617
rect 344926 63543 344928 63552
rect 344980 63543 344982 63552
rect 344928 63514 344980 63520
rect 343732 8696 343784 8702
rect 343732 8638 343784 8644
rect 343640 4684 343692 4690
rect 343640 4626 343692 4632
rect 344284 4684 344336 4690
rect 344284 4626 344336 4632
rect 343088 3188 343140 3194
rect 343088 3130 343140 3136
rect 341892 2984 341944 2990
rect 341892 2926 341944 2932
rect 341904 480 341932 2926
rect 343100 480 343128 3130
rect 344296 480 344324 4626
rect 345032 4622 345060 335582
rect 345124 7206 345152 340068
rect 345216 340054 345690 340082
rect 345952 340054 346334 340082
rect 346412 340054 346978 340082
rect 347148 340054 347530 340082
rect 347792 340054 348174 340082
rect 345216 8566 345244 340054
rect 345952 335646 345980 340054
rect 346308 337272 346360 337278
rect 346308 337214 346360 337220
rect 345940 335640 345992 335646
rect 345940 335582 345992 335588
rect 345938 123312 345994 123321
rect 345938 123247 345940 123256
rect 345992 123247 345994 123256
rect 345940 123218 345992 123224
rect 346216 110764 346268 110770
rect 346216 110706 346268 110712
rect 346228 110537 346256 110706
rect 346214 110528 346270 110537
rect 346214 110463 346270 110472
rect 346320 76514 346348 337214
rect 346228 76486 346348 76514
rect 346228 76022 346256 76486
rect 346216 76016 346268 76022
rect 346216 75958 346268 75964
rect 346308 75948 346360 75954
rect 346308 75890 346360 75896
rect 346216 63640 346268 63646
rect 346214 63608 346216 63617
rect 346268 63608 346270 63617
rect 346214 63543 346270 63552
rect 345204 8560 345256 8566
rect 345204 8502 345256 8508
rect 345112 7200 345164 7206
rect 345112 7142 345164 7148
rect 345020 4616 345072 4622
rect 345020 4558 345072 4564
rect 346320 746 346348 75890
rect 346412 7138 346440 340054
rect 347148 331242 347176 340054
rect 346596 331214 347176 331242
rect 346596 311846 346624 331214
rect 346584 311840 346636 311846
rect 346584 311782 346636 311788
rect 346584 309188 346636 309194
rect 346584 309130 346636 309136
rect 346596 299470 346624 309130
rect 346584 299464 346636 299470
rect 346584 299406 346636 299412
rect 346584 289876 346636 289882
rect 346584 289818 346636 289824
rect 346596 280158 346624 289818
rect 346584 280152 346636 280158
rect 346584 280094 346636 280100
rect 346584 270564 346636 270570
rect 346584 270506 346636 270512
rect 346596 260846 346624 270506
rect 347686 267744 347742 267753
rect 347686 267679 347742 267688
rect 346584 260840 346636 260846
rect 346584 260782 346636 260788
rect 347700 258097 347728 267679
rect 347686 258088 347742 258097
rect 347686 258023 347742 258032
rect 346584 251252 346636 251258
rect 346584 251194 346636 251200
rect 346596 241505 346624 251194
rect 346582 241496 346638 241505
rect 346582 241431 346638 241440
rect 346766 241496 346822 241505
rect 346766 241431 346822 241440
rect 346780 231878 346808 241431
rect 346584 231872 346636 231878
rect 346584 231814 346636 231820
rect 346768 231872 346820 231878
rect 346768 231814 346820 231820
rect 346596 222193 346624 231814
rect 346582 222184 346638 222193
rect 346582 222119 346638 222128
rect 346766 222184 346822 222193
rect 346766 222119 346822 222128
rect 346780 212566 346808 222119
rect 346584 212560 346636 212566
rect 346584 212502 346636 212508
rect 346768 212560 346820 212566
rect 346768 212502 346820 212508
rect 346596 202881 346624 212502
rect 346582 202872 346638 202881
rect 346582 202807 346638 202816
rect 346766 202872 346822 202881
rect 346766 202807 346822 202816
rect 346780 193254 346808 202807
rect 346584 193248 346636 193254
rect 346584 193190 346636 193196
rect 346768 193248 346820 193254
rect 346768 193190 346820 193196
rect 346596 176662 346624 193190
rect 346584 176656 346636 176662
rect 346584 176598 346636 176604
rect 346584 176520 346636 176526
rect 346584 176462 346636 176468
rect 346596 157350 346624 176462
rect 346584 157344 346636 157350
rect 346584 157286 346636 157292
rect 346584 157208 346636 157214
rect 346584 157150 346636 157156
rect 346596 138122 346624 157150
rect 346504 138094 346624 138122
rect 346504 137986 346532 138094
rect 346504 137958 346624 137986
rect 346596 118726 346624 137958
rect 346584 118720 346636 118726
rect 346584 118662 346636 118668
rect 346584 118584 346636 118590
rect 346584 118526 346636 118532
rect 346596 99498 346624 118526
rect 346504 99470 346624 99498
rect 346504 99362 346532 99470
rect 346504 99334 346624 99362
rect 346596 86970 346624 99334
rect 346584 86964 346636 86970
rect 346584 86906 346636 86912
rect 346584 80028 346636 80034
rect 346584 79970 346636 79976
rect 346596 66230 346624 79970
rect 346584 66224 346636 66230
rect 346584 66166 346636 66172
rect 346676 66224 346728 66230
rect 346676 66166 346728 66172
rect 346490 63880 346546 63889
rect 346490 63815 346546 63824
rect 346504 63646 346532 63815
rect 346492 63640 346544 63646
rect 346492 63582 346544 63588
rect 346688 60704 346716 66166
rect 346596 60676 346716 60704
rect 346596 33810 346624 60676
rect 346504 33782 346624 33810
rect 346504 27606 346532 33782
rect 346492 27600 346544 27606
rect 346492 27542 346544 27548
rect 346492 18012 346544 18018
rect 346492 17954 346544 17960
rect 346504 9654 346532 17954
rect 347688 16856 347740 16862
rect 347686 16824 347688 16833
rect 347740 16824 347742 16833
rect 347686 16759 347742 16768
rect 346492 9648 346544 9654
rect 346492 9590 346544 9596
rect 346492 7268 346544 7274
rect 346492 7210 346544 7216
rect 346400 7132 346452 7138
rect 346400 7074 346452 7080
rect 346504 3398 346532 7210
rect 347792 4826 347820 340054
rect 348804 336802 348832 340068
rect 349264 340054 349370 340082
rect 349632 340054 350014 340082
rect 347964 336796 348016 336802
rect 347964 336738 348016 336744
rect 348792 336796 348844 336802
rect 348792 336738 348844 336744
rect 347976 333985 348004 336738
rect 349160 335640 349212 335646
rect 349160 335582 349212 335588
rect 347962 333976 348018 333985
rect 347962 333911 348018 333920
rect 348238 333976 348294 333985
rect 348238 333911 348294 333920
rect 348252 324358 348280 333911
rect 348056 324352 348108 324358
rect 348056 324294 348108 324300
rect 348240 324352 348292 324358
rect 348240 324294 348292 324300
rect 348068 321638 348096 324294
rect 348056 321632 348108 321638
rect 348056 321574 348108 321580
rect 347964 321564 348016 321570
rect 347964 321506 348016 321512
rect 347976 299606 348004 321506
rect 347964 299600 348016 299606
rect 347964 299542 348016 299548
rect 347964 299396 348016 299402
rect 347964 299338 348016 299344
rect 347976 298110 348004 299338
rect 347964 298104 348016 298110
rect 347964 298046 348016 298052
rect 348056 288448 348108 288454
rect 348056 288390 348108 288396
rect 348068 280158 348096 288390
rect 348056 280152 348108 280158
rect 348056 280094 348108 280100
rect 348148 280152 348200 280158
rect 348148 280094 348200 280100
rect 348160 270586 348188 280094
rect 348160 270558 348280 270586
rect 348252 267782 348280 270558
rect 347872 267776 347924 267782
rect 347870 267744 347872 267753
rect 348240 267776 348292 267782
rect 347924 267744 347926 267753
rect 348240 267718 348292 267724
rect 347870 267679 347926 267688
rect 348054 258088 348110 258097
rect 348054 258023 348110 258032
rect 348068 250102 348096 258023
rect 348056 250096 348108 250102
rect 348056 250038 348108 250044
rect 348056 241528 348108 241534
rect 348056 241470 348108 241476
rect 348068 230586 348096 241470
rect 347964 230580 348016 230586
rect 347964 230522 348016 230528
rect 348056 230580 348108 230586
rect 348056 230522 348108 230528
rect 347976 225010 348004 230522
rect 347964 225004 348016 225010
rect 347964 224946 348016 224952
rect 348056 224868 348108 224874
rect 348056 224810 348108 224816
rect 348068 217410 348096 224810
rect 348068 217382 348188 217410
rect 348160 212566 348188 217382
rect 347964 212560 348016 212566
rect 347964 212502 348016 212508
rect 348148 212560 348200 212566
rect 348148 212502 348200 212508
rect 347976 205698 348004 212502
rect 347964 205692 348016 205698
rect 347964 205634 348016 205640
rect 348056 205624 348108 205630
rect 348056 205566 348108 205572
rect 348068 198098 348096 205566
rect 348068 198070 348188 198098
rect 348160 193254 348188 198070
rect 347964 193248 348016 193254
rect 347964 193190 348016 193196
rect 348148 193248 348200 193254
rect 348148 193190 348200 193196
rect 347976 183598 348004 193190
rect 347964 183592 348016 183598
rect 347964 183534 348016 183540
rect 348056 183592 348108 183598
rect 348056 183534 348108 183540
rect 348068 180810 348096 183534
rect 348056 180804 348108 180810
rect 348056 180746 348108 180752
rect 347964 162920 348016 162926
rect 347964 162862 348016 162868
rect 347976 153218 348004 162862
rect 347976 153190 348096 153218
rect 348068 144906 348096 153190
rect 347964 144900 348016 144906
rect 347964 144842 348016 144848
rect 348056 144900 348108 144906
rect 348056 144842 348108 144848
rect 347976 134065 348004 144842
rect 347962 134056 348018 134065
rect 347962 133991 348018 134000
rect 347962 133920 348018 133929
rect 347962 133855 348018 133864
rect 347976 125662 348004 133855
rect 347964 125656 348016 125662
rect 347964 125598 348016 125604
rect 348056 125520 348108 125526
rect 348056 125462 348108 125468
rect 348068 114578 348096 125462
rect 348056 114572 348108 114578
rect 348056 114514 348108 114520
rect 348056 113212 348108 113218
rect 348056 113154 348108 113160
rect 348068 104922 348096 113154
rect 347872 104916 347924 104922
rect 347872 104858 347924 104864
rect 348056 104916 348108 104922
rect 348056 104858 348108 104864
rect 347884 85610 347912 104858
rect 347872 85604 347924 85610
rect 347872 85546 347924 85552
rect 348056 85604 348108 85610
rect 348056 85546 348108 85552
rect 348068 77382 348096 85546
rect 348056 77376 348108 77382
rect 348056 77318 348108 77324
rect 347964 77308 348016 77314
rect 347964 77250 348016 77256
rect 347976 60858 348004 77250
rect 347964 60852 348016 60858
rect 347964 60794 348016 60800
rect 347964 60716 348016 60722
rect 347964 60658 348016 60664
rect 347976 46986 348004 60658
rect 347964 46980 348016 46986
rect 347964 46922 348016 46928
rect 348148 46980 348200 46986
rect 348148 46922 348200 46928
rect 348160 35970 348188 46922
rect 347872 35964 347924 35970
rect 347872 35906 347924 35912
rect 348148 35964 348200 35970
rect 348148 35906 348200 35912
rect 347884 26246 347912 35906
rect 347872 26240 347924 26246
rect 347872 26182 347924 26188
rect 347964 19440 348016 19446
rect 347964 19382 348016 19388
rect 347976 12510 348004 19382
rect 347964 12504 348016 12510
rect 347964 12446 348016 12452
rect 347872 12436 347924 12442
rect 347872 12378 347924 12384
rect 347884 7614 347912 12378
rect 347872 7608 347924 7614
rect 347872 7550 347924 7556
rect 347964 7336 348016 7342
rect 347964 7278 348016 7284
rect 347780 4820 347832 4826
rect 347780 4762 347832 4768
rect 347872 4820 347924 4826
rect 347872 4762 347924 4768
rect 346676 4140 346728 4146
rect 346676 4082 346728 4088
rect 346492 3392 346544 3398
rect 346492 3334 346544 3340
rect 345480 740 345532 746
rect 345480 682 345532 688
rect 346308 740 346360 746
rect 346308 682 346360 688
rect 345492 480 345520 682
rect 346688 480 346716 4082
rect 347884 480 347912 4762
rect 347976 3330 348004 7278
rect 349068 6860 349120 6866
rect 349068 6802 349120 6808
rect 347964 3324 348016 3330
rect 347964 3266 348016 3272
rect 349080 480 349108 6802
rect 349172 4894 349200 335582
rect 349264 8430 349292 340054
rect 349632 335646 349660 340054
rect 349620 335640 349672 335646
rect 349620 335582 349672 335588
rect 350540 335640 350592 335646
rect 350540 335582 350592 335588
rect 349802 40488 349858 40497
rect 349802 40423 349858 40432
rect 349816 40225 349844 40423
rect 349802 40216 349858 40225
rect 349802 40151 349858 40160
rect 349252 8424 349304 8430
rect 349252 8366 349304 8372
rect 350552 4962 350580 335582
rect 350644 7682 350672 340068
rect 350736 340054 351210 340082
rect 351472 340054 351854 340082
rect 351932 340054 352498 340082
rect 352668 340054 353050 340082
rect 353312 340054 353694 340082
rect 353956 340054 354246 340082
rect 354784 340054 354890 340082
rect 355152 340054 355534 340082
rect 356086 340054 356192 340082
rect 350736 8362 350764 340054
rect 351472 335646 351500 340054
rect 351460 335640 351512 335646
rect 351460 335582 351512 335588
rect 351826 269104 351882 269113
rect 351826 269039 351882 269048
rect 351840 259486 351868 269039
rect 351828 259480 351880 259486
rect 351828 259422 351880 259428
rect 351826 240136 351882 240145
rect 351826 240071 351882 240080
rect 351840 234530 351868 240071
rect 351828 234524 351880 234530
rect 351828 234466 351880 234472
rect 351826 230480 351882 230489
rect 351826 230415 351882 230424
rect 351840 220862 351868 230415
rect 351828 220856 351880 220862
rect 351828 220798 351880 220804
rect 351828 211132 351880 211138
rect 351828 211074 351880 211080
rect 351840 201521 351868 211074
rect 351826 201512 351882 201521
rect 351826 201447 351882 201456
rect 351826 104816 351882 104825
rect 351826 104751 351882 104760
rect 351840 95130 351868 104751
rect 351828 95124 351880 95130
rect 351828 95066 351880 95072
rect 350998 29472 351054 29481
rect 350998 29407 351054 29416
rect 351012 29209 351040 29407
rect 350998 29200 351054 29209
rect 350998 29135 351054 29144
rect 350724 8356 350776 8362
rect 350724 8298 350776 8304
rect 350632 7676 350684 7682
rect 350632 7618 350684 7624
rect 351828 7608 351880 7614
rect 351828 7550 351880 7556
rect 350540 4956 350592 4962
rect 350540 4898 350592 4904
rect 349160 4888 349212 4894
rect 349160 4830 349212 4836
rect 351368 4888 351420 4894
rect 351368 4830 351420 4836
rect 350264 3052 350316 3058
rect 350264 2994 350316 3000
rect 350276 480 350304 2994
rect 351380 480 351408 4830
rect 351840 2990 351868 7550
rect 351932 7070 351960 340054
rect 352668 333334 352696 340054
rect 353208 337136 353260 337142
rect 353208 337078 353260 337084
rect 352012 333328 352064 333334
rect 352012 333270 352064 333276
rect 352656 333328 352708 333334
rect 352656 333270 352708 333276
rect 352024 328522 352052 333270
rect 352024 328494 352144 328522
rect 352116 325689 352144 328494
rect 352102 325680 352158 325689
rect 352102 325615 352158 325624
rect 352286 325680 352342 325689
rect 352286 325615 352342 325624
rect 352300 316062 352328 325615
rect 352104 316056 352156 316062
rect 352102 316024 352104 316033
rect 352288 316056 352340 316062
rect 352156 316024 352158 316033
rect 352102 315959 352158 315968
rect 352286 316024 352288 316033
rect 352340 316024 352342 316033
rect 352286 315959 352342 315968
rect 352300 306406 352328 315959
rect 352104 306400 352156 306406
rect 352104 306342 352156 306348
rect 352288 306400 352340 306406
rect 352288 306342 352340 306348
rect 352116 298110 352144 306342
rect 352104 298104 352156 298110
rect 352104 298046 352156 298052
rect 352104 287972 352156 287978
rect 352104 287914 352156 287920
rect 352116 287065 352144 287914
rect 352102 287056 352158 287065
rect 352102 286991 352158 287000
rect 352286 287056 352342 287065
rect 352286 286991 352342 287000
rect 352300 280158 352328 286991
rect 352104 280152 352156 280158
rect 352104 280094 352156 280100
rect 352288 280152 352340 280158
rect 352288 280094 352340 280100
rect 352116 269113 352144 280094
rect 352102 269104 352158 269113
rect 352102 269039 352158 269048
rect 352012 259480 352064 259486
rect 352012 259422 352064 259428
rect 352024 251258 352052 259422
rect 352012 251252 352064 251258
rect 352012 251194 352064 251200
rect 352104 251252 352156 251258
rect 352104 251194 352156 251200
rect 352116 246378 352144 251194
rect 352024 246350 352144 246378
rect 352024 240145 352052 246350
rect 352010 240136 352066 240145
rect 352010 240071 352066 240080
rect 352104 234524 352156 234530
rect 352104 234466 352156 234472
rect 352116 230489 352144 234466
rect 352102 230480 352158 230489
rect 352102 230415 352158 230424
rect 352012 220856 352064 220862
rect 352012 220798 352064 220804
rect 352024 212566 352052 220798
rect 352012 212560 352064 212566
rect 352104 212560 352156 212566
rect 352064 212508 352104 212514
rect 352012 212502 352156 212508
rect 352024 212486 352144 212502
rect 352024 211138 352052 212486
rect 352012 211132 352064 211138
rect 352012 211074 352064 211080
rect 352102 201512 352158 201521
rect 352102 201447 352104 201456
rect 352156 201447 352158 201456
rect 352104 201418 352156 201424
rect 352104 193180 352156 193186
rect 352104 193122 352156 193128
rect 352116 191842 352144 193122
rect 352116 191814 352236 191842
rect 352208 183598 352236 191814
rect 352012 183592 352064 183598
rect 352012 183534 352064 183540
rect 352196 183592 352248 183598
rect 352196 183534 352248 183540
rect 352024 180810 352052 183534
rect 352012 180804 352064 180810
rect 352012 180746 352064 180752
rect 352104 162920 352156 162926
rect 352104 162862 352156 162868
rect 352116 153218 352144 162862
rect 352024 153190 352144 153218
rect 352024 144906 352052 153190
rect 352012 144900 352064 144906
rect 352012 144842 352064 144848
rect 352196 144900 352248 144906
rect 352196 144842 352248 144848
rect 352208 137714 352236 144842
rect 352116 137686 352236 137714
rect 352116 125769 352144 137686
rect 352102 125760 352158 125769
rect 352102 125695 352158 125704
rect 352010 125624 352066 125633
rect 352010 125559 352066 125568
rect 352024 119354 352052 125559
rect 352024 119326 352144 119354
rect 352116 109698 352144 119326
rect 352024 109670 352144 109698
rect 352024 104825 352052 109670
rect 352010 104816 352066 104825
rect 352010 104751 352066 104760
rect 352196 95124 352248 95130
rect 352196 95066 352248 95072
rect 352208 85610 352236 95066
rect 352104 85604 352156 85610
rect 352104 85546 352156 85552
rect 352196 85604 352248 85610
rect 352196 85546 352248 85552
rect 352116 77382 352144 85546
rect 352104 77376 352156 77382
rect 352104 77318 352156 77324
rect 352012 66292 352064 66298
rect 352012 66234 352064 66240
rect 352024 66178 352052 66234
rect 352024 66150 352144 66178
rect 352116 48414 352144 66150
rect 352104 48408 352156 48414
rect 352104 48350 352156 48356
rect 352012 48340 352064 48346
rect 352012 48282 352064 48288
rect 352024 37330 352052 48282
rect 352012 37324 352064 37330
rect 352012 37266 352064 37272
rect 352104 37324 352156 37330
rect 352104 37266 352156 37272
rect 352116 37210 352144 37266
rect 352116 37182 352328 37210
rect 352300 19258 352328 37182
rect 352208 19230 352328 19258
rect 352208 14074 352236 19230
rect 352196 14068 352248 14074
rect 352196 14010 352248 14016
rect 351920 7064 351972 7070
rect 351920 7006 351972 7012
rect 353220 3738 353248 337078
rect 353312 5030 353340 340054
rect 353956 328506 353984 340054
rect 354680 335640 354732 335646
rect 354680 335582 354732 335588
rect 353576 328500 353628 328506
rect 353576 328442 353628 328448
rect 353944 328500 353996 328506
rect 353944 328442 353996 328448
rect 353588 309194 353616 328442
rect 353484 309188 353536 309194
rect 353484 309130 353536 309136
rect 353576 309188 353628 309194
rect 353576 309130 353628 309136
rect 353496 299606 353524 309130
rect 353484 299600 353536 299606
rect 353484 299542 353536 299548
rect 353484 299396 353536 299402
rect 353484 299338 353536 299344
rect 353496 298110 353524 299338
rect 353484 298104 353536 298110
rect 353484 298046 353536 298052
rect 353576 298104 353628 298110
rect 353576 298046 353628 298052
rect 353588 280158 353616 298046
rect 353484 280152 353536 280158
rect 353484 280094 353536 280100
rect 353576 280152 353628 280158
rect 353576 280094 353628 280100
rect 353496 263634 353524 280094
rect 353484 263628 353536 263634
rect 353484 263570 353536 263576
rect 353576 263492 353628 263498
rect 353576 263434 353628 263440
rect 353588 251190 353616 263434
rect 353576 251184 353628 251190
rect 353576 251126 353628 251132
rect 353576 241528 353628 241534
rect 353576 241470 353628 241476
rect 353588 230586 353616 241470
rect 353484 230580 353536 230586
rect 353484 230522 353536 230528
rect 353576 230580 353628 230586
rect 353576 230522 353628 230528
rect 353496 225010 353524 230522
rect 353484 225004 353536 225010
rect 353484 224946 353536 224952
rect 353576 224868 353628 224874
rect 353576 224810 353628 224816
rect 353588 217410 353616 224810
rect 353588 217382 353708 217410
rect 353680 212566 353708 217382
rect 353484 212560 353536 212566
rect 353668 212560 353720 212566
rect 353536 212508 353616 212514
rect 353484 212502 353616 212508
rect 353668 212502 353720 212508
rect 353496 212486 353616 212502
rect 353588 198098 353616 212486
rect 353588 198070 353708 198098
rect 353680 193254 353708 198070
rect 353484 193248 353536 193254
rect 353484 193190 353536 193196
rect 353668 193248 353720 193254
rect 353668 193190 353720 193196
rect 353496 183598 353524 193190
rect 353484 183592 353536 183598
rect 353484 183534 353536 183540
rect 353576 183592 353628 183598
rect 353576 183534 353628 183540
rect 353588 180810 353616 183534
rect 353576 180804 353628 180810
rect 353576 180746 353628 180752
rect 353484 162920 353536 162926
rect 353484 162862 353536 162868
rect 353496 153218 353524 162862
rect 353496 153190 353616 153218
rect 353588 144906 353616 153190
rect 353484 144900 353536 144906
rect 353484 144842 353536 144848
rect 353576 144900 353628 144906
rect 353576 144842 353628 144848
rect 353496 134065 353524 144842
rect 353482 134056 353538 134065
rect 353482 133991 353538 134000
rect 353482 133920 353538 133929
rect 353482 133855 353484 133864
rect 353536 133855 353538 133864
rect 353484 133826 353536 133832
rect 353576 124228 353628 124234
rect 353576 124170 353628 124176
rect 353588 114646 353616 124170
rect 354588 123276 354640 123282
rect 354588 123218 354640 123224
rect 354600 123185 354628 123218
rect 354586 123176 354642 123185
rect 354586 123111 354642 123120
rect 353576 114640 353628 114646
rect 353576 114582 353628 114588
rect 353484 114572 353536 114578
rect 353484 114514 353536 114520
rect 353496 114481 353524 114514
rect 353482 114472 353538 114481
rect 353482 114407 353538 114416
rect 353574 114336 353630 114345
rect 353574 114271 353630 114280
rect 353588 103494 353616 114271
rect 353576 103488 353628 103494
rect 353576 103430 353628 103436
rect 353484 93900 353536 93906
rect 353484 93842 353536 93848
rect 353496 84182 353524 93842
rect 354586 87272 354642 87281
rect 354586 87207 354642 87216
rect 354600 87174 354628 87207
rect 354588 87168 354640 87174
rect 354588 87110 354640 87116
rect 353484 84176 353536 84182
rect 353484 84118 353536 84124
rect 353392 84108 353444 84114
rect 353392 84050 353444 84056
rect 353404 66337 353432 84050
rect 353390 66328 353446 66337
rect 353390 66263 353446 66272
rect 353666 66056 353722 66065
rect 353666 65991 353722 66000
rect 353680 56574 353708 65991
rect 353484 56568 353536 56574
rect 353484 56510 353536 56516
rect 353668 56568 353720 56574
rect 353668 56510 353720 56516
rect 353496 47002 353524 56510
rect 353496 46974 353616 47002
rect 353588 45558 353616 46974
rect 353576 45552 353628 45558
rect 353576 45494 353628 45500
rect 353576 37256 353628 37262
rect 353576 37198 353628 37204
rect 353588 32450 353616 37198
rect 353588 32422 353708 32450
rect 353680 12186 353708 32422
rect 353404 12158 353708 12186
rect 353404 7002 353432 12158
rect 353392 6996 353444 7002
rect 353392 6938 353444 6944
rect 354692 5098 354720 335582
rect 354784 14482 354812 340054
rect 355152 335646 355180 340054
rect 355140 335640 355192 335646
rect 355140 335582 355192 335588
rect 355506 63880 355562 63889
rect 355506 63815 355508 63824
rect 355560 63815 355562 63824
rect 355508 63786 355560 63792
rect 355966 17232 356022 17241
rect 355966 17167 356022 17176
rect 355980 16862 356008 17167
rect 355968 16856 356020 16862
rect 355968 16798 356020 16804
rect 354772 14476 354824 14482
rect 354772 14418 354824 14424
rect 356164 7750 356192 340054
rect 356256 340054 356730 340082
rect 356256 9926 356284 340054
rect 357360 338434 357388 340068
rect 357452 340054 357926 340082
rect 358280 340054 358570 340082
rect 358832 340054 359214 340082
rect 359476 340054 359766 340082
rect 360304 340054 360410 340082
rect 360672 340054 361054 340082
rect 356704 338428 356756 338434
rect 356704 338370 356756 338376
rect 357348 338428 357400 338434
rect 357348 338370 357400 338376
rect 356716 336734 356744 338370
rect 357348 337136 357400 337142
rect 357348 337078 357400 337084
rect 356520 336728 356572 336734
rect 356520 336670 356572 336676
rect 356704 336728 356756 336734
rect 356704 336670 356756 336676
rect 356532 335306 356560 336670
rect 356520 335300 356572 335306
rect 356520 335242 356572 335248
rect 356520 317484 356572 317490
rect 356520 317426 356572 317432
rect 356532 304314 356560 317426
rect 356532 304286 356652 304314
rect 356624 289898 356652 304286
rect 356440 289870 356652 289898
rect 356440 289814 356468 289870
rect 356428 289808 356480 289814
rect 356428 289750 356480 289756
rect 356520 289740 356572 289746
rect 356520 289682 356572 289688
rect 356532 288425 356560 289682
rect 356518 288416 356574 288425
rect 356518 288351 356574 288360
rect 356702 288416 356758 288425
rect 356702 288351 356758 288360
rect 356716 277438 356744 288351
rect 356428 277432 356480 277438
rect 356428 277374 356480 277380
rect 356704 277432 356756 277438
rect 356704 277374 356756 277380
rect 356440 273358 356468 277374
rect 356428 273352 356480 273358
rect 356428 273294 356480 273300
rect 356428 270496 356480 270502
rect 356428 270438 356480 270444
rect 356440 263702 356468 270438
rect 356428 263696 356480 263702
rect 356428 263638 356480 263644
rect 356520 263560 356572 263566
rect 356520 263502 356572 263508
rect 356532 259570 356560 263502
rect 356440 259542 356560 259570
rect 356440 258058 356468 259542
rect 356428 258052 356480 258058
rect 356428 257994 356480 258000
rect 356612 258052 356664 258058
rect 356612 257994 356664 258000
rect 356624 248441 356652 257994
rect 356426 248432 356482 248441
rect 356336 248396 356388 248402
rect 356426 248367 356428 248376
rect 356336 248338 356388 248344
rect 356480 248367 356482 248376
rect 356610 248432 356666 248441
rect 356610 248367 356666 248376
rect 356428 248338 356480 248344
rect 356348 238785 356376 248338
rect 356334 238776 356390 238785
rect 356334 238711 356390 238720
rect 356518 238776 356574 238785
rect 356518 238711 356574 238720
rect 356532 238678 356560 238711
rect 356520 238672 356572 238678
rect 356520 238614 356572 238620
rect 356612 238672 356664 238678
rect 356612 238614 356664 238620
rect 356624 233866 356652 238614
rect 356532 233838 356652 233866
rect 356532 212634 356560 233838
rect 356520 212628 356572 212634
rect 356520 212570 356572 212576
rect 356428 212560 356480 212566
rect 356426 212528 356428 212537
rect 356480 212528 356482 212537
rect 356426 212463 356482 212472
rect 356610 212528 356666 212537
rect 356610 212463 356666 212472
rect 356624 204898 356652 212463
rect 356440 204870 356652 204898
rect 356440 202722 356468 204870
rect 356440 202694 356560 202722
rect 356532 193322 356560 202694
rect 356520 193316 356572 193322
rect 356520 193258 356572 193264
rect 356428 193248 356480 193254
rect 356428 193190 356480 193196
rect 356440 183598 356468 193190
rect 356428 183592 356480 183598
rect 356428 183534 356480 183540
rect 356520 183592 356572 183598
rect 356520 183534 356572 183540
rect 356532 167142 356560 183534
rect 356520 167136 356572 167142
rect 356520 167078 356572 167084
rect 356428 166932 356480 166938
rect 356428 166874 356480 166880
rect 356440 161362 356468 166874
rect 356428 161356 356480 161362
rect 356428 161298 356480 161304
rect 356428 151836 356480 151842
rect 356428 151778 356480 151784
rect 356440 144945 356468 151778
rect 356426 144936 356482 144945
rect 356426 144871 356482 144880
rect 356426 144800 356482 144809
rect 356426 144735 356482 144744
rect 356440 134065 356468 144735
rect 356426 134056 356482 134065
rect 356426 133991 356482 134000
rect 356426 133920 356482 133929
rect 356426 133855 356428 133864
rect 356480 133855 356482 133864
rect 356428 133826 356480 133832
rect 356428 124228 356480 124234
rect 356428 124170 356480 124176
rect 356440 114646 356468 124170
rect 356428 114640 356480 114646
rect 356428 114582 356480 114588
rect 356520 114572 356572 114578
rect 356520 114514 356572 114520
rect 356532 104802 356560 114514
rect 356532 104774 356652 104802
rect 356624 103494 356652 104774
rect 356612 103488 356664 103494
rect 356612 103430 356664 103436
rect 356428 103420 356480 103426
rect 356428 103362 356480 103368
rect 356440 94081 356468 103362
rect 356426 94072 356482 94081
rect 356426 94007 356482 94016
rect 356426 93936 356482 93945
rect 356426 93871 356482 93880
rect 356440 89758 356468 93871
rect 356428 89752 356480 89758
rect 356428 89694 356480 89700
rect 356520 89616 356572 89622
rect 356520 89558 356572 89564
rect 356532 84182 356560 89558
rect 356520 84176 356572 84182
rect 356520 84118 356572 84124
rect 356520 84040 356572 84046
rect 356520 83982 356572 83988
rect 356532 82822 356560 83982
rect 356520 82816 356572 82822
rect 356520 82758 356572 82764
rect 356428 73228 356480 73234
rect 356428 73170 356480 73176
rect 356440 64870 356468 73170
rect 356428 64864 356480 64870
rect 356428 64806 356480 64812
rect 356612 64864 356664 64870
rect 356612 64806 356664 64812
rect 356624 63510 356652 64806
rect 356612 63504 356664 63510
rect 356612 63446 356664 63452
rect 356520 45620 356572 45626
rect 356520 45562 356572 45568
rect 356532 40798 356560 45562
rect 356520 40792 356572 40798
rect 356520 40734 356572 40740
rect 356612 35964 356664 35970
rect 356612 35906 356664 35912
rect 356624 31142 356652 35906
rect 356612 31136 356664 31142
rect 356612 31078 356664 31084
rect 356520 26376 356572 26382
rect 356520 26318 356572 26324
rect 356532 24857 356560 26318
rect 356334 24848 356390 24857
rect 356334 24783 356390 24792
rect 356518 24848 356574 24857
rect 356518 24783 356574 24792
rect 356348 15230 356376 24783
rect 356336 15224 356388 15230
rect 356336 15166 356388 15172
rect 356428 15224 356480 15230
rect 356428 15166 356480 15172
rect 356244 9920 356296 9926
rect 356244 9862 356296 9868
rect 356152 7744 356204 7750
rect 356152 7686 356204 7692
rect 354956 6044 355008 6050
rect 354956 5986 355008 5992
rect 354680 5092 354732 5098
rect 354680 5034 354732 5040
rect 353300 5024 353352 5030
rect 353300 4966 353352 4972
rect 352564 3732 352616 3738
rect 352564 3674 352616 3680
rect 353208 3732 353260 3738
rect 353208 3674 353260 3680
rect 351828 2984 351880 2990
rect 351828 2926 351880 2932
rect 352576 480 352604 3674
rect 353760 3392 353812 3398
rect 353760 3334 353812 3340
rect 353772 480 353800 3334
rect 354968 480 354996 5986
rect 356440 5166 356468 15166
rect 356428 5160 356480 5166
rect 356428 5102 356480 5108
rect 356060 4616 356112 4622
rect 356060 4558 356112 4564
rect 356072 3466 356100 4558
rect 356060 3460 356112 3466
rect 356060 3402 356112 3408
rect 356150 3360 356206 3369
rect 356150 3295 356206 3304
rect 356164 480 356192 3295
rect 357360 480 357388 337078
rect 357452 7818 357480 340054
rect 358280 335646 358308 340054
rect 357624 335640 357676 335646
rect 357624 335582 357676 335588
rect 358268 335640 358320 335646
rect 358268 335582 358320 335588
rect 357636 327078 357664 335582
rect 357624 327072 357676 327078
rect 357624 327014 357676 327020
rect 357532 317484 357584 317490
rect 357532 317426 357584 317432
rect 357544 316033 357572 317426
rect 357530 316024 357586 316033
rect 357530 315959 357586 315968
rect 357714 316024 357770 316033
rect 357714 315959 357770 315968
rect 357728 306406 357756 315959
rect 357532 306400 357584 306406
rect 357532 306342 357584 306348
rect 357716 306400 357768 306406
rect 357716 306342 357768 306348
rect 357544 299282 357572 306342
rect 357544 299254 357664 299282
rect 357636 298058 357664 299254
rect 357544 298030 357664 298058
rect 357544 296721 357572 298030
rect 357530 296712 357586 296721
rect 357530 296647 357586 296656
rect 357806 296712 357862 296721
rect 357806 296647 357862 296656
rect 357820 278798 357848 296647
rect 357624 278792 357676 278798
rect 357624 278734 357676 278740
rect 357808 278792 357860 278798
rect 357808 278734 357860 278740
rect 357636 273358 357664 278734
rect 357624 273352 357676 273358
rect 357624 273294 357676 273300
rect 357624 273216 357676 273222
rect 357624 273158 357676 273164
rect 357636 253994 357664 273158
rect 357544 253966 357664 253994
rect 357544 253858 357572 253966
rect 357544 253830 357664 253858
rect 357636 241482 357664 253830
rect 357636 241454 357756 241482
rect 357728 234666 357756 241454
rect 357716 234660 357768 234666
rect 357716 234602 357768 234608
rect 357624 234592 357676 234598
rect 357624 234534 357676 234540
rect 357636 222170 357664 234534
rect 357636 222142 357756 222170
rect 357728 215354 357756 222142
rect 357716 215348 357768 215354
rect 357716 215290 357768 215296
rect 357624 215280 357676 215286
rect 357624 215222 357676 215228
rect 357636 196058 357664 215222
rect 357544 196030 357664 196058
rect 357544 195922 357572 196030
rect 357544 195894 357664 195922
rect 357636 186454 357664 195894
rect 357624 186448 357676 186454
rect 357624 186390 357676 186396
rect 357624 179444 357676 179450
rect 357624 179386 357676 179392
rect 357636 179330 357664 179386
rect 357636 179302 357756 179330
rect 357728 144945 357756 179302
rect 357530 144936 357586 144945
rect 357530 144871 357532 144880
rect 357584 144871 357586 144880
rect 357714 144936 357770 144945
rect 357714 144871 357716 144880
rect 357532 144842 357584 144848
rect 357768 144871 357770 144880
rect 357716 144842 357768 144848
rect 357728 137714 357756 144842
rect 357636 137686 357756 137714
rect 357636 125769 357664 137686
rect 357622 125760 357678 125769
rect 357622 125695 357678 125704
rect 357622 125624 357678 125633
rect 357622 125559 357678 125568
rect 357636 118794 357664 125559
rect 357624 118788 357676 118794
rect 357624 118730 357676 118736
rect 357624 118652 357676 118658
rect 357624 118594 357676 118600
rect 357636 106282 357664 118594
rect 357624 106276 357676 106282
rect 357624 106218 357676 106224
rect 357716 96552 357768 96558
rect 357716 96494 357768 96500
rect 357728 87009 357756 96494
rect 357530 87000 357586 87009
rect 357530 86935 357586 86944
rect 357714 87000 357770 87009
rect 357714 86935 357770 86944
rect 357544 86902 357572 86935
rect 357532 86896 357584 86902
rect 357532 86838 357584 86844
rect 357716 86896 357768 86902
rect 357716 86838 357768 86844
rect 357728 84182 357756 86838
rect 357716 84176 357768 84182
rect 357716 84118 357768 84124
rect 357716 74588 357768 74594
rect 357716 74530 357768 74536
rect 357728 64938 357756 74530
rect 357624 64932 357676 64938
rect 357624 64874 357676 64880
rect 357716 64932 357768 64938
rect 357716 64874 357768 64880
rect 357636 41478 357664 64874
rect 357624 41472 357676 41478
rect 357624 41414 357676 41420
rect 357532 35964 357584 35970
rect 357532 35906 357584 35912
rect 357544 26246 357572 35906
rect 357532 26240 357584 26246
rect 357532 26182 357584 26188
rect 357440 7812 357492 7818
rect 357440 7754 357492 7760
rect 358832 5234 358860 340054
rect 359476 328506 359504 340054
rect 360108 337068 360160 337074
rect 360108 337010 360160 337016
rect 359096 328500 359148 328506
rect 359096 328442 359148 328448
rect 359464 328500 359516 328506
rect 359464 328442 359516 328448
rect 359108 321638 359136 328442
rect 359096 321632 359148 321638
rect 359096 321574 359148 321580
rect 359004 321564 359056 321570
rect 359004 321506 359056 321512
rect 359016 318730 359044 321506
rect 359016 318702 359136 318730
rect 359108 292618 359136 318702
rect 359016 292590 359136 292618
rect 359016 282826 359044 292590
rect 359016 282798 359136 282826
rect 359108 280158 359136 282798
rect 359004 280152 359056 280158
rect 359004 280094 359056 280100
rect 359096 280152 359148 280158
rect 359096 280094 359148 280100
rect 359016 270745 359044 280094
rect 359002 270736 359058 270745
rect 359002 270671 359058 270680
rect 359186 270464 359242 270473
rect 359186 270399 359242 270408
rect 359200 260914 359228 270399
rect 359096 260908 359148 260914
rect 359096 260850 359148 260856
rect 359188 260908 359240 260914
rect 359188 260850 359240 260856
rect 359108 249966 359136 260850
rect 359096 249960 359148 249966
rect 359096 249902 359148 249908
rect 359004 249892 359056 249898
rect 359004 249834 359056 249840
rect 359016 249801 359044 249834
rect 359002 249792 359058 249801
rect 359002 249727 359058 249736
rect 359278 249792 359334 249801
rect 359278 249727 359334 249736
rect 359292 240174 359320 249727
rect 359096 240168 359148 240174
rect 359096 240110 359148 240116
rect 359280 240168 359332 240174
rect 359280 240110 359332 240116
rect 359108 233918 359136 240110
rect 359096 233912 359148 233918
rect 359096 233854 359148 233860
rect 359280 233912 359332 233918
rect 359280 233854 359332 233860
rect 359292 229129 359320 233854
rect 359094 229120 359150 229129
rect 359094 229055 359150 229064
rect 359278 229120 359334 229129
rect 359278 229055 359334 229064
rect 359108 220862 359136 229055
rect 358912 220856 358964 220862
rect 358912 220798 358964 220804
rect 359096 220856 359148 220862
rect 359096 220798 359148 220804
rect 358924 218006 358952 220798
rect 358912 218000 358964 218006
rect 358912 217942 358964 217948
rect 359004 218000 359056 218006
rect 359004 217942 359056 217948
rect 359016 209658 359044 217942
rect 359016 209630 359228 209658
rect 359200 200297 359228 209630
rect 359186 200288 359242 200297
rect 359186 200223 359242 200232
rect 359094 198792 359150 198801
rect 359094 198727 359150 198736
rect 359108 197334 359136 198727
rect 359096 197328 359148 197334
rect 359096 197270 359148 197276
rect 359096 187740 359148 187746
rect 359096 187682 359148 187688
rect 359108 179314 359136 187682
rect 359096 179308 359148 179314
rect 359096 179250 359148 179256
rect 359188 179308 359240 179314
rect 359188 179250 359240 179256
rect 359200 144945 359228 179250
rect 359002 144936 359058 144945
rect 359002 144871 359004 144880
rect 359056 144871 359058 144880
rect 359186 144936 359242 144945
rect 359186 144871 359188 144880
rect 359004 144842 359056 144848
rect 359240 144871 359242 144880
rect 359188 144842 359240 144848
rect 359200 139890 359228 144842
rect 359108 139862 359228 139890
rect 359108 124273 359136 139862
rect 359094 124264 359150 124273
rect 359094 124199 359150 124208
rect 359186 114472 359242 114481
rect 359186 114407 359242 114416
rect 359200 89690 359228 114407
rect 359004 89684 359056 89690
rect 359004 89626 359056 89632
rect 359188 89684 359240 89690
rect 359188 89626 359240 89632
rect 359016 84182 359044 89626
rect 359004 84176 359056 84182
rect 359004 84118 359056 84124
rect 359280 77988 359332 77994
rect 359280 77930 359332 77936
rect 359292 73166 359320 77930
rect 359188 73160 359240 73166
rect 359188 73102 359240 73108
rect 359280 73160 359332 73166
rect 359280 73102 359332 73108
rect 359200 63510 359228 73102
rect 359188 63504 359240 63510
rect 359188 63446 359240 63452
rect 359188 53848 359240 53854
rect 359188 53790 359240 53796
rect 359200 48414 359228 53790
rect 359188 48408 359240 48414
rect 359188 48350 359240 48356
rect 359096 45620 359148 45626
rect 359096 45562 359148 45568
rect 359108 35902 359136 45562
rect 358912 35896 358964 35902
rect 358912 35838 358964 35844
rect 359096 35896 359148 35902
rect 359096 35838 359148 35844
rect 358924 26246 358952 35838
rect 358912 26240 358964 26246
rect 358912 26182 358964 26188
rect 359004 26172 359056 26178
rect 359004 26114 359056 26120
rect 359016 8362 359044 26114
rect 358912 8356 358964 8362
rect 358912 8298 358964 8304
rect 359004 8356 359056 8362
rect 359004 8298 359056 8304
rect 358924 7886 358952 8298
rect 358912 7880 358964 7886
rect 358912 7822 358964 7828
rect 358820 5228 358872 5234
rect 358820 5170 358872 5176
rect 358544 4956 358596 4962
rect 358544 4898 358596 4904
rect 358556 480 358584 4898
rect 360120 626 360148 337010
rect 360200 335640 360252 335646
rect 360200 335582 360252 335588
rect 360212 5914 360240 335582
rect 360304 9790 360332 340054
rect 360672 335646 360700 340054
rect 360660 335640 360712 335646
rect 360660 335582 360712 335588
rect 360384 63844 360436 63850
rect 360384 63786 360436 63792
rect 360396 63617 360424 63786
rect 360382 63608 360438 63617
rect 360382 63543 360438 63552
rect 360292 9784 360344 9790
rect 360292 9726 360344 9732
rect 361592 7954 361620 340068
rect 361776 340054 362250 340082
rect 362512 340054 362894 340082
rect 363064 340054 363446 340082
rect 363800 340054 364090 340082
rect 364352 340054 364734 340082
rect 361672 335640 361724 335646
rect 361672 335582 361724 335588
rect 361684 9314 361712 335582
rect 361776 9722 361804 340054
rect 362512 335646 362540 340054
rect 362500 335640 362552 335646
rect 362500 335582 362552 335588
rect 362960 335640 363012 335646
rect 362960 335582 363012 335588
rect 361764 9716 361816 9722
rect 361764 9658 361816 9664
rect 361672 9308 361724 9314
rect 361672 9250 361724 9256
rect 361580 7948 361632 7954
rect 361580 7890 361632 7896
rect 360200 5908 360252 5914
rect 360200 5850 360252 5856
rect 362132 5908 362184 5914
rect 362132 5850 362184 5856
rect 360936 3324 360988 3330
rect 360936 3266 360988 3272
rect 359752 598 360148 626
rect 359752 480 359780 598
rect 360948 480 360976 3266
rect 362144 480 362172 5850
rect 362972 4622 363000 335582
rect 363064 8022 363092 340054
rect 363604 336864 363656 336870
rect 363604 336806 363656 336812
rect 363052 8016 363104 8022
rect 363052 7958 363104 7964
rect 362960 4616 363012 4622
rect 362960 4558 363012 4564
rect 363616 3262 363644 336806
rect 363696 336796 363748 336802
rect 363696 336738 363748 336744
rect 363708 4010 363736 336738
rect 363800 335646 363828 340054
rect 363788 335640 363840 335646
rect 363788 335582 363840 335588
rect 364352 212838 364380 340054
rect 364812 328506 364840 340190
rect 365916 337686 365944 340068
rect 366008 340054 366574 340082
rect 365904 337680 365956 337686
rect 365904 337622 365956 337628
rect 366008 328522 366036 340054
rect 366916 337680 366968 337686
rect 366916 337622 366968 337628
rect 366456 337000 366508 337006
rect 366456 336942 366508 336948
rect 366364 336932 366416 336938
rect 366364 336874 366416 336880
rect 364616 328500 364668 328506
rect 364616 328442 364668 328448
rect 364800 328500 364852 328506
rect 364800 328442 364852 328448
rect 365916 328494 366036 328522
rect 364628 309194 364656 328442
rect 365916 318782 365944 328494
rect 365812 318776 365864 318782
rect 365812 318718 365864 318724
rect 365904 318776 365956 318782
rect 365904 318718 365956 318724
rect 365824 317422 365852 318718
rect 365812 317416 365864 317422
rect 365812 317358 365864 317364
rect 365904 317416 365956 317422
rect 365904 317358 365956 317364
rect 364524 309188 364576 309194
rect 364524 309130 364576 309136
rect 364616 309188 364668 309194
rect 364616 309130 364668 309136
rect 364536 307766 364564 309130
rect 364524 307760 364576 307766
rect 364524 307702 364576 307708
rect 364616 298172 364668 298178
rect 364616 298114 364668 298120
rect 364628 298058 364656 298114
rect 364536 298030 364656 298058
rect 364536 291378 364564 298030
rect 365916 292618 365944 317358
rect 365824 292590 365944 292618
rect 365824 292482 365852 292590
rect 365824 292454 365944 292482
rect 364524 291372 364576 291378
rect 364524 291314 364576 291320
rect 364616 284980 364668 284986
rect 364616 284922 364668 284928
rect 364628 280158 364656 284922
rect 365916 280158 365944 292454
rect 364524 280152 364576 280158
rect 364524 280094 364576 280100
rect 364616 280152 364668 280158
rect 364616 280094 364668 280100
rect 365904 280152 365956 280158
rect 365904 280094 365956 280100
rect 365996 280152 366048 280158
rect 365996 280094 366048 280100
rect 364536 270745 364564 280094
rect 366008 273204 366036 280094
rect 365916 273176 366036 273204
rect 364522 270736 364578 270745
rect 364522 270671 364578 270680
rect 364614 270464 364670 270473
rect 364614 270399 364670 270408
rect 364628 249898 364656 270399
rect 365916 253994 365944 273176
rect 365824 253966 365944 253994
rect 365824 253858 365852 253966
rect 365824 253830 365944 253858
rect 364524 249892 364576 249898
rect 364524 249834 364576 249840
rect 364616 249892 364668 249898
rect 364616 249834 364668 249840
rect 364536 244322 364564 249834
rect 364524 244316 364576 244322
rect 364524 244258 364576 244264
rect 364616 244180 364668 244186
rect 364616 244122 364668 244128
rect 364628 231878 364656 244122
rect 364616 231872 364668 231878
rect 364616 231814 364668 231820
rect 364524 231804 364576 231810
rect 364524 231746 364576 231752
rect 364536 229106 364564 231746
rect 364536 229078 364748 229106
rect 364720 220862 364748 229078
rect 364432 220856 364484 220862
rect 364432 220798 364484 220804
rect 364708 220856 364760 220862
rect 364708 220798 364760 220804
rect 364340 212832 364392 212838
rect 364340 212774 364392 212780
rect 364444 212566 364472 220798
rect 364432 212560 364484 212566
rect 364432 212502 364484 212508
rect 364340 212424 364392 212430
rect 364340 212366 364392 212372
rect 364156 208412 364208 208418
rect 364156 208354 364208 208360
rect 364168 202910 364196 208354
rect 364156 202904 364208 202910
rect 364156 202846 364208 202852
rect 364352 181082 364380 212366
rect 364616 202904 364668 202910
rect 364616 202846 364668 202852
rect 364628 196110 364656 202846
rect 365916 196654 365944 253830
rect 365720 196648 365772 196654
rect 365720 196590 365772 196596
rect 365904 196648 365956 196654
rect 365904 196590 365956 196596
rect 364616 196104 364668 196110
rect 364616 196046 364668 196052
rect 364800 196104 364852 196110
rect 364800 196046 364852 196052
rect 364812 190505 364840 196046
rect 365732 191865 365760 196590
rect 365718 191856 365774 191865
rect 365718 191791 365774 191800
rect 365902 191856 365958 191865
rect 365902 191791 365958 191800
rect 364614 190496 364670 190505
rect 364536 190466 364614 190482
rect 364524 190460 364614 190466
rect 364576 190454 364614 190460
rect 364614 190431 364670 190440
rect 364798 190496 364854 190505
rect 364798 190431 364854 190440
rect 364524 190402 364576 190408
rect 364536 190371 364564 190402
rect 364524 186312 364576 186318
rect 364524 186254 364576 186260
rect 364340 181076 364392 181082
rect 364340 181018 364392 181024
rect 364340 180872 364392 180878
rect 364340 180814 364392 180820
rect 364536 180826 364564 186254
rect 365916 182170 365944 191791
rect 365720 182164 365772 182170
rect 365720 182106 365772 182112
rect 365904 182164 365956 182170
rect 365904 182106 365956 182112
rect 364352 5846 364380 180814
rect 364536 180798 364656 180826
rect 364628 176798 364656 180798
rect 364616 176792 364668 176798
rect 364616 176734 364668 176740
rect 364616 176656 364668 176662
rect 364616 176598 364668 176604
rect 364628 156754 364656 176598
rect 365732 172553 365760 182106
rect 365718 172544 365774 172553
rect 365718 172479 365774 172488
rect 365902 172544 365958 172553
rect 365902 172479 365958 172488
rect 365720 169992 365772 169998
rect 365718 169960 365720 169969
rect 365772 169960 365774 169969
rect 365718 169895 365774 169904
rect 365916 157298 365944 172479
rect 365824 157270 365944 157298
rect 365824 157026 365852 157270
rect 365824 156998 365944 157026
rect 364536 156726 364656 156754
rect 364536 147694 364564 156726
rect 364524 147688 364576 147694
rect 364524 147630 364576 147636
rect 364616 147620 364668 147626
rect 364616 147562 364668 147568
rect 364628 144906 364656 147562
rect 364524 144900 364576 144906
rect 364524 144842 364576 144848
rect 364616 144900 364668 144906
rect 364616 144842 364668 144848
rect 364536 125662 364564 144842
rect 365916 138666 365944 156998
rect 365916 138638 366036 138666
rect 366008 135318 366036 138638
rect 365996 135312 366048 135318
rect 365996 135254 366048 135260
rect 365904 135244 365956 135250
rect 365904 135186 365956 135192
rect 365916 133906 365944 135186
rect 365916 133878 366036 133906
rect 366008 125662 366036 133878
rect 364524 125656 364576 125662
rect 364524 125598 364576 125604
rect 365904 125656 365956 125662
rect 365904 125598 365956 125604
rect 365996 125656 366048 125662
rect 365996 125598 366048 125604
rect 364616 125520 364668 125526
rect 364616 125462 364668 125468
rect 364628 114458 364656 125462
rect 365916 124166 365944 125598
rect 365904 124160 365956 124166
rect 365904 124102 365956 124108
rect 365904 118652 365956 118658
rect 365904 118594 365956 118600
rect 364628 114430 364748 114458
rect 364720 109138 364748 114430
rect 364524 109132 364576 109138
rect 364524 109074 364576 109080
rect 364708 109132 364760 109138
rect 364708 109074 364760 109080
rect 364536 103766 364564 109074
rect 364524 103760 364576 103766
rect 364524 103702 364576 103708
rect 364708 103760 364760 103766
rect 364708 103702 364760 103708
rect 364720 93838 364748 103702
rect 364708 93832 364760 93838
rect 364708 93774 364760 93780
rect 365626 87272 365682 87281
rect 365626 87207 365628 87216
rect 365680 87207 365682 87216
rect 365628 87178 365680 87184
rect 364524 84244 364576 84250
rect 364524 84186 364576 84192
rect 364536 74526 364564 84186
rect 365916 80102 365944 118594
rect 365904 80096 365956 80102
rect 365904 80038 365956 80044
rect 365904 79960 365956 79966
rect 365904 79902 365956 79908
rect 364524 74520 364576 74526
rect 364524 74462 364576 74468
rect 364524 64932 364576 64938
rect 364524 64874 364576 64880
rect 364536 60874 364564 64874
rect 364536 60846 364656 60874
rect 364628 59786 364656 60846
rect 365916 60738 365944 79902
rect 365824 60710 365944 60738
rect 365824 60602 365852 60710
rect 365824 60574 365944 60602
rect 364536 59758 364656 59786
rect 364536 53122 364564 59758
rect 364536 53094 364656 53122
rect 364628 36038 364656 53094
rect 365916 47002 365944 60574
rect 365824 46974 365944 47002
rect 365824 40746 365852 46974
rect 365824 40718 365944 40746
rect 364616 36032 364668 36038
rect 364616 35974 364668 35980
rect 364524 35964 364576 35970
rect 364524 35906 364576 35912
rect 364536 31090 364564 35906
rect 364536 31062 364840 31090
rect 364812 26246 364840 31062
rect 365916 27554 365944 40718
rect 365916 27526 366036 27554
rect 364800 26240 364852 26246
rect 364800 26182 364852 26188
rect 366008 22778 366036 27526
rect 365720 22772 365772 22778
rect 365720 22714 365772 22720
rect 365996 22772 366048 22778
rect 365996 22714 366048 22720
rect 364800 17468 364852 17474
rect 364800 17410 364852 17416
rect 364812 8362 364840 17410
rect 365732 10538 365760 22714
rect 365720 10532 365772 10538
rect 365720 10474 365772 10480
rect 364432 8356 364484 8362
rect 364432 8298 364484 8304
rect 364800 8356 364852 8362
rect 364800 8298 364852 8304
rect 364444 8090 364472 8298
rect 364432 8084 364484 8090
rect 364432 8026 364484 8032
rect 364340 5840 364392 5846
rect 364340 5782 364392 5788
rect 365720 5024 365772 5030
rect 365720 4966 365772 4972
rect 363696 4004 363748 4010
rect 363696 3946 363748 3952
rect 364524 4004 364576 4010
rect 364524 3946 364576 3952
rect 363604 3256 363656 3262
rect 363604 3198 363656 3204
rect 363328 2984 363380 2990
rect 363328 2926 363380 2932
rect 363340 480 363368 2926
rect 364536 480 364564 3946
rect 365732 480 365760 4966
rect 366376 3126 366404 336874
rect 366468 4010 366496 336942
rect 366456 4004 366508 4010
rect 366456 3946 366508 3952
rect 366364 3120 366416 3126
rect 366364 3062 366416 3068
rect 366928 480 366956 337622
rect 367112 8158 367140 340068
rect 367204 340054 367770 340082
rect 367204 10674 367232 340054
rect 367848 328506 367876 340190
rect 368584 340054 368966 340082
rect 367284 328500 367336 328506
rect 367284 328442 367336 328448
rect 367836 328500 367888 328506
rect 367836 328442 367888 328448
rect 367296 328386 367324 328442
rect 367296 328358 367508 328386
rect 367480 309194 367508 328358
rect 367376 309188 367428 309194
rect 367376 309130 367428 309136
rect 367468 309188 367520 309194
rect 367468 309130 367520 309136
rect 367388 292670 367416 309130
rect 367376 292664 367428 292670
rect 367376 292606 367428 292612
rect 367376 292528 367428 292534
rect 367376 292470 367428 292476
rect 367388 273358 367416 292470
rect 367376 273352 367428 273358
rect 367376 273294 367428 273300
rect 367376 273216 367428 273222
rect 367376 273158 367428 273164
rect 367388 253994 367416 273158
rect 367296 253966 367416 253994
rect 367296 253858 367324 253966
rect 367296 253830 367416 253858
rect 367388 241482 367416 253830
rect 367388 241454 367508 241482
rect 367480 234666 367508 241454
rect 367468 234660 367520 234666
rect 367468 234602 367520 234608
rect 367376 234592 367428 234598
rect 367376 234534 367428 234540
rect 367388 222170 367416 234534
rect 367388 222142 367508 222170
rect 367480 215354 367508 222142
rect 367468 215348 367520 215354
rect 367468 215290 367520 215296
rect 367376 215280 367428 215286
rect 367376 215222 367428 215228
rect 367388 202858 367416 215222
rect 367388 202830 367508 202858
rect 367480 196042 367508 202830
rect 367468 196036 367520 196042
rect 367468 195978 367520 195984
rect 367376 195968 367428 195974
rect 367376 195910 367428 195916
rect 367388 135425 367416 195910
rect 368296 169992 368348 169998
rect 368294 169960 368296 169969
rect 368348 169960 368350 169969
rect 368294 169895 368350 169904
rect 367374 135416 367430 135425
rect 367374 135351 367430 135360
rect 367374 135280 367430 135289
rect 367374 135215 367376 135224
rect 367428 135215 367430 135224
rect 367560 135244 367612 135250
rect 367376 135186 367428 135192
rect 367560 135186 367612 135192
rect 367572 125633 367600 135186
rect 367374 125624 367430 125633
rect 367374 125559 367430 125568
rect 367558 125624 367614 125633
rect 367558 125559 367614 125568
rect 367388 99498 367416 125559
rect 367296 99470 367416 99498
rect 367296 99362 367324 99470
rect 367296 99334 367416 99362
rect 367388 80084 367416 99334
rect 367388 80056 367508 80084
rect 367480 79948 367508 80056
rect 367388 79920 367508 79948
rect 367388 55457 367416 79920
rect 367374 55448 367430 55457
rect 367374 55383 367430 55392
rect 367282 55312 367338 55321
rect 367282 55247 367338 55256
rect 367296 55214 367324 55247
rect 367284 55208 367336 55214
rect 367284 55150 367336 55156
rect 367376 55208 367428 55214
rect 367376 55150 367428 55156
rect 367388 45665 367416 55150
rect 367374 45656 367430 45665
rect 367374 45591 367430 45600
rect 367466 45520 367522 45529
rect 367466 45455 367522 45464
rect 367480 35970 367508 45455
rect 367376 35964 367428 35970
rect 367376 35906 367428 35912
rect 367468 35964 367520 35970
rect 367468 35906 367520 35912
rect 367388 31906 367416 35906
rect 367388 31878 367508 31906
rect 367480 31090 367508 31878
rect 367296 31062 367508 31090
rect 367296 26194 367324 31062
rect 367296 26166 367416 26194
rect 367192 10668 367244 10674
rect 367192 10610 367244 10616
rect 367388 10606 367416 26166
rect 367376 10600 367428 10606
rect 367376 10542 367428 10548
rect 368584 8226 368612 340054
rect 369596 337754 369624 340068
rect 369872 340054 370254 340082
rect 369584 337748 369636 337754
rect 369584 337690 369636 337696
rect 369768 280152 369820 280158
rect 369768 280094 369820 280100
rect 369780 274854 369808 280094
rect 369768 274848 369820 274854
rect 369768 274790 369820 274796
rect 369768 233912 369820 233918
rect 369768 233854 369820 233860
rect 369780 220862 369808 233854
rect 369768 220856 369820 220862
rect 369768 220798 369820 220804
rect 368572 8220 368624 8226
rect 368572 8162 368624 8168
rect 367100 8152 367152 8158
rect 367100 8094 367152 8100
rect 369872 5982 369900 340054
rect 370332 328506 370360 340190
rect 371436 337414 371464 340068
rect 371424 337408 371476 337414
rect 371424 337350 371476 337356
rect 371528 328574 371556 340190
rect 372646 340054 372752 340082
rect 372528 337408 372580 337414
rect 372528 337350 372580 337356
rect 371516 328568 371568 328574
rect 371516 328510 371568 328516
rect 370136 328500 370188 328506
rect 370136 328442 370188 328448
rect 370320 328500 370372 328506
rect 370320 328442 370372 328448
rect 371332 328500 371384 328506
rect 371332 328442 371384 328448
rect 370148 299470 370176 328442
rect 371344 323626 371372 328442
rect 371344 323598 371464 323626
rect 371436 318782 371464 323598
rect 371332 318776 371384 318782
rect 371332 318718 371384 318724
rect 371424 318776 371476 318782
rect 371424 318718 371476 318724
rect 371344 317422 371372 318718
rect 371332 317416 371384 317422
rect 371332 317358 371384 317364
rect 371332 309120 371384 309126
rect 371332 309062 371384 309068
rect 371344 304314 371372 309062
rect 371344 304286 371464 304314
rect 370044 299464 370096 299470
rect 370044 299406 370096 299412
rect 370136 299464 370188 299470
rect 370136 299406 370188 299412
rect 370056 298110 370084 299406
rect 370044 298104 370096 298110
rect 370044 298046 370096 298052
rect 371436 292482 371464 304286
rect 371344 292454 371464 292482
rect 371344 292210 371372 292454
rect 371344 292182 371464 292210
rect 370044 288448 370096 288454
rect 370044 288390 370096 288396
rect 370056 282946 370084 288390
rect 370044 282940 370096 282946
rect 370044 282882 370096 282888
rect 370136 282804 370188 282810
rect 370136 282746 370188 282752
rect 370148 280158 370176 282746
rect 371436 280158 371464 292182
rect 370136 280152 370188 280158
rect 370136 280094 370188 280100
rect 371424 280152 371476 280158
rect 371424 280094 371476 280100
rect 371516 280152 371568 280158
rect 371516 280094 371568 280100
rect 370136 274848 370188 274854
rect 370136 274790 370188 274796
rect 370148 267753 370176 274790
rect 371528 273170 371556 280094
rect 371436 273142 371556 273170
rect 369950 267744 370006 267753
rect 369950 267679 370006 267688
rect 370134 267744 370190 267753
rect 370134 267679 370190 267688
rect 369964 258097 369992 267679
rect 369950 258088 370006 258097
rect 369950 258023 370006 258032
rect 370134 258088 370190 258097
rect 370134 258023 370190 258032
rect 370148 254046 370176 258023
rect 370136 254040 370188 254046
rect 371436 253994 371464 273142
rect 370136 253982 370188 253988
rect 371344 253966 371464 253994
rect 371344 253858 371372 253966
rect 371344 253830 371464 253858
rect 370044 248532 370096 248538
rect 370044 248474 370096 248480
rect 370056 248402 370084 248474
rect 370044 248396 370096 248402
rect 370044 248338 370096 248344
rect 370320 248396 370372 248402
rect 370320 248338 370372 248344
rect 370332 233918 370360 248338
rect 370320 233912 370372 233918
rect 370320 233854 370372 233860
rect 369952 220856 370004 220862
rect 369952 220798 370004 220804
rect 369964 212498 369992 220798
rect 369952 212492 370004 212498
rect 369952 212434 370004 212440
rect 369952 202904 370004 202910
rect 369952 202846 370004 202852
rect 369964 201482 369992 202846
rect 369952 201476 370004 201482
rect 369952 201418 370004 201424
rect 369952 193180 370004 193186
rect 369952 193122 370004 193128
rect 369964 186266 369992 193122
rect 369964 186238 370176 186266
rect 370148 173942 370176 186238
rect 371146 180976 371202 180985
rect 371146 180911 371202 180920
rect 371160 180713 371188 180911
rect 371146 180704 371202 180713
rect 371146 180639 371202 180648
rect 371436 176610 371464 253830
rect 371344 176582 371464 176610
rect 371344 176338 371372 176582
rect 371344 176310 371464 176338
rect 370044 173936 370096 173942
rect 370044 173878 370096 173884
rect 370136 173936 370188 173942
rect 370136 173878 370188 173884
rect 370056 169402 370084 173878
rect 370056 169374 370176 169402
rect 370148 164218 370176 169374
rect 370136 164212 370188 164218
rect 370136 164154 370188 164160
rect 371436 157298 371464 176310
rect 371344 157270 371464 157298
rect 371344 157026 371372 157270
rect 371344 156998 371464 157026
rect 370044 154624 370096 154630
rect 370044 154566 370096 154572
rect 370056 147694 370084 154566
rect 370044 147688 370096 147694
rect 370044 147630 370096 147636
rect 370136 147620 370188 147626
rect 370136 147562 370188 147568
rect 370148 144906 370176 147562
rect 370136 144900 370188 144906
rect 370136 144842 370188 144848
rect 370228 144900 370280 144906
rect 370228 144842 370280 144848
rect 370240 135289 370268 144842
rect 371436 138122 371464 156998
rect 371344 138094 371464 138122
rect 371344 137714 371372 138094
rect 371344 137686 371464 137714
rect 370042 135280 370098 135289
rect 370042 135215 370098 135224
rect 370226 135280 370282 135289
rect 370226 135215 370282 135224
rect 370056 130370 370084 135215
rect 370056 130342 370268 130370
rect 370240 128194 370268 130342
rect 370148 128166 370268 128194
rect 370148 125594 370176 128166
rect 371436 125594 371464 137686
rect 369952 125588 370004 125594
rect 369952 125530 370004 125536
rect 370136 125588 370188 125594
rect 370136 125530 370188 125536
rect 371424 125588 371476 125594
rect 371424 125530 371476 125536
rect 371516 125588 371568 125594
rect 371516 125530 371568 125536
rect 369964 114646 369992 125530
rect 371528 118674 371556 125530
rect 371436 118646 371556 118674
rect 369952 114640 370004 114646
rect 369952 114582 370004 114588
rect 370044 114572 370096 114578
rect 370044 114514 370096 114520
rect 370056 106350 370084 114514
rect 370044 106344 370096 106350
rect 370044 106286 370096 106292
rect 370136 106208 370188 106214
rect 370136 106150 370188 106156
rect 370148 103494 370176 106150
rect 370136 103488 370188 103494
rect 370136 103430 370188 103436
rect 370320 103488 370372 103494
rect 370320 103430 370372 103436
rect 370332 76022 370360 103430
rect 371436 99498 371464 118646
rect 371344 99470 371464 99498
rect 371344 99362 371372 99470
rect 371344 99334 371464 99362
rect 370044 76016 370096 76022
rect 370044 75958 370096 75964
rect 370320 76016 370372 76022
rect 370320 75958 370372 75964
rect 370056 66434 370084 75958
rect 370044 66428 370096 66434
rect 370044 66370 370096 66376
rect 370044 66292 370096 66298
rect 370044 66234 370096 66240
rect 370056 60874 370084 66234
rect 370056 60846 370176 60874
rect 370148 59786 370176 60846
rect 371436 60738 371464 99334
rect 371344 60710 371464 60738
rect 371344 60602 371372 60710
rect 371344 60574 371464 60602
rect 370056 59758 370176 59786
rect 370056 46986 370084 59758
rect 371436 47002 371464 60574
rect 370044 46980 370096 46986
rect 370044 46922 370096 46928
rect 370136 46980 370188 46986
rect 370136 46922 370188 46928
rect 371344 46974 371464 47002
rect 370148 35970 370176 46922
rect 371344 40746 371372 46974
rect 371344 40718 371464 40746
rect 370044 35964 370096 35970
rect 370044 35906 370096 35912
rect 370136 35964 370188 35970
rect 370136 35906 370188 35912
rect 370056 12510 370084 35906
rect 371436 28966 371464 40718
rect 371240 28960 371292 28966
rect 371240 28902 371292 28908
rect 371424 28960 371476 28966
rect 371424 28902 371476 28908
rect 371252 19394 371280 28902
rect 371252 19366 371372 19394
rect 370044 12504 370096 12510
rect 370044 12446 370096 12452
rect 371344 12458 371372 19366
rect 369952 12436 370004 12442
rect 371344 12430 371464 12458
rect 369952 12378 370004 12384
rect 369964 9654 369992 12378
rect 371436 9738 371464 12430
rect 371252 9710 371464 9738
rect 371252 9654 371280 9710
rect 369952 9648 370004 9654
rect 369952 9590 370004 9596
rect 371240 9648 371292 9654
rect 371240 9590 371292 9596
rect 369860 5976 369912 5982
rect 369860 5918 369912 5924
rect 369216 5840 369268 5846
rect 369216 5782 369268 5788
rect 368020 3120 368072 3126
rect 368020 3062 368072 3068
rect 368032 480 368060 3062
rect 369228 480 369256 5782
rect 370412 3256 370464 3262
rect 370412 3198 370464 3204
rect 370424 480 370452 3198
rect 372540 2990 372568 337350
rect 372618 181248 372674 181257
rect 372618 181183 372620 181192
rect 372672 181183 372674 181192
rect 372620 181154 372672 181160
rect 372724 7546 372752 340054
rect 373276 337482 373304 340068
rect 373460 340054 373842 340082
rect 374104 340054 374486 340082
rect 373264 337476 373316 337482
rect 373264 337418 373316 337424
rect 373460 331242 373488 340054
rect 372816 331214 373488 331242
rect 372712 7540 372764 7546
rect 372712 7482 372764 7488
rect 372816 6186 372844 331214
rect 373908 87236 373960 87242
rect 373908 87178 373960 87184
rect 373920 87145 373948 87178
rect 373906 87136 373962 87145
rect 373906 87071 373962 87080
rect 373906 29336 373962 29345
rect 373906 29271 373962 29280
rect 373920 28937 373948 29271
rect 373906 28928 373962 28937
rect 373906 28863 373962 28872
rect 374104 7478 374132 340054
rect 375116 337822 375144 340068
rect 375392 340054 375682 340082
rect 375852 340054 376326 340082
rect 375104 337816 375156 337822
rect 375104 337758 375156 337764
rect 374644 337748 374696 337754
rect 374644 337690 374696 337696
rect 374092 7472 374144 7478
rect 374092 7414 374144 7420
rect 372804 6180 372856 6186
rect 372804 6122 372856 6128
rect 372896 6180 372948 6186
rect 372896 6122 372948 6128
rect 372908 4434 372936 6122
rect 372816 4406 372936 4434
rect 371608 2984 371660 2990
rect 371608 2926 371660 2932
rect 372528 2984 372580 2990
rect 372528 2926 372580 2932
rect 371620 480 371648 2926
rect 372816 480 372844 4406
rect 374656 3074 374684 337690
rect 375288 337476 375340 337482
rect 375288 337418 375340 337424
rect 375196 280152 375248 280158
rect 375196 280094 375248 280100
rect 375208 269074 375236 280094
rect 375196 269068 375248 269074
rect 375196 269010 375248 269016
rect 375194 204504 375250 204513
rect 375194 204439 375250 204448
rect 375208 204406 375236 204439
rect 375196 204400 375248 204406
rect 375196 204342 375248 204348
rect 374564 3058 374684 3074
rect 375196 3120 375248 3126
rect 375196 3062 375248 3068
rect 374552 3052 374684 3058
rect 374604 3046 374684 3052
rect 374552 2994 374604 3000
rect 374000 1964 374052 1970
rect 374000 1906 374052 1912
rect 374012 480 374040 1906
rect 375208 480 375236 3062
rect 375300 1970 375328 337418
rect 375392 6254 375420 340054
rect 375852 328386 375880 340054
rect 376024 337816 376076 337822
rect 376024 337758 376076 337764
rect 375760 328358 375880 328386
rect 375760 318850 375788 328358
rect 375564 318844 375616 318850
rect 375564 318786 375616 318792
rect 375748 318844 375800 318850
rect 375748 318786 375800 318792
rect 375576 318730 375604 318786
rect 375576 318702 375696 318730
rect 375668 299418 375696 318702
rect 375484 299390 375696 299418
rect 375484 298110 375512 299390
rect 375472 298104 375524 298110
rect 375472 298046 375524 298052
rect 375472 289808 375524 289814
rect 375472 289750 375524 289756
rect 375484 282878 375512 289750
rect 375472 282872 375524 282878
rect 375472 282814 375524 282820
rect 375656 282804 375708 282810
rect 375656 282746 375708 282752
rect 375668 280158 375696 282746
rect 375656 280152 375708 280158
rect 375656 280094 375708 280100
rect 375656 269068 375708 269074
rect 375656 269010 375708 269016
rect 375668 267753 375696 269010
rect 375470 267744 375526 267753
rect 375470 267679 375526 267688
rect 375654 267744 375710 267753
rect 375654 267679 375710 267688
rect 375484 258097 375512 267679
rect 375470 258088 375526 258097
rect 375470 258023 375526 258032
rect 375654 258088 375710 258097
rect 375654 258023 375710 258032
rect 375668 254046 375696 258023
rect 375656 254040 375708 254046
rect 375656 253982 375708 253988
rect 375564 248532 375616 248538
rect 375564 248474 375616 248480
rect 375576 248402 375604 248474
rect 375564 248396 375616 248402
rect 375564 248338 375616 248344
rect 375564 242820 375616 242826
rect 375564 242762 375616 242768
rect 375576 220862 375604 242762
rect 375472 220856 375524 220862
rect 375472 220798 375524 220804
rect 375564 220856 375616 220862
rect 375564 220798 375616 220804
rect 375484 220726 375512 220798
rect 375472 220720 375524 220726
rect 375472 220662 375524 220668
rect 375840 220720 375892 220726
rect 375840 220662 375892 220668
rect 375852 211177 375880 220662
rect 375654 211168 375710 211177
rect 375654 211103 375710 211112
rect 375838 211168 375894 211177
rect 375838 211103 375894 211112
rect 375668 196110 375696 211103
rect 375656 196104 375708 196110
rect 375656 196046 375708 196052
rect 375564 193248 375616 193254
rect 375564 193190 375616 193196
rect 375576 186266 375604 193190
rect 375576 186238 375696 186266
rect 375470 157584 375526 157593
rect 375470 157519 375526 157528
rect 375484 157321 375512 157519
rect 375470 157312 375526 157321
rect 375470 157247 375526 157256
rect 375668 154578 375696 186238
rect 375576 154562 375696 154578
rect 375564 154556 375696 154562
rect 375616 154550 375696 154556
rect 375564 154498 375616 154504
rect 375576 154467 375604 154498
rect 375564 147620 375616 147626
rect 375564 147562 375616 147568
rect 375576 144922 375604 147562
rect 375576 144906 375696 144922
rect 375564 144900 375708 144906
rect 375616 144894 375656 144900
rect 375564 144842 375616 144848
rect 375656 144842 375708 144848
rect 375576 128330 375604 144842
rect 375576 128302 375696 128330
rect 375668 99498 375696 128302
rect 375576 99470 375696 99498
rect 375576 93566 375604 99470
rect 375564 93560 375616 93566
rect 375564 93502 375616 93508
rect 375656 85604 375708 85610
rect 375656 85546 375708 85552
rect 375668 85490 375696 85546
rect 375576 85462 375696 85490
rect 375576 80084 375604 85462
rect 375576 80056 375788 80084
rect 375760 75970 375788 80056
rect 375576 75942 375788 75970
rect 375576 75886 375604 75942
rect 375564 75880 375616 75886
rect 375564 75822 375616 75828
rect 375564 56636 375616 56642
rect 375564 56578 375616 56584
rect 375576 56506 375604 56578
rect 375564 56500 375616 56506
rect 375564 56442 375616 56448
rect 375656 51740 375708 51746
rect 375656 51682 375708 51688
rect 375668 35986 375696 51682
rect 375576 35958 375696 35986
rect 375576 35902 375604 35958
rect 375564 35896 375616 35902
rect 375564 35838 375616 35844
rect 375748 35896 375800 35902
rect 375748 35838 375800 35844
rect 375760 9722 375788 35838
rect 375472 9716 375524 9722
rect 375472 9658 375524 9664
rect 375748 9716 375800 9722
rect 375748 9658 375800 9664
rect 375484 7410 375512 9658
rect 375472 7404 375524 7410
rect 375472 7346 375524 7352
rect 375380 6248 375432 6254
rect 375380 6190 375432 6196
rect 376036 3534 376064 337758
rect 376956 337550 376984 340068
rect 376944 337544 376996 337550
rect 376944 337486 376996 337492
rect 377048 335646 377076 340190
rect 378166 340054 378364 340082
rect 377036 335640 377088 335646
rect 377036 335582 377088 335588
rect 378232 335640 378284 335646
rect 378232 335582 378284 335588
rect 377036 327140 377088 327146
rect 377036 327082 377088 327088
rect 377048 318850 377076 327082
rect 376944 318844 376996 318850
rect 376944 318786 376996 318792
rect 377036 318844 377088 318850
rect 377036 318786 377088 318792
rect 376956 317422 376984 318786
rect 376944 317416 376996 317422
rect 376944 317358 376996 317364
rect 376944 307828 376996 307834
rect 376944 307770 376996 307776
rect 376956 299470 376984 307770
rect 376944 299464 376996 299470
rect 376944 299406 376996 299412
rect 376944 289876 376996 289882
rect 376944 289818 376996 289824
rect 376956 273222 376984 289818
rect 376944 273216 376996 273222
rect 376944 273158 376996 273164
rect 376944 273080 376996 273086
rect 376944 273022 376996 273028
rect 376956 253910 376984 273022
rect 376944 253904 376996 253910
rect 376944 253846 376996 253852
rect 376944 253768 376996 253774
rect 376944 253710 376996 253716
rect 376956 234598 376984 253710
rect 376944 234592 376996 234598
rect 376944 234534 376996 234540
rect 376944 234456 376996 234462
rect 376944 234398 376996 234404
rect 376956 215286 376984 234398
rect 376944 215280 376996 215286
rect 376944 215222 376996 215228
rect 376944 215144 376996 215150
rect 376944 215086 376996 215092
rect 376956 195974 376984 215086
rect 376944 195968 376996 195974
rect 376944 195910 376996 195916
rect 376944 195832 376996 195838
rect 376944 195774 376996 195780
rect 376956 169114 376984 195774
rect 376944 169108 376996 169114
rect 376944 169050 376996 169056
rect 377128 169108 377180 169114
rect 377128 169050 377180 169056
rect 377140 164257 377168 169050
rect 376942 164248 376998 164257
rect 376942 164183 376944 164192
rect 376996 164183 376998 164192
rect 377126 164248 377182 164257
rect 377126 164183 377182 164192
rect 376944 164154 376996 164160
rect 376944 154624 376996 154630
rect 376944 154566 376996 154572
rect 376956 138038 376984 154566
rect 376944 138032 376996 138038
rect 376944 137974 376996 137980
rect 376944 137896 376996 137902
rect 376944 137838 376996 137844
rect 376956 99498 376984 137838
rect 376864 99470 376984 99498
rect 376864 99362 376892 99470
rect 376864 99334 376984 99362
rect 376956 80102 376984 99334
rect 376944 80096 376996 80102
rect 376944 80038 376996 80044
rect 376944 79960 376996 79966
rect 376944 79902 376996 79908
rect 376956 67726 376984 79902
rect 376944 67720 376996 67726
rect 376944 67662 376996 67668
rect 376852 67652 376904 67658
rect 376852 67594 376904 67600
rect 376864 38690 376892 67594
rect 376852 38684 376904 38690
rect 376852 38626 376904 38632
rect 376944 38684 376996 38690
rect 376944 38626 376996 38632
rect 376956 29050 376984 38626
rect 376864 29022 376984 29050
rect 376864 27606 376892 29022
rect 376852 27600 376904 27606
rect 376852 27542 376904 27548
rect 377036 27600 377088 27606
rect 377036 27542 377088 27548
rect 377048 9994 377076 27542
rect 377036 9988 377088 9994
rect 377036 9930 377088 9936
rect 378244 6390 378272 335582
rect 378336 10334 378364 340054
rect 378428 340054 378810 340082
rect 379072 340054 379362 340082
rect 379624 340054 380006 340082
rect 378324 10328 378376 10334
rect 378324 10270 378376 10276
rect 378232 6384 378284 6390
rect 378232 6326 378284 6332
rect 376392 5092 376444 5098
rect 376392 5034 376444 5040
rect 376024 3528 376076 3534
rect 376024 3470 376076 3476
rect 375288 1964 375340 1970
rect 375288 1906 375340 1912
rect 376404 480 376432 5034
rect 378428 3738 378456 340054
rect 379072 335646 379100 340054
rect 379060 335640 379112 335646
rect 379060 335582 379112 335588
rect 379334 170096 379390 170105
rect 379518 170096 379574 170105
rect 379390 170054 379518 170082
rect 379334 170031 379390 170040
rect 379518 170031 379574 170040
rect 379624 10470 379652 340054
rect 380636 337618 380664 340068
rect 380912 340054 381202 340082
rect 380624 337612 380676 337618
rect 380624 337554 380676 337560
rect 380806 220824 380862 220833
rect 380806 220759 380862 220768
rect 380820 211177 380848 220759
rect 380806 211168 380862 211177
rect 380806 211103 380862 211112
rect 380808 22228 380860 22234
rect 380808 22170 380860 22176
rect 379612 10464 379664 10470
rect 379612 10406 379664 10412
rect 380820 6730 380848 22170
rect 380808 6724 380860 6730
rect 380808 6666 380860 6672
rect 379980 6248 380032 6254
rect 379980 6190 380032 6196
rect 378416 3732 378468 3738
rect 378416 3674 378468 3680
rect 378784 3052 378836 3058
rect 378784 2994 378836 3000
rect 377588 2984 377640 2990
rect 377588 2926 377640 2932
rect 377600 480 377628 2926
rect 378796 480 378824 2994
rect 379992 480 380020 6190
rect 380912 5302 380940 340054
rect 381280 338042 381308 340190
rect 381188 338014 381308 338042
rect 381188 331158 381216 338014
rect 382476 336802 382504 340068
rect 382660 340054 383042 340082
rect 383686 340054 383792 340082
rect 381544 336796 381596 336802
rect 381544 336738 381596 336744
rect 382464 336796 382516 336802
rect 382464 336738 382516 336744
rect 381176 331152 381228 331158
rect 381176 331094 381228 331100
rect 381084 328500 381136 328506
rect 381136 328460 381216 328488
rect 381084 328442 381136 328448
rect 381188 319025 381216 328460
rect 381174 319016 381230 319025
rect 381174 318951 381230 318960
rect 381082 318880 381138 318889
rect 381082 318815 381138 318824
rect 381096 317422 381124 318815
rect 381084 317416 381136 317422
rect 381084 317358 381136 317364
rect 381360 317416 381412 317422
rect 381360 317358 381412 317364
rect 381372 289882 381400 317358
rect 381084 289876 381136 289882
rect 381084 289818 381136 289824
rect 381360 289876 381412 289882
rect 381360 289818 381412 289824
rect 381096 282946 381124 289818
rect 381084 282940 381136 282946
rect 381084 282882 381136 282888
rect 381176 282804 381228 282810
rect 381176 282746 381228 282752
rect 381188 280090 381216 282746
rect 381176 280084 381228 280090
rect 381176 280026 381228 280032
rect 381084 270564 381136 270570
rect 381084 270506 381136 270512
rect 381096 270434 381124 270506
rect 381084 270428 381136 270434
rect 381084 270370 381136 270376
rect 381176 260908 381228 260914
rect 381176 260850 381228 260856
rect 381188 260794 381216 260850
rect 381188 260766 381308 260794
rect 381280 251326 381308 260766
rect 381268 251320 381320 251326
rect 381268 251262 381320 251268
rect 381084 251252 381136 251258
rect 381084 251194 381136 251200
rect 381096 244322 381124 251194
rect 381084 244316 381136 244322
rect 381084 244258 381136 244264
rect 381176 244180 381228 244186
rect 381176 244122 381228 244128
rect 381188 241482 381216 244122
rect 381096 241454 381216 241482
rect 381096 240122 381124 241454
rect 381096 240094 381216 240122
rect 381188 234666 381216 240094
rect 381176 234660 381228 234666
rect 381176 234602 381228 234608
rect 381084 234592 381136 234598
rect 381084 234534 381136 234540
rect 381096 225010 381124 234534
rect 381084 225004 381136 225010
rect 381084 224946 381136 224952
rect 381176 224868 381228 224874
rect 381176 224810 381228 224816
rect 381188 222170 381216 224810
rect 381096 222142 381216 222170
rect 381096 220833 381124 222142
rect 381082 220824 381138 220833
rect 381082 220759 381138 220768
rect 380990 211168 381046 211177
rect 380990 211103 381046 211112
rect 381004 205578 381032 211103
rect 381004 205550 381216 205578
rect 381188 202858 381216 205550
rect 381096 202830 381216 202858
rect 381096 186266 381124 202830
rect 381096 186238 381216 186266
rect 381188 154578 381216 186238
rect 381096 154562 381216 154578
rect 381084 154556 381216 154562
rect 381136 154550 381216 154556
rect 381084 154498 381136 154504
rect 381096 154467 381124 154498
rect 381084 147620 381136 147626
rect 381084 147562 381136 147568
rect 381096 144922 381124 147562
rect 381096 144894 381216 144922
rect 381188 144838 381216 144894
rect 381176 144832 381228 144838
rect 381176 144774 381228 144780
rect 381084 135312 381136 135318
rect 381084 135254 381136 135260
rect 381096 128330 381124 135254
rect 381096 128302 381216 128330
rect 381188 125594 381216 128302
rect 381176 125588 381228 125594
rect 381176 125530 381228 125536
rect 381176 116000 381228 116006
rect 381176 115942 381228 115948
rect 381188 99498 381216 115942
rect 381096 99470 381216 99498
rect 381096 89826 381124 99470
rect 381084 89820 381136 89826
rect 381084 89762 381136 89768
rect 380992 87032 381044 87038
rect 380992 86974 381044 86980
rect 381004 85542 381032 86974
rect 380992 85536 381044 85542
rect 380992 85478 381044 85484
rect 381084 75948 381136 75954
rect 381084 75890 381136 75896
rect 381096 67590 381124 75890
rect 381084 67584 381136 67590
rect 381084 67526 381136 67532
rect 381084 57996 381136 58002
rect 381084 57938 381136 57944
rect 381096 53122 381124 57938
rect 381096 53094 381308 53122
rect 381280 50946 381308 53094
rect 381188 50918 381308 50946
rect 381188 48278 381216 50918
rect 380992 48272 381044 48278
rect 380992 48214 381044 48220
rect 381176 48272 381228 48278
rect 381176 48214 381228 48220
rect 381004 41290 381032 48214
rect 381004 41262 381124 41290
rect 381096 29034 381124 41262
rect 381084 29028 381136 29034
rect 381084 28970 381136 28976
rect 381176 29028 381228 29034
rect 381176 28970 381228 28976
rect 381188 22234 381216 28970
rect 381176 22228 381228 22234
rect 381176 22170 381228 22176
rect 380900 5296 380952 5302
rect 380900 5238 380952 5244
rect 381556 3602 381584 336738
rect 382660 336734 382688 340054
rect 382924 336796 382976 336802
rect 382924 336738 382976 336744
rect 382648 336728 382700 336734
rect 382648 336670 382700 336676
rect 382464 336660 382516 336666
rect 382464 336602 382516 336608
rect 382476 327078 382504 336602
rect 382464 327072 382516 327078
rect 382464 327014 382516 327020
rect 382464 317552 382516 317558
rect 382464 317494 382516 317500
rect 382476 317422 382504 317494
rect 382464 317416 382516 317422
rect 382464 317358 382516 317364
rect 382464 307828 382516 307834
rect 382464 307770 382516 307776
rect 382476 298042 382504 307770
rect 382464 298036 382516 298042
rect 382464 297978 382516 297984
rect 382556 298036 382608 298042
rect 382556 297978 382608 297984
rect 382568 292482 382596 297978
rect 382476 292454 382596 292482
rect 382476 280158 382504 292454
rect 382464 280152 382516 280158
rect 382464 280094 382516 280100
rect 382464 270564 382516 270570
rect 382464 270506 382516 270512
rect 382476 260846 382504 270506
rect 382464 260840 382516 260846
rect 382464 260782 382516 260788
rect 382464 251252 382516 251258
rect 382464 251194 382516 251200
rect 382476 241505 382504 251194
rect 382278 241496 382334 241505
rect 382278 241431 382334 241440
rect 382462 241496 382518 241505
rect 382462 241431 382518 241440
rect 382292 231878 382320 241431
rect 382280 231872 382332 231878
rect 382280 231814 382332 231820
rect 382464 231872 382516 231878
rect 382464 231814 382516 231820
rect 382476 222193 382504 231814
rect 382278 222184 382334 222193
rect 382278 222119 382334 222128
rect 382462 222184 382518 222193
rect 382462 222119 382518 222128
rect 382292 212566 382320 222119
rect 382280 212560 382332 212566
rect 382280 212502 382332 212508
rect 382464 212560 382516 212566
rect 382464 212502 382516 212508
rect 382476 202881 382504 212502
rect 382278 202872 382334 202881
rect 382278 202807 382334 202816
rect 382462 202872 382518 202881
rect 382462 202807 382518 202816
rect 382292 193254 382320 202807
rect 382280 193248 382332 193254
rect 382280 193190 382332 193196
rect 382464 193248 382516 193254
rect 382464 193190 382516 193196
rect 382476 183666 382504 193190
rect 382464 183660 382516 183666
rect 382464 183602 382516 183608
rect 382464 183524 382516 183530
rect 382464 183466 382516 183472
rect 382476 182209 382504 183466
rect 382278 182200 382334 182209
rect 382278 182135 382334 182144
rect 382462 182200 382518 182209
rect 382462 182135 382518 182144
rect 382188 181212 382240 181218
rect 382188 181154 382240 181160
rect 382200 180985 382228 181154
rect 382186 180976 382242 180985
rect 382186 180911 382242 180920
rect 382292 167686 382320 182135
rect 382280 167680 382332 167686
rect 382280 167622 382332 167628
rect 382464 154624 382516 154630
rect 382464 154566 382516 154572
rect 382476 138038 382504 154566
rect 382464 138032 382516 138038
rect 382464 137974 382516 137980
rect 382464 137896 382516 137902
rect 382464 137838 382516 137844
rect 382476 99498 382504 137838
rect 382384 99470 382504 99498
rect 382384 99362 382412 99470
rect 382384 99334 382504 99362
rect 382476 86970 382504 99334
rect 382464 86964 382516 86970
rect 382464 86906 382516 86912
rect 382464 75948 382516 75954
rect 382464 75890 382516 75896
rect 382476 51134 382504 75890
rect 382464 51128 382516 51134
rect 382464 51070 382516 51076
rect 382372 48340 382424 48346
rect 382372 48282 382424 48288
rect 382384 38690 382412 48282
rect 382372 38684 382424 38690
rect 382372 38626 382424 38632
rect 382464 38684 382516 38690
rect 382464 38626 382516 38632
rect 382476 29050 382504 38626
rect 382384 29022 382504 29050
rect 382384 27606 382412 29022
rect 382372 27600 382424 27606
rect 382372 27542 382424 27548
rect 382648 27600 382700 27606
rect 382648 27542 382700 27548
rect 382660 13122 382688 27542
rect 382648 13116 382700 13122
rect 382648 13058 382700 13064
rect 382936 3670 382964 336738
rect 383660 134088 383712 134094
rect 383658 134056 383660 134065
rect 383712 134056 383714 134065
rect 383658 133991 383714 134000
rect 383566 63744 383622 63753
rect 383566 63679 383622 63688
rect 383580 63481 383608 63679
rect 383566 63472 383622 63481
rect 383566 63407 383622 63416
rect 383566 40216 383622 40225
rect 383566 40151 383622 40160
rect 383580 40089 383608 40151
rect 383566 40080 383622 40089
rect 383566 40015 383622 40024
rect 383566 29608 383622 29617
rect 383566 29543 383622 29552
rect 383580 29209 383608 29543
rect 383566 29200 383622 29209
rect 383566 29135 383622 29144
rect 383764 10402 383792 340054
rect 384040 340054 384330 340082
rect 384500 340054 384882 340082
rect 385144 340054 385526 340082
rect 384040 337550 384068 340054
rect 384028 337544 384080 337550
rect 384028 337486 384080 337492
rect 384500 331242 384528 340054
rect 383856 331214 384528 331242
rect 383752 10396 383804 10402
rect 383752 10338 383804 10344
rect 383856 5438 383884 331214
rect 384946 204504 385002 204513
rect 384946 204439 385002 204448
rect 384960 204406 384988 204439
rect 384948 204400 385000 204406
rect 384948 204342 385000 204348
rect 384946 87272 385002 87281
rect 384946 87207 385002 87216
rect 384960 86873 384988 87207
rect 384946 86864 385002 86873
rect 384946 86799 385002 86808
rect 385144 6662 385172 340054
rect 385684 337952 385736 337958
rect 385684 337894 385736 337900
rect 385222 134192 385278 134201
rect 385222 134127 385278 134136
rect 385236 134094 385264 134127
rect 385224 134088 385276 134094
rect 385224 134030 385276 134036
rect 385132 6656 385184 6662
rect 385132 6598 385184 6604
rect 383844 5432 383896 5438
rect 383844 5374 383896 5380
rect 383568 5160 383620 5166
rect 383568 5102 383620 5108
rect 382924 3664 382976 3670
rect 382924 3606 382976 3612
rect 381544 3596 381596 3602
rect 381544 3538 381596 3544
rect 382372 3528 382424 3534
rect 382372 3470 382424 3476
rect 381176 3188 381228 3194
rect 381176 3130 381228 3136
rect 381188 480 381216 3130
rect 382384 480 382412 3470
rect 383580 480 383608 5102
rect 384672 2916 384724 2922
rect 384672 2858 384724 2864
rect 384684 480 384712 2858
rect 385696 2854 385724 337894
rect 386156 336802 386184 340068
rect 386432 340054 386722 340082
rect 386892 340054 387366 340082
rect 386144 336796 386196 336802
rect 386144 336738 386196 336744
rect 386432 6458 386460 340054
rect 386892 328506 386920 340054
rect 387996 337890 388024 340068
rect 387984 337884 388036 337890
rect 387984 337826 388036 337832
rect 388088 331242 388116 340190
rect 389206 340054 389312 340082
rect 389088 337544 389140 337550
rect 389088 337486 389140 337492
rect 387996 331214 388116 331242
rect 386696 328500 386748 328506
rect 386696 328442 386748 328448
rect 386880 328500 386932 328506
rect 386880 328442 386932 328448
rect 386708 318782 386736 328442
rect 387996 321638 388024 331214
rect 387984 321632 388036 321638
rect 387984 321574 388036 321580
rect 388076 321428 388128 321434
rect 388076 321370 388128 321376
rect 386696 318776 386748 318782
rect 386696 318718 386748 318724
rect 386696 309188 386748 309194
rect 386696 309130 386748 309136
rect 386708 292618 386736 309130
rect 388088 292618 388116 321370
rect 386616 292590 386736 292618
rect 387904 292590 388116 292618
rect 386616 287094 386644 292590
rect 387904 292482 387932 292590
rect 387904 292454 388024 292482
rect 386604 287088 386656 287094
rect 386604 287030 386656 287036
rect 386708 278798 386736 278829
rect 386696 278792 386748 278798
rect 386616 278740 386696 278746
rect 386616 278734 386748 278740
rect 386616 278718 386736 278734
rect 386616 273290 386644 278718
rect 386604 273284 386656 273290
rect 386604 273226 386656 273232
rect 386604 269204 386656 269210
rect 386604 269146 386656 269152
rect 386616 264314 386644 269146
rect 386604 264308 386656 264314
rect 386604 264250 386656 264256
rect 386512 259480 386564 259486
rect 386512 259422 386564 259428
rect 386524 251190 386552 259422
rect 387996 253910 388024 292454
rect 387984 253904 388036 253910
rect 387984 253846 388036 253852
rect 387984 253768 388036 253774
rect 387984 253710 388036 253716
rect 386512 251184 386564 251190
rect 386512 251126 386564 251132
rect 386880 251184 386932 251190
rect 386880 251126 386932 251132
rect 386892 231878 386920 251126
rect 387996 234598 388024 253710
rect 387984 234592 388036 234598
rect 387984 234534 388036 234540
rect 387984 234456 388036 234462
rect 387984 234398 388036 234404
rect 386604 231872 386656 231878
rect 386602 231840 386604 231849
rect 386880 231872 386932 231878
rect 386656 231840 386658 231849
rect 386602 231775 386658 231784
rect 386878 231840 386880 231849
rect 386932 231840 386934 231849
rect 386878 231775 386934 231784
rect 386892 212566 386920 231775
rect 387996 215286 388024 234398
rect 387984 215280 388036 215286
rect 387984 215222 388036 215228
rect 387984 215144 388036 215150
rect 387984 215086 388036 215092
rect 386604 212560 386656 212566
rect 386604 212502 386656 212508
rect 386880 212560 386932 212566
rect 386880 212502 386932 212508
rect 386616 209778 386644 212502
rect 386604 209772 386656 209778
rect 386604 209714 386656 209720
rect 386788 209772 386840 209778
rect 386788 209714 386840 209720
rect 386800 200138 386828 209714
rect 386800 200122 386920 200138
rect 386604 200116 386656 200122
rect 386800 200116 386932 200122
rect 386800 200110 386880 200116
rect 386604 200058 386656 200064
rect 386880 200058 386932 200064
rect 386616 198694 386644 200058
rect 386604 198688 386656 198694
rect 386604 198630 386656 198636
rect 387996 195974 388024 215086
rect 387984 195968 388036 195974
rect 387984 195910 388036 195916
rect 387984 195832 388036 195838
rect 387984 195774 388036 195780
rect 386604 186312 386656 186318
rect 386604 186254 386656 186260
rect 386616 180826 386644 186254
rect 386616 180798 386736 180826
rect 386708 176798 386736 180798
rect 386696 176792 386748 176798
rect 387996 176746 388024 195774
rect 386696 176734 386748 176740
rect 387904 176718 388024 176746
rect 386696 176656 386748 176662
rect 386696 176598 386748 176604
rect 387904 176610 387932 176718
rect 386708 164218 386736 176598
rect 387904 176582 388024 176610
rect 386696 164212 386748 164218
rect 386696 164154 386748 164160
rect 386788 164212 386840 164218
rect 386788 164154 386840 164160
rect 386800 154601 386828 164154
rect 387996 157486 388024 176582
rect 387984 157480 388036 157486
rect 387984 157422 388036 157428
rect 387984 157344 388036 157350
rect 387984 157286 388036 157292
rect 386602 154592 386658 154601
rect 386602 154527 386604 154536
rect 386656 154527 386658 154536
rect 386786 154592 386842 154601
rect 386786 154527 386788 154536
rect 386604 154498 386656 154504
rect 386840 154527 386842 154536
rect 386788 154498 386840 154504
rect 386800 135425 386828 154498
rect 386786 135416 386842 135425
rect 386786 135351 386842 135360
rect 386602 135280 386658 135289
rect 386602 135215 386658 135224
rect 386616 133890 386644 135215
rect 386604 133884 386656 133890
rect 386604 133826 386656 133832
rect 386696 122936 386748 122942
rect 386616 122884 386696 122890
rect 386616 122878 386748 122884
rect 386616 122862 386736 122878
rect 386616 121446 386644 122862
rect 386604 121440 386656 121446
rect 386604 121382 386656 121388
rect 387996 118810 388024 157286
rect 387904 118782 388024 118810
rect 387904 118674 387932 118782
rect 387904 118646 388024 118674
rect 386880 103556 386932 103562
rect 386880 103498 386932 103504
rect 386892 103442 386920 103498
rect 386800 103414 386920 103442
rect 386800 93974 386828 103414
rect 387996 96778 388024 118646
rect 387996 96750 388116 96778
rect 388088 96665 388116 96750
rect 388074 96656 388130 96665
rect 388074 96591 388130 96600
rect 387982 96520 388038 96529
rect 387982 96455 388038 96464
rect 386788 93968 386840 93974
rect 386788 93910 386840 93916
rect 386880 93900 386932 93906
rect 386880 93842 386932 93848
rect 386892 86850 386920 93842
rect 386616 86822 386920 86850
rect 386616 77450 386644 86822
rect 387996 80102 388024 96455
rect 387984 80096 388036 80102
rect 387984 80038 388036 80044
rect 387984 79960 388036 79966
rect 387984 79902 388036 79908
rect 386604 77444 386656 77450
rect 386604 77386 386656 77392
rect 386604 77308 386656 77314
rect 386604 77250 386656 77256
rect 386616 61470 386644 77250
rect 386604 61464 386656 61470
rect 386604 61406 386656 61412
rect 386788 61464 386840 61470
rect 386788 61406 386840 61412
rect 386800 48362 386828 61406
rect 387996 60738 388024 79902
rect 387904 60710 388024 60738
rect 387904 60602 387932 60710
rect 387904 60574 388024 60602
rect 387996 57934 388024 60574
rect 387892 57928 387944 57934
rect 387892 57870 387944 57876
rect 387984 57928 388036 57934
rect 387984 57870 388036 57876
rect 386708 48334 386828 48362
rect 386708 48278 386736 48334
rect 386696 48272 386748 48278
rect 386696 48214 386748 48220
rect 386788 48272 386840 48278
rect 386788 48214 386840 48220
rect 386800 29102 386828 48214
rect 387904 38570 387932 57870
rect 387904 38542 388116 38570
rect 386788 29096 386840 29102
rect 386788 29038 386840 29044
rect 388088 29034 388116 38542
rect 386696 29028 386748 29034
rect 386696 28970 386748 28976
rect 387892 29028 387944 29034
rect 387892 28970 387944 28976
rect 388076 29028 388128 29034
rect 388076 28970 388128 28976
rect 386708 22114 386736 28970
rect 387904 22250 387932 28970
rect 387812 22222 387932 22250
rect 386708 22086 386828 22114
rect 386800 21978 386828 22086
rect 386616 21950 386828 21978
rect 387812 21978 387840 22222
rect 387812 21950 387932 21978
rect 386616 14634 386644 21950
rect 386616 14606 386736 14634
rect 386708 14362 386736 14606
rect 386524 14334 386736 14362
rect 386524 6798 386552 14334
rect 386512 6792 386564 6798
rect 386512 6734 386564 6740
rect 387904 6526 387932 21950
rect 387892 6520 387944 6526
rect 387892 6462 387944 6468
rect 386420 6452 386472 6458
rect 386420 6394 386472 6400
rect 387064 5228 387116 5234
rect 387064 5170 387116 5176
rect 385868 3732 385920 3738
rect 385868 3674 385920 3680
rect 385684 2848 385736 2854
rect 385684 2790 385736 2796
rect 385880 480 385908 3674
rect 387076 480 387104 5170
rect 389100 3670 389128 337486
rect 389284 9042 389312 340054
rect 389744 337958 389772 340068
rect 389836 340054 390402 340082
rect 390664 340054 391046 340082
rect 389732 337952 389784 337958
rect 389732 337894 389784 337900
rect 389836 335730 389864 340054
rect 389916 336796 389968 336802
rect 389916 336738 389968 336744
rect 389376 335702 389864 335730
rect 389272 9036 389324 9042
rect 389272 8978 389324 8984
rect 389376 6594 389404 335702
rect 389928 335594 389956 336738
rect 389836 335566 389956 335594
rect 389364 6588 389416 6594
rect 389364 6530 389416 6536
rect 389836 3806 389864 335566
rect 390664 9178 390692 340054
rect 391204 337884 391256 337890
rect 391204 337826 391256 337832
rect 390652 9172 390704 9178
rect 390652 9114 390704 9120
rect 390652 5296 390704 5302
rect 390652 5238 390704 5244
rect 389824 3800 389876 3806
rect 389824 3742 389876 3748
rect 388260 3664 388312 3670
rect 388260 3606 388312 3612
rect 389088 3664 389140 3670
rect 389088 3606 389140 3612
rect 388272 480 388300 3606
rect 389456 3596 389508 3602
rect 389456 3538 389508 3544
rect 389468 480 389496 3538
rect 390664 480 390692 5238
rect 391216 3942 391244 337826
rect 391584 337618 391612 340068
rect 391952 340054 392242 340082
rect 391572 337612 391624 337618
rect 391572 337554 391624 337560
rect 391952 5506 391980 340054
rect 392320 338042 392348 340190
rect 392320 338014 392440 338042
rect 392412 328522 392440 338014
rect 393228 337612 393280 337618
rect 393228 337554 393280 337560
rect 392320 328494 392440 328522
rect 392320 328438 392348 328494
rect 393240 328438 393268 337554
rect 393424 336802 393452 340068
rect 393516 340054 394082 340082
rect 394726 340054 394832 340082
rect 393412 336796 393464 336802
rect 393412 336738 393464 336744
rect 392308 328432 392360 328438
rect 392308 328374 392360 328380
rect 393228 328432 393280 328438
rect 393228 328374 393280 328380
rect 392400 318844 392452 318850
rect 392400 318786 392452 318792
rect 393228 318844 393280 318850
rect 393228 318786 393280 318792
rect 392412 318730 392440 318786
rect 392412 318702 392532 318730
rect 392504 310962 392532 318702
rect 392032 310956 392084 310962
rect 392032 310898 392084 310904
rect 392492 310956 392544 310962
rect 392492 310898 392544 310904
rect 392044 298194 392072 310898
rect 392044 298166 392164 298194
rect 392136 296698 392164 298166
rect 392136 296670 392256 296698
rect 392228 292602 392256 296670
rect 392216 292596 392268 292602
rect 392216 292538 392268 292544
rect 392124 292528 392176 292534
rect 392124 292470 392176 292476
rect 392136 278769 392164 292470
rect 393240 278769 393268 318786
rect 392122 278760 392178 278769
rect 392122 278695 392178 278704
rect 393226 278760 393282 278769
rect 393226 278695 393282 278704
rect 393410 278760 393466 278769
rect 393410 278695 393466 278704
rect 392214 278624 392270 278633
rect 392214 278559 392270 278568
rect 392228 264314 392256 278559
rect 393424 269142 393452 278695
rect 393228 269136 393280 269142
rect 393226 269104 393228 269113
rect 393412 269136 393464 269142
rect 393280 269104 393282 269113
rect 393226 269039 393282 269048
rect 393410 269104 393412 269113
rect 393464 269104 393466 269113
rect 393410 269039 393466 269048
rect 392216 264308 392268 264314
rect 392216 264250 392268 264256
rect 393424 259486 393452 269039
rect 392032 259480 392084 259486
rect 392032 259422 392084 259428
rect 393228 259480 393280 259486
rect 393228 259422 393280 259428
rect 393412 259480 393464 259486
rect 393412 259422 393464 259428
rect 392044 241534 392072 259422
rect 393240 251326 393268 259422
rect 393228 251320 393280 251326
rect 393228 251262 393280 251268
rect 393136 251116 393188 251122
rect 393136 251058 393188 251064
rect 393148 249801 393176 251058
rect 392950 249792 393006 249801
rect 392950 249727 393006 249736
rect 393134 249792 393190 249801
rect 393134 249727 393190 249736
rect 392032 241528 392084 241534
rect 392124 241528 392176 241534
rect 392032 241470 392084 241476
rect 392122 241496 392124 241505
rect 392176 241496 392178 241505
rect 392122 241431 392178 241440
rect 392306 241496 392362 241505
rect 392306 241431 392362 241440
rect 392320 240145 392348 241431
rect 392964 240174 392992 249727
rect 392952 240168 393004 240174
rect 392306 240136 392362 240145
rect 392306 240071 392362 240080
rect 392490 240136 392546 240145
rect 392952 240110 393004 240116
rect 393228 240168 393280 240174
rect 393228 240110 393280 240116
rect 392490 240071 392546 240080
rect 392504 231554 392532 240071
rect 392320 231526 392532 231554
rect 392320 222222 392348 231526
rect 392124 222216 392176 222222
rect 392122 222184 392124 222193
rect 392308 222216 392360 222222
rect 392176 222184 392178 222193
rect 392308 222158 392360 222164
rect 392122 222119 392178 222128
rect 392214 222048 392270 222057
rect 392214 221983 392270 221992
rect 392228 202858 392256 221983
rect 392136 202830 392256 202858
rect 392136 193254 392164 202830
rect 392124 193248 392176 193254
rect 392124 193190 392176 193196
rect 392216 193248 392268 193254
rect 392216 193190 392268 193196
rect 392228 176746 392256 193190
rect 392136 176718 392256 176746
rect 392136 154737 392164 176718
rect 393240 164286 393268 240110
rect 393228 164280 393280 164286
rect 393228 164222 393280 164228
rect 393228 164144 393280 164150
rect 393228 164086 393280 164092
rect 393240 162858 393268 164086
rect 393228 162852 393280 162858
rect 393228 162794 393280 162800
rect 392122 154728 392178 154737
rect 392122 154663 392178 154672
rect 392122 154592 392178 154601
rect 392122 154527 392124 154536
rect 392176 154527 392178 154536
rect 392124 154498 392176 154504
rect 392124 147620 392176 147626
rect 392124 147562 392176 147568
rect 392136 144922 392164 147562
rect 393228 145036 393280 145042
rect 393228 144978 393280 144984
rect 392136 144894 392256 144922
rect 392228 138281 392256 144894
rect 393240 143546 393268 144978
rect 393228 143540 393280 143546
rect 393228 143482 393280 143488
rect 392214 138272 392270 138281
rect 392214 138207 392270 138216
rect 392122 135280 392178 135289
rect 392122 135215 392178 135224
rect 392136 125610 392164 135215
rect 393228 133952 393280 133958
rect 393228 133894 393280 133900
rect 393240 125769 393268 133894
rect 393226 125760 393282 125769
rect 393226 125695 393282 125704
rect 393226 125624 393282 125633
rect 392136 125582 392256 125610
rect 392228 119354 392256 125582
rect 393226 125559 393282 125568
rect 392136 119326 392256 119354
rect 392136 118674 392164 119326
rect 392136 118646 392256 118674
rect 392228 118402 392256 118646
rect 392136 118374 392256 118402
rect 392136 109018 392164 118374
rect 393240 114714 393268 125559
rect 393228 114708 393280 114714
rect 393228 114650 393280 114656
rect 393228 114572 393280 114578
rect 393228 114514 393280 114520
rect 392136 108990 392348 109018
rect 392320 106282 392348 108990
rect 392032 106276 392084 106282
rect 392032 106218 392084 106224
rect 392308 106276 392360 106282
rect 392308 106218 392360 106224
rect 392044 96665 392072 106218
rect 393240 104854 393268 114514
rect 393228 104848 393280 104854
rect 393228 104790 393280 104796
rect 393136 98728 393188 98734
rect 393136 98670 393188 98676
rect 392030 96656 392086 96665
rect 392030 96591 392086 96600
rect 392214 96656 392270 96665
rect 392214 96591 392270 96600
rect 392228 77382 392256 96591
rect 393148 86850 393176 98670
rect 393148 86822 393268 86850
rect 392216 77376 392268 77382
rect 392216 77318 392268 77324
rect 392124 77308 392176 77314
rect 392124 77250 392176 77256
rect 392136 70258 392164 77250
rect 392136 70230 392256 70258
rect 392228 51134 392256 70230
rect 393240 66230 393268 86822
rect 393228 66224 393280 66230
rect 393228 66166 393280 66172
rect 393136 66156 393188 66162
rect 393136 66098 393188 66104
rect 392216 51128 392268 51134
rect 392216 51070 392268 51076
rect 392124 51060 392176 51066
rect 392124 51002 392176 51008
rect 392136 48278 392164 51002
rect 393148 48346 393176 66098
rect 393320 63844 393372 63850
rect 393320 63786 393372 63792
rect 393332 63753 393360 63786
rect 393318 63744 393374 63753
rect 393318 63679 393374 63688
rect 393136 48340 393188 48346
rect 393136 48282 393188 48288
rect 393228 48340 393280 48346
rect 393228 48282 393280 48288
rect 392124 48272 392176 48278
rect 392124 48214 392176 48220
rect 393240 39114 393268 48282
rect 393148 39086 393268 39114
rect 392216 35964 392268 35970
rect 392216 35906 392268 35912
rect 392228 26246 392256 35906
rect 393148 29034 393176 39086
rect 393136 29028 393188 29034
rect 393136 28970 393188 28976
rect 393228 29028 393280 29034
rect 393228 28970 393280 28976
rect 393240 27606 393268 28970
rect 393228 27600 393280 27606
rect 393228 27542 393280 27548
rect 392216 26240 392268 26246
rect 392216 26182 392268 26188
rect 393228 18012 393280 18018
rect 393228 17954 393280 17960
rect 392216 16652 392268 16658
rect 392216 16594 392268 16600
rect 392228 14686 392256 16594
rect 392032 14680 392084 14686
rect 392032 14622 392084 14628
rect 392216 14680 392268 14686
rect 392216 14622 392268 14628
rect 392044 9246 392072 14622
rect 393240 12510 393268 17954
rect 393228 12504 393280 12510
rect 393228 12446 393280 12452
rect 393044 12436 393096 12442
rect 393044 12378 393096 12384
rect 393056 9654 393084 12378
rect 393044 9648 393096 9654
rect 393044 9590 393096 9596
rect 392032 9240 392084 9246
rect 392032 9182 392084 9188
rect 391940 5500 391992 5506
rect 391940 5442 391992 5448
rect 393516 4554 393544 340054
rect 394804 9110 394832 340054
rect 395264 338026 395292 340068
rect 395356 340054 395922 340082
rect 396184 340054 396566 340082
rect 395252 338020 395304 338026
rect 395252 337962 395304 337968
rect 395356 335730 395384 340054
rect 395436 336932 395488 336938
rect 395436 336874 395488 336880
rect 394896 335702 395384 335730
rect 394792 9104 394844 9110
rect 394792 9046 394844 9052
rect 394240 5364 394292 5370
rect 394240 5306 394292 5312
rect 393504 4548 393556 4554
rect 393504 4490 393556 4496
rect 391204 3936 391256 3942
rect 391204 3878 391256 3884
rect 391848 3664 391900 3670
rect 391848 3606 391900 3612
rect 391860 480 391888 3606
rect 393044 604 393096 610
rect 393044 546 393096 552
rect 393056 480 393084 546
rect 394252 480 394280 5306
rect 394896 4486 394924 335702
rect 395448 331242 395476 336874
rect 395356 331214 395476 331242
rect 394884 4480 394936 4486
rect 394884 4422 394936 4428
rect 395356 3806 395384 331214
rect 395894 29200 395950 29209
rect 396078 29200 396134 29209
rect 395950 29158 396078 29186
rect 395894 29135 395950 29144
rect 396078 29135 396134 29144
rect 396184 7274 396212 340054
rect 397104 337890 397132 340068
rect 397472 340054 397762 340082
rect 397092 337884 397144 337890
rect 397092 337826 397144 337832
rect 396724 336796 396776 336802
rect 396724 336738 396776 336744
rect 396172 7268 396224 7274
rect 396172 7210 396224 7216
rect 396736 3942 396764 336738
rect 397472 280226 397500 340054
rect 397840 328438 397868 340190
rect 398944 336870 398972 340068
rect 399036 340054 399602 340082
rect 398932 336864 398984 336870
rect 398932 336806 398984 336812
rect 397828 328432 397880 328438
rect 397828 328374 397880 328380
rect 397920 318844 397972 318850
rect 397920 318786 397972 318792
rect 397932 311914 397960 318786
rect 397552 311908 397604 311914
rect 397552 311850 397604 311856
rect 397920 311908 397972 311914
rect 397920 311850 397972 311856
rect 397564 302138 397592 311850
rect 397564 302110 397684 302138
rect 397656 299418 397684 302110
rect 397656 299390 397776 299418
rect 397748 298110 397776 299390
rect 397736 298104 397788 298110
rect 397736 298046 397788 298052
rect 397736 288448 397788 288454
rect 397736 288390 397788 288396
rect 397460 280220 397512 280226
rect 397460 280162 397512 280168
rect 397460 280084 397512 280090
rect 397460 280026 397512 280032
rect 397472 4418 397500 280026
rect 397748 278798 397776 288390
rect 397644 278792 397696 278798
rect 397644 278734 397696 278740
rect 397736 278792 397788 278798
rect 397736 278734 397788 278740
rect 397656 278594 397684 278734
rect 397644 278588 397696 278594
rect 397644 278530 397696 278536
rect 397920 269136 397972 269142
rect 397920 269078 397972 269084
rect 397932 260914 397960 269078
rect 397644 260908 397696 260914
rect 397644 260850 397696 260856
rect 397920 260908 397972 260914
rect 397920 260850 397972 260856
rect 397656 259434 397684 260850
rect 397656 259406 397776 259434
rect 397748 253978 397776 259406
rect 397736 253972 397788 253978
rect 397736 253914 397788 253920
rect 397552 249824 397604 249830
rect 397552 249766 397604 249772
rect 397564 245002 397592 249766
rect 397552 244996 397604 245002
rect 397552 244938 397604 244944
rect 397644 240168 397696 240174
rect 397644 240110 397696 240116
rect 397656 234734 397684 240110
rect 397644 234728 397696 234734
rect 397644 234670 397696 234676
rect 397644 234592 397696 234598
rect 397644 234534 397696 234540
rect 397656 227066 397684 234534
rect 397564 227038 397684 227066
rect 397564 215268 397592 227038
rect 397564 215240 397776 215268
rect 397748 202858 397776 215240
rect 397748 202830 397960 202858
rect 397932 193254 397960 202830
rect 397736 193248 397788 193254
rect 397736 193190 397788 193196
rect 397920 193248 397972 193254
rect 397920 193190 397972 193196
rect 397748 176662 397776 193190
rect 397736 176656 397788 176662
rect 397736 176598 397788 176604
rect 397736 173936 397788 173942
rect 397736 173878 397788 173884
rect 397748 164218 397776 173878
rect 397736 164212 397788 164218
rect 397736 164154 397788 164160
rect 397736 154624 397788 154630
rect 397736 154566 397788 154572
rect 397748 144974 397776 154566
rect 397736 144968 397788 144974
rect 397736 144910 397788 144916
rect 397736 143608 397788 143614
rect 397736 143550 397788 143556
rect 397748 124234 397776 143550
rect 397736 124228 397788 124234
rect 397736 124170 397788 124176
rect 397920 124228 397972 124234
rect 397920 124170 397972 124176
rect 397932 115977 397960 124170
rect 397734 115968 397790 115977
rect 397734 115903 397790 115912
rect 397918 115968 397974 115977
rect 397918 115903 397974 115912
rect 397748 114510 397776 115903
rect 397736 114504 397788 114510
rect 397736 114446 397788 114452
rect 397644 104984 397696 104990
rect 397644 104926 397696 104932
rect 397656 104854 397684 104926
rect 397644 104848 397696 104854
rect 397644 104790 397696 104796
rect 397828 104780 397880 104786
rect 397828 104722 397880 104728
rect 397840 99362 397868 104722
rect 397748 99334 397868 99362
rect 397748 80186 397776 99334
rect 397656 80158 397776 80186
rect 397656 80050 397684 80158
rect 397656 80022 397776 80050
rect 397748 56658 397776 80022
rect 398748 76288 398800 76294
rect 398746 76256 398748 76265
rect 398800 76256 398802 76265
rect 398746 76191 398802 76200
rect 397748 56630 397868 56658
rect 397840 56574 397868 56630
rect 397828 56568 397880 56574
rect 397828 56510 397880 56516
rect 397736 46980 397788 46986
rect 397736 46922 397788 46928
rect 397748 22114 397776 46922
rect 397656 22086 397776 22114
rect 397656 19310 397684 22086
rect 397644 19304 397696 19310
rect 397644 19246 397696 19252
rect 397552 9716 397604 9722
rect 397552 9658 397604 9664
rect 397564 7342 397592 9658
rect 397552 7336 397604 7342
rect 397552 7278 397604 7284
rect 397828 5432 397880 5438
rect 397828 5374 397880 5380
rect 397460 4412 397512 4418
rect 397460 4354 397512 4360
rect 396724 3936 396776 3942
rect 396724 3878 396776 3884
rect 395344 3800 395396 3806
rect 395344 3742 395396 3748
rect 396632 3392 396684 3398
rect 396632 3334 396684 3340
rect 395436 2848 395488 2854
rect 395436 2790 395488 2796
rect 395448 480 395476 2790
rect 396644 480 396672 3334
rect 397840 480 397868 5374
rect 399036 4350 399064 340054
rect 400232 338094 400260 340068
rect 400220 338088 400272 338094
rect 400220 338030 400272 338036
rect 400784 336938 400812 340068
rect 400876 340054 401442 340082
rect 401704 340054 402086 340082
rect 400772 336932 400824 336938
rect 400772 336874 400824 336880
rect 400876 335594 400904 340054
rect 401048 336796 401100 336802
rect 401048 336738 401100 336744
rect 400600 335566 400904 335594
rect 400600 328438 400628 335566
rect 401060 331242 401088 336738
rect 400876 331214 401088 331242
rect 400312 328432 400364 328438
rect 400312 328374 400364 328380
rect 400588 328432 400640 328438
rect 400588 328374 400640 328380
rect 400324 327078 400352 328374
rect 400312 327072 400364 327078
rect 400312 327014 400364 327020
rect 400496 318844 400548 318850
rect 400496 318786 400548 318792
rect 400508 315994 400536 318786
rect 400496 315988 400548 315994
rect 400496 315930 400548 315936
rect 400496 299464 400548 299470
rect 400496 299406 400548 299412
rect 400508 282878 400536 299406
rect 400496 282872 400548 282878
rect 400496 282814 400548 282820
rect 400496 282736 400548 282742
rect 400496 282678 400548 282684
rect 400508 273306 400536 282678
rect 400416 273278 400536 273306
rect 400416 273222 400444 273278
rect 400404 273216 400456 273222
rect 400404 273158 400456 273164
rect 400588 273216 400640 273222
rect 400588 273158 400640 273164
rect 400600 270502 400628 273158
rect 400588 270496 400640 270502
rect 400588 270438 400640 270444
rect 400496 260908 400548 260914
rect 400496 260850 400548 260856
rect 400508 253994 400536 260850
rect 400416 253966 400536 253994
rect 400416 253910 400444 253966
rect 400404 253904 400456 253910
rect 400404 253846 400456 253852
rect 400588 253904 400640 253910
rect 400588 253846 400640 253852
rect 400600 251190 400628 253846
rect 400588 251184 400640 251190
rect 400588 251126 400640 251132
rect 400496 241528 400548 241534
rect 400496 241470 400548 241476
rect 400508 234682 400536 241470
rect 400416 234654 400536 234682
rect 400416 234598 400444 234654
rect 400404 234592 400456 234598
rect 400404 234534 400456 234540
rect 400588 234592 400640 234598
rect 400588 234534 400640 234540
rect 400600 231849 400628 234534
rect 400402 231840 400458 231849
rect 400402 231775 400458 231784
rect 400586 231840 400642 231849
rect 400586 231775 400642 231784
rect 400416 222222 400444 231775
rect 400404 222216 400456 222222
rect 400310 222184 400366 222193
rect 400496 222216 400548 222222
rect 400404 222158 400456 222164
rect 400494 222184 400496 222193
rect 400548 222184 400550 222193
rect 400310 222119 400366 222128
rect 400494 222119 400550 222128
rect 400324 212566 400352 222119
rect 400312 212560 400364 212566
rect 400312 212502 400364 212508
rect 400588 212560 400640 212566
rect 400588 212502 400640 212508
rect 400600 205578 400628 212502
rect 400508 205550 400628 205578
rect 400508 202842 400536 205550
rect 400496 202836 400548 202842
rect 400496 202778 400548 202784
rect 400588 202836 400640 202842
rect 400588 202778 400640 202784
rect 400600 167074 400628 202778
rect 400404 167068 400456 167074
rect 400404 167010 400456 167016
rect 400588 167068 400640 167074
rect 400588 167010 400640 167016
rect 400416 166954 400444 167010
rect 400416 166926 400536 166954
rect 400508 164218 400536 166926
rect 400496 164212 400548 164218
rect 400496 164154 400548 164160
rect 400496 157344 400548 157350
rect 400496 157286 400548 157292
rect 400508 154578 400536 157286
rect 400508 154550 400628 154578
rect 400600 147694 400628 154550
rect 400404 147688 400456 147694
rect 400588 147688 400640 147694
rect 400456 147636 400536 147642
rect 400404 147630 400536 147636
rect 400588 147630 400640 147636
rect 400416 147614 400536 147630
rect 400508 144906 400536 147614
rect 400496 144900 400548 144906
rect 400496 144842 400548 144848
rect 400496 137964 400548 137970
rect 400496 137906 400548 137912
rect 400508 135266 400536 137906
rect 400508 135238 400628 135266
rect 400600 125662 400628 135238
rect 400496 125656 400548 125662
rect 400496 125598 400548 125604
rect 400588 125656 400640 125662
rect 400588 125598 400640 125604
rect 400508 116006 400536 125598
rect 400404 116000 400456 116006
rect 400404 115942 400456 115948
rect 400496 116000 400548 116006
rect 400496 115942 400548 115948
rect 400416 111058 400444 115942
rect 400416 111030 400536 111058
rect 400508 104854 400536 111030
rect 400496 104848 400548 104854
rect 400496 104790 400548 104796
rect 400588 95260 400640 95266
rect 400588 95202 400640 95208
rect 400600 67658 400628 95202
rect 400496 67652 400548 67658
rect 400496 67594 400548 67600
rect 400588 67652 400640 67658
rect 400588 67594 400640 67600
rect 400508 60738 400536 67594
rect 400508 60710 400628 60738
rect 400600 47190 400628 60710
rect 400588 47184 400640 47190
rect 400588 47126 400640 47132
rect 400588 45620 400640 45626
rect 400588 45562 400640 45568
rect 400600 45506 400628 45562
rect 400600 45490 400720 45506
rect 400600 45484 400732 45490
rect 400600 45478 400680 45484
rect 400680 45426 400732 45432
rect 400680 37188 400732 37194
rect 400680 37130 400732 37136
rect 400692 28898 400720 37130
rect 400496 28892 400548 28898
rect 400496 28834 400548 28840
rect 400680 28892 400732 28898
rect 400680 28834 400732 28840
rect 400508 12510 400536 28834
rect 400496 12504 400548 12510
rect 400496 12446 400548 12452
rect 400404 12436 400456 12442
rect 400404 12378 400456 12384
rect 399024 4344 399076 4350
rect 399024 4286 399076 4292
rect 400416 4282 400444 12378
rect 400404 4276 400456 4282
rect 400404 4218 400456 4224
rect 400220 3936 400272 3942
rect 400220 3878 400272 3884
rect 399024 3800 399076 3806
rect 399024 3742 399076 3748
rect 399036 480 399064 3742
rect 400232 480 400260 3878
rect 400876 3874 400904 331214
rect 401704 8974 401732 340054
rect 402624 338026 402652 340068
rect 403084 340054 403282 340082
rect 402612 338020 402664 338026
rect 402612 337962 402664 337968
rect 402886 134328 402942 134337
rect 402886 134263 402942 134272
rect 402900 133929 402928 134263
rect 402886 133920 402942 133929
rect 402886 133855 402942 133864
rect 402980 40384 403032 40390
rect 402978 40352 402980 40361
rect 403032 40352 403034 40361
rect 402978 40287 403034 40296
rect 401692 8968 401744 8974
rect 401692 8910 401744 8916
rect 401324 5500 401376 5506
rect 401324 5442 401376 5448
rect 400864 3868 400916 3874
rect 400864 3810 400916 3816
rect 401336 480 401364 5442
rect 403084 4214 403112 340054
rect 403912 337346 403940 340068
rect 403900 337340 403952 337346
rect 403900 337282 403952 337288
rect 404464 336870 404492 340068
rect 404556 340054 405122 340082
rect 405766 340054 405872 340082
rect 404452 336864 404504 336870
rect 404452 336806 404504 336812
rect 404556 4758 404584 340054
rect 405004 337884 405056 337890
rect 405004 337826 405056 337832
rect 404544 4752 404596 4758
rect 404544 4694 404596 4700
rect 404912 4752 404964 4758
rect 404912 4694 404964 4700
rect 403072 4208 403124 4214
rect 403072 4150 403124 4156
rect 402520 3868 402572 3874
rect 402520 3810 402572 3816
rect 403716 3868 403768 3874
rect 403716 3810 403768 3816
rect 402532 480 402560 3810
rect 403728 480 403756 3810
rect 404924 480 404952 4694
rect 405016 4214 405044 337826
rect 405740 157752 405792 157758
rect 405738 157720 405740 157729
rect 405792 157720 405794 157729
rect 405738 157655 405794 157664
rect 405646 134328 405702 134337
rect 405702 134286 405780 134314
rect 405646 134263 405702 134272
rect 405752 134201 405780 134286
rect 405738 134192 405794 134201
rect 405738 134127 405794 134136
rect 405648 76288 405700 76294
rect 405646 76256 405648 76265
rect 405700 76256 405702 76265
rect 405646 76191 405702 76200
rect 405646 63880 405702 63889
rect 405646 63815 405648 63824
rect 405700 63815 405702 63824
rect 405648 63786 405700 63792
rect 405738 16960 405794 16969
rect 405738 16895 405794 16904
rect 405752 16833 405780 16895
rect 405738 16824 405794 16833
rect 405738 16759 405794 16768
rect 405844 7614 405872 340054
rect 406304 337822 406332 340068
rect 406672 340054 406962 340082
rect 406292 337816 406344 337822
rect 406292 337758 406344 337764
rect 406672 335646 406700 340054
rect 407500 337278 407528 340068
rect 407764 337952 407816 337958
rect 407764 337894 407816 337900
rect 407488 337272 407540 337278
rect 407488 337214 407540 337220
rect 405924 335640 405976 335646
rect 405924 335582 405976 335588
rect 406660 335640 406712 335646
rect 406660 335582 406712 335588
rect 405832 7608 405884 7614
rect 405832 7550 405884 7556
rect 405936 4690 405964 335582
rect 407776 251190 407804 337894
rect 408144 336802 408172 340068
rect 408512 340054 408802 340082
rect 408132 336796 408184 336802
rect 408132 336738 408184 336744
rect 407672 251184 407724 251190
rect 407672 251126 407724 251132
rect 407764 251184 407816 251190
rect 407764 251126 407816 251132
rect 407684 249801 407712 251126
rect 407486 249792 407542 249801
rect 407486 249727 407542 249736
rect 407670 249792 407726 249801
rect 407670 249727 407726 249736
rect 407500 240174 407528 249727
rect 407488 240168 407540 240174
rect 407488 240110 407540 240116
rect 407764 240168 407816 240174
rect 407764 240110 407816 240116
rect 407776 124166 407804 240110
rect 408408 164212 408460 164218
rect 408408 164154 408460 164160
rect 408420 154601 408448 164154
rect 408406 154592 408462 154601
rect 408406 154527 408462 154536
rect 407764 124160 407816 124166
rect 407764 124102 407816 124108
rect 407764 114572 407816 114578
rect 407764 114514 407816 114520
rect 407776 104854 407804 114514
rect 407764 104848 407816 104854
rect 407764 104790 407816 104796
rect 407856 87032 407908 87038
rect 407776 86980 407856 86986
rect 407776 86974 407908 86980
rect 407776 86958 407896 86974
rect 407776 85542 407804 86958
rect 407764 85536 407816 85542
rect 407764 85478 407816 85484
rect 407764 75948 407816 75954
rect 407764 75890 407816 75896
rect 407776 66230 407804 75890
rect 407764 66224 407816 66230
rect 407764 66166 407816 66172
rect 407764 56636 407816 56642
rect 407764 56578 407816 56584
rect 407776 46918 407804 56578
rect 407764 46912 407816 46918
rect 407764 46854 407816 46860
rect 407764 37324 407816 37330
rect 407764 37266 407816 37272
rect 407776 27606 407804 37266
rect 407764 27600 407816 27606
rect 407764 27542 407816 27548
rect 407856 9716 407908 9722
rect 407856 9658 407908 9664
rect 405924 4684 405976 4690
rect 405924 4626 405976 4632
rect 407868 4282 407896 9658
rect 408512 4826 408540 340054
rect 408880 331242 408908 340190
rect 409788 337816 409840 337822
rect 409788 337758 409840 337764
rect 409144 337272 409196 337278
rect 409144 337214 409196 337220
rect 408696 331214 408908 331242
rect 408696 321638 408724 331214
rect 408684 321632 408736 321638
rect 408684 321574 408736 321580
rect 408776 321496 408828 321502
rect 408776 321438 408828 321444
rect 408788 315994 408816 321438
rect 408776 315988 408828 315994
rect 408776 315930 408828 315936
rect 408776 302116 408828 302122
rect 408776 302058 408828 302064
rect 408788 292670 408816 302058
rect 408776 292664 408828 292670
rect 408776 292606 408828 292612
rect 408684 292528 408736 292534
rect 408684 292470 408736 292476
rect 408696 288386 408724 292470
rect 408684 288380 408736 288386
rect 408684 288322 408736 288328
rect 408776 278792 408828 278798
rect 408776 278734 408828 278740
rect 408788 273358 408816 278734
rect 408776 273352 408828 273358
rect 408776 273294 408828 273300
rect 408684 273216 408736 273222
rect 408684 273158 408736 273164
rect 408696 263634 408724 273158
rect 408684 263628 408736 263634
rect 408684 263570 408736 263576
rect 408776 263492 408828 263498
rect 408776 263434 408828 263440
rect 408788 258058 408816 263434
rect 408776 258052 408828 258058
rect 408776 257994 408828 258000
rect 408960 258052 409012 258058
rect 408960 257994 409012 258000
rect 408972 248441 409000 257994
rect 408774 248432 408830 248441
rect 408774 248367 408830 248376
rect 408958 248432 409014 248441
rect 408958 248367 409014 248376
rect 408788 229106 408816 248367
rect 408696 229078 408816 229106
rect 408696 224942 408724 229078
rect 408684 224936 408736 224942
rect 408684 224878 408736 224884
rect 408868 224936 408920 224942
rect 408868 224878 408920 224884
rect 408880 222170 408908 224878
rect 408788 222142 408908 222170
rect 408788 215354 408816 222142
rect 408776 215348 408828 215354
rect 408776 215290 408828 215296
rect 408776 212560 408828 212566
rect 408776 212502 408828 212508
rect 408788 205578 408816 212502
rect 408696 205550 408816 205578
rect 408696 202881 408724 205550
rect 408682 202872 408738 202881
rect 408682 202807 408738 202816
rect 408958 202872 409014 202881
rect 408958 202807 409014 202816
rect 408972 193254 409000 202807
rect 408776 193248 408828 193254
rect 408776 193190 408828 193196
rect 408960 193248 409012 193254
rect 408960 193190 409012 193196
rect 408788 186266 408816 193190
rect 408696 186238 408816 186266
rect 408696 183569 408724 186238
rect 408682 183560 408738 183569
rect 408682 183495 408738 183504
rect 408958 183560 409014 183569
rect 408958 183495 409014 183504
rect 408972 173942 409000 183495
rect 408776 173936 408828 173942
rect 408776 173878 408828 173884
rect 408960 173936 409012 173942
rect 408960 173878 409012 173884
rect 408788 166954 408816 173878
rect 408604 166926 408816 166954
rect 408604 164218 408632 166926
rect 408592 164212 408644 164218
rect 408592 164154 408644 164160
rect 408682 154592 408738 154601
rect 408682 154527 408738 154536
rect 408696 147642 408724 154527
rect 408696 147614 408908 147642
rect 408880 140078 408908 147614
rect 408868 140072 408920 140078
rect 408868 140014 408920 140020
rect 409052 140072 409104 140078
rect 409052 140014 409104 140020
rect 409064 135289 409092 140014
rect 408866 135280 408922 135289
rect 408866 135215 408922 135224
rect 409050 135280 409106 135289
rect 409050 135215 409106 135224
rect 408880 125769 408908 135215
rect 408866 125760 408922 125769
rect 408866 125695 408922 125704
rect 408682 125624 408738 125633
rect 408682 125559 408738 125568
rect 408696 119354 408724 125559
rect 408604 119326 408724 119354
rect 408604 114646 408632 119326
rect 408592 114640 408644 114646
rect 408592 114582 408644 114588
rect 408776 114640 408828 114646
rect 408776 114582 408828 114588
rect 408788 114510 408816 114582
rect 408776 114504 408828 114510
rect 408776 114446 408828 114452
rect 408684 104916 408736 104922
rect 408684 104858 408736 104864
rect 408696 104802 408724 104858
rect 408696 104774 408816 104802
rect 408788 100094 408816 104774
rect 408776 100088 408828 100094
rect 408776 100030 408828 100036
rect 408776 89684 408828 89690
rect 408776 89626 408828 89632
rect 408788 86986 408816 89626
rect 408788 86958 408908 86986
rect 408880 85542 408908 86958
rect 408868 85536 408920 85542
rect 408868 85478 408920 85484
rect 408684 76016 408736 76022
rect 408684 75958 408736 75964
rect 408696 75886 408724 75958
rect 408684 75880 408736 75886
rect 408684 75822 408736 75828
rect 408776 66292 408828 66298
rect 408776 66234 408828 66240
rect 408788 66178 408816 66234
rect 408696 66150 408816 66178
rect 408696 60738 408724 66150
rect 408696 60710 408816 60738
rect 408788 56658 408816 60710
rect 408696 56630 408816 56658
rect 408696 51134 408724 56630
rect 408684 51128 408736 51134
rect 408684 51070 408736 51076
rect 408776 51060 408828 51066
rect 408776 51002 408828 51008
rect 408788 47002 408816 51002
rect 408696 46974 408816 47002
rect 408696 45558 408724 46974
rect 408684 45552 408736 45558
rect 408684 45494 408736 45500
rect 408776 45552 408828 45558
rect 408776 45494 408828 45500
rect 408788 31822 408816 45494
rect 408776 31816 408828 31822
rect 408776 31758 408828 31764
rect 408684 31748 408736 31754
rect 408684 31690 408736 31696
rect 408696 27577 408724 31690
rect 408682 27568 408738 27577
rect 408682 27503 408738 27512
rect 408774 27432 408830 27441
rect 408774 27367 408830 27376
rect 408788 6866 408816 27367
rect 408776 6860 408828 6866
rect 408776 6802 408828 6808
rect 408500 4820 408552 4826
rect 408500 4762 408552 4768
rect 407856 4276 407908 4282
rect 407856 4218 407908 4224
rect 405004 4208 405056 4214
rect 405004 4150 405056 4156
rect 408408 4072 408460 4078
rect 408408 4014 408460 4020
rect 408316 3664 408368 3670
rect 408314 3632 408316 3641
rect 408368 3632 408370 3641
rect 408314 3567 408370 3576
rect 408420 3466 408448 4014
rect 409156 4010 409184 337214
rect 409144 4004 409196 4010
rect 409144 3946 409196 3952
rect 408592 3664 408644 3670
rect 408590 3632 408592 3641
rect 408644 3632 408646 3641
rect 408590 3567 408646 3576
rect 409800 3466 409828 337758
rect 409984 337754 410012 340068
rect 410076 340054 410642 340082
rect 409972 337748 410024 337754
rect 409972 337690 410024 337696
rect 410076 4894 410104 340054
rect 411180 337346 411208 340068
rect 411824 337890 411852 340068
rect 411916 340054 412482 340082
rect 411812 337884 411864 337890
rect 411812 337826 411864 337832
rect 411168 337340 411220 337346
rect 411168 337282 411220 337288
rect 410616 336864 410668 336870
rect 410616 336806 410668 336812
rect 410524 336796 410576 336802
rect 410524 336738 410576 336744
rect 410064 4888 410116 4894
rect 410064 4830 410116 4836
rect 408408 3460 408460 3466
rect 408408 3402 408460 3408
rect 408500 3460 408552 3466
rect 408500 3402 408552 3408
rect 409788 3460 409840 3466
rect 409788 3402 409840 3408
rect 407304 3392 407356 3398
rect 407304 3334 407356 3340
rect 406108 3324 406160 3330
rect 406108 3266 406160 3272
rect 406120 480 406148 3266
rect 407316 480 407344 3334
rect 408512 480 408540 3402
rect 409696 3392 409748 3398
rect 410536 3369 410564 336738
rect 409696 3334 409748 3340
rect 410522 3360 410578 3369
rect 408592 3052 408644 3058
rect 408592 2994 408644 3000
rect 408604 2922 408632 2994
rect 408592 2916 408644 2922
rect 408592 2858 408644 2864
rect 409708 480 409736 3334
rect 410522 3295 410578 3304
rect 410628 3126 410656 336806
rect 411916 335594 411944 340054
rect 412088 338088 412140 338094
rect 412088 338030 412140 338036
rect 411364 335566 411944 335594
rect 411364 6050 411392 335566
rect 412100 331242 412128 338030
rect 412548 337748 412600 337754
rect 412548 337690 412600 337696
rect 411916 331214 412128 331242
rect 411352 6044 411404 6050
rect 411352 5986 411404 5992
rect 410892 4072 410944 4078
rect 410892 4014 410944 4020
rect 410616 3120 410668 3126
rect 410616 3062 410668 3068
rect 410904 480 410932 4014
rect 411916 3262 411944 331214
rect 412454 40488 412510 40497
rect 412454 40423 412510 40432
rect 412468 40390 412496 40423
rect 412456 40384 412508 40390
rect 412456 40326 412508 40332
rect 412560 4146 412588 337690
rect 413020 336802 413048 340068
rect 413284 337884 413336 337890
rect 413284 337826 413336 337832
rect 413008 336796 413060 336802
rect 413008 336738 413060 336744
rect 412088 4140 412140 4146
rect 412088 4082 412140 4088
rect 412548 4140 412600 4146
rect 412548 4082 412600 4088
rect 411904 3256 411956 3262
rect 411904 3198 411956 3204
rect 412100 480 412128 4082
rect 413296 3058 413324 337826
rect 413468 337272 413520 337278
rect 413468 337214 413520 337220
rect 413376 336932 413428 336938
rect 413376 336874 413428 336880
rect 413388 4078 413416 336874
rect 413376 4072 413428 4078
rect 413376 4014 413428 4020
rect 413284 3052 413336 3058
rect 413284 2994 413336 3000
rect 413376 3052 413428 3058
rect 413376 2994 413428 3000
rect 413388 1714 413416 2994
rect 413480 2990 413508 337214
rect 413664 337142 413692 340068
rect 414124 340054 414322 340082
rect 413652 337136 413704 337142
rect 413652 337078 413704 337084
rect 413926 40488 413982 40497
rect 413926 40423 413982 40432
rect 413940 40225 413968 40423
rect 413926 40216 413982 40225
rect 413926 40151 413982 40160
rect 414124 4962 414152 340054
rect 414664 337136 414716 337142
rect 414664 337078 414716 337084
rect 414112 4956 414164 4962
rect 414112 4898 414164 4904
rect 414676 4146 414704 337078
rect 414860 337074 414888 340068
rect 415504 337958 415532 340068
rect 415596 340054 416162 340082
rect 416424 340054 416714 340082
rect 415492 337952 415544 337958
rect 415492 337894 415544 337900
rect 414848 337068 414900 337074
rect 414848 337010 414900 337016
rect 415308 157752 415360 157758
rect 415306 157720 415308 157729
rect 415360 157720 415362 157729
rect 415306 157655 415362 157664
rect 415398 87136 415454 87145
rect 415398 87071 415400 87080
rect 415452 87071 415454 87080
rect 415400 87042 415452 87048
rect 415596 5914 415624 340054
rect 416136 337884 416188 337890
rect 416136 337826 416188 337832
rect 416044 336796 416096 336802
rect 416044 336738 416096 336744
rect 415584 5908 415636 5914
rect 415584 5850 415636 5856
rect 414664 4140 414716 4146
rect 414664 4082 414716 4088
rect 415676 4140 415728 4146
rect 415676 4082 415728 4088
rect 414480 4072 414532 4078
rect 414480 4014 414532 4020
rect 413468 2984 413520 2990
rect 413468 2926 413520 2932
rect 413296 1686 413416 1714
rect 413296 480 413324 1686
rect 414492 480 414520 4014
rect 415688 480 415716 4082
rect 416056 2922 416084 336738
rect 416148 4078 416176 337826
rect 416424 336870 416452 340054
rect 416688 338020 416740 338026
rect 416688 337962 416740 337968
rect 416412 336864 416464 336870
rect 416412 336806 416464 336812
rect 416700 4146 416728 337962
rect 417344 337006 417372 340068
rect 417436 340054 418002 340082
rect 417332 337000 417384 337006
rect 417332 336942 417384 336948
rect 417436 335594 417464 340054
rect 418540 337686 418568 340068
rect 419184 338094 419212 340068
rect 419644 340054 419842 340082
rect 419172 338088 419224 338094
rect 419172 338030 419224 338036
rect 418528 337680 418580 337686
rect 418528 337622 418580 337628
rect 417608 337204 417660 337210
rect 417608 337146 417660 337152
rect 416792 335566 417464 335594
rect 416792 331226 416820 335566
rect 417620 334234 417648 337146
rect 417436 334206 417648 334234
rect 416780 331220 416832 331226
rect 416780 331162 416832 331168
rect 416964 331220 417016 331226
rect 416964 331162 417016 331168
rect 416976 328438 417004 331162
rect 416964 328432 417016 328438
rect 416964 328374 417016 328380
rect 416872 318844 416924 318850
rect 416872 318786 416924 318792
rect 416884 311930 416912 318786
rect 416792 311902 416912 311930
rect 416792 311846 416820 311902
rect 416780 311840 416832 311846
rect 416780 311782 416832 311788
rect 416964 311840 417016 311846
rect 416964 311782 417016 311788
rect 416976 309126 417004 311782
rect 416964 309120 417016 309126
rect 416964 309062 417016 309068
rect 416872 299532 416924 299538
rect 416872 299474 416924 299480
rect 416884 294658 416912 299474
rect 416884 294630 417004 294658
rect 416976 282826 417004 294630
rect 416884 282798 417004 282826
rect 416884 280158 416912 282798
rect 416872 280152 416924 280158
rect 416872 280094 416924 280100
rect 416964 270564 417016 270570
rect 416964 270506 417016 270512
rect 416976 263514 417004 270506
rect 416884 263486 417004 263514
rect 416884 260846 416912 263486
rect 416872 260840 416924 260846
rect 416872 260782 416924 260788
rect 416964 251252 417016 251258
rect 416964 251194 417016 251200
rect 416976 244202 417004 251194
rect 416884 244174 417004 244202
rect 416884 241505 416912 244174
rect 416870 241496 416926 241505
rect 416870 241431 416926 241440
rect 417146 241496 417202 241505
rect 417146 241431 417202 241440
rect 417160 231878 417188 241431
rect 416964 231872 417016 231878
rect 416964 231814 417016 231820
rect 417148 231872 417200 231878
rect 417148 231814 417200 231820
rect 416976 224890 417004 231814
rect 416884 224862 417004 224890
rect 416884 222193 416912 224862
rect 416870 222184 416926 222193
rect 416870 222119 416926 222128
rect 417146 222184 417202 222193
rect 417146 222119 417202 222128
rect 417160 212566 417188 222119
rect 416964 212560 417016 212566
rect 416964 212502 417016 212508
rect 417148 212560 417200 212566
rect 417148 212502 417200 212508
rect 416976 205578 417004 212502
rect 416884 205550 417004 205578
rect 416884 202881 416912 205550
rect 416870 202872 416926 202881
rect 416870 202807 416926 202816
rect 417146 202872 417202 202881
rect 417146 202807 417202 202816
rect 417160 193254 417188 202807
rect 416964 193248 417016 193254
rect 416964 193190 417016 193196
rect 417148 193248 417200 193254
rect 417148 193190 417200 193196
rect 416976 186266 417004 193190
rect 416884 186238 417004 186266
rect 416884 183530 416912 186238
rect 416872 183524 416924 183530
rect 416872 183466 416924 183472
rect 416964 183524 417016 183530
rect 416964 183466 417016 183472
rect 416976 166954 417004 183466
rect 416884 166926 417004 166954
rect 416884 164218 416912 166926
rect 416872 164212 416924 164218
rect 416872 164154 416924 164160
rect 416964 164212 417016 164218
rect 416964 164154 417016 164160
rect 416976 147642 417004 164154
rect 416884 147614 417004 147642
rect 416884 138038 416912 147614
rect 416872 138032 416924 138038
rect 416872 137974 416924 137980
rect 416780 137964 416832 137970
rect 416780 137906 416832 137912
rect 416792 135289 416820 137906
rect 416778 135280 416834 135289
rect 416778 135215 416834 135224
rect 416962 135280 417018 135289
rect 416962 135215 417018 135224
rect 416976 128330 417004 135215
rect 416884 128302 417004 128330
rect 416884 118726 416912 128302
rect 416872 118720 416924 118726
rect 416872 118662 416924 118668
rect 416780 118652 416832 118658
rect 416780 118594 416832 118600
rect 416792 115977 416820 118594
rect 416778 115968 416834 115977
rect 416778 115903 416834 115912
rect 416962 115968 417018 115977
rect 416962 115903 417018 115912
rect 416976 109018 417004 115903
rect 416884 108990 417004 109018
rect 416884 99414 416912 108990
rect 416872 99408 416924 99414
rect 416872 99350 416924 99356
rect 416780 99340 416832 99346
rect 416780 99282 416832 99288
rect 416792 96665 416820 99282
rect 416778 96656 416834 96665
rect 416778 96591 416834 96600
rect 416962 96656 417018 96665
rect 416962 96591 417018 96600
rect 416976 89706 417004 96591
rect 416884 89678 417004 89706
rect 416884 77382 416912 89678
rect 416872 77376 416924 77382
rect 416872 77318 416924 77324
rect 416964 77376 417016 77382
rect 416964 77318 417016 77324
rect 416976 70514 417004 77318
rect 416964 70508 417016 70514
rect 416964 70450 417016 70456
rect 416872 70372 416924 70378
rect 416872 70314 416924 70320
rect 416884 67590 416912 70314
rect 416872 67584 416924 67590
rect 416872 67526 416924 67532
rect 417056 67584 417108 67590
rect 417056 67526 417108 67532
rect 417068 58018 417096 67526
rect 416976 57990 417096 58018
rect 416976 57934 417004 57990
rect 416964 57928 417016 57934
rect 416964 57870 417016 57876
rect 416872 48408 416924 48414
rect 416872 48350 416924 48356
rect 416884 48278 416912 48350
rect 416872 48272 416924 48278
rect 416872 48214 416924 48220
rect 417056 48272 417108 48278
rect 417056 48214 417108 48220
rect 417068 38706 417096 48214
rect 416976 38678 417096 38706
rect 416976 31822 417004 38678
rect 416964 31816 417016 31822
rect 416964 31758 417016 31764
rect 416872 31748 416924 31754
rect 416872 31690 416924 31696
rect 416884 22114 416912 31690
rect 416792 22098 416912 22114
rect 416780 22092 416912 22098
rect 416832 22086 416912 22092
rect 416964 22092 417016 22098
rect 416780 22034 416832 22040
rect 416964 22034 417016 22040
rect 416976 11966 417004 22034
rect 416964 11960 417016 11966
rect 416964 11902 417016 11908
rect 416964 11824 417016 11830
rect 416964 11766 417016 11772
rect 416976 5030 417004 11766
rect 416964 5024 417016 5030
rect 416964 4966 417016 4972
rect 416688 4140 416740 4146
rect 416688 4082 416740 4088
rect 416136 4072 416188 4078
rect 416136 4014 416188 4020
rect 417436 3330 417464 334206
rect 418066 204504 418122 204513
rect 418066 204439 418122 204448
rect 418080 204105 418108 204439
rect 418066 204096 418122 204105
rect 418066 204031 418122 204040
rect 418066 169960 418122 169969
rect 418066 169895 418122 169904
rect 418080 169561 418108 169895
rect 418066 169552 418122 169561
rect 418066 169487 418122 169496
rect 417882 134328 417938 134337
rect 417882 134263 417938 134272
rect 417896 134178 417924 134263
rect 418250 134192 418306 134201
rect 417896 134150 418250 134178
rect 418250 134127 418306 134136
rect 418066 110664 418122 110673
rect 418066 110599 418122 110608
rect 418080 110265 418108 110599
rect 418066 110256 418122 110265
rect 418066 110191 418122 110200
rect 418066 76256 418122 76265
rect 418066 76191 418122 76200
rect 418080 76106 418108 76191
rect 418158 76120 418214 76129
rect 418080 76078 418158 76106
rect 418158 76055 418214 76064
rect 418066 63880 418122 63889
rect 418066 63815 418122 63824
rect 418080 63730 418108 63815
rect 418158 63744 418214 63753
rect 418080 63702 418158 63730
rect 418158 63679 418214 63688
rect 418066 16960 418122 16969
rect 418250 16960 418306 16969
rect 418122 16918 418250 16946
rect 418066 16895 418122 16904
rect 418250 16895 418306 16904
rect 419644 5846 419672 340054
rect 420276 338088 420328 338094
rect 420276 338030 420328 338036
rect 420184 337068 420236 337074
rect 420184 337010 420236 337016
rect 419632 5840 419684 5846
rect 419632 5782 419684 5788
rect 419172 4140 419224 4146
rect 419172 4082 419224 4088
rect 416780 3324 416832 3330
rect 416780 3266 416832 3272
rect 417424 3324 417476 3330
rect 417424 3266 417476 3272
rect 417976 3324 418028 3330
rect 417976 3266 418028 3272
rect 416792 3126 416820 3266
rect 416780 3120 416832 3126
rect 416780 3062 416832 3068
rect 416872 3120 416924 3126
rect 416872 3062 416924 3068
rect 416044 2916 416096 2922
rect 416044 2858 416096 2864
rect 416884 480 416912 3062
rect 417988 480 418016 3266
rect 419184 480 419212 4082
rect 420196 2854 420224 337010
rect 420288 4146 420316 338030
rect 420380 337958 420408 340068
rect 420368 337952 420420 337958
rect 420368 337894 420420 337900
rect 420828 337680 420880 337686
rect 420828 337622 420880 337628
rect 420840 4146 420868 337622
rect 421024 337414 421052 340068
rect 421116 340054 421682 340082
rect 421012 337408 421064 337414
rect 421012 337350 421064 337356
rect 421116 6186 421144 340054
rect 422220 337482 422248 340068
rect 422208 337476 422260 337482
rect 422208 337418 422260 337424
rect 422208 337272 422260 337278
rect 422208 337214 422260 337220
rect 422116 22568 422168 22574
rect 422116 22510 422168 22516
rect 422128 9722 422156 22510
rect 422116 9716 422168 9722
rect 422116 9658 422168 9664
rect 421104 6180 421156 6186
rect 421104 6122 421156 6128
rect 422220 4146 422248 337214
rect 422864 337142 422892 340068
rect 423232 340054 423522 340082
rect 422852 337136 422904 337142
rect 422852 337078 422904 337084
rect 423232 335646 423260 340054
rect 424060 337210 424088 340068
rect 424244 340054 424718 340082
rect 425164 340054 425270 340082
rect 424048 337204 424100 337210
rect 424048 337146 424100 337152
rect 423588 337136 423640 337142
rect 423588 337078 423640 337084
rect 422300 335640 422352 335646
rect 422300 335582 422352 335588
rect 423220 335640 423272 335646
rect 423220 335582 423272 335588
rect 422312 331226 422340 335582
rect 422300 331220 422352 331226
rect 422300 331162 422352 331168
rect 422484 331220 422536 331226
rect 422484 331162 422536 331168
rect 422496 328438 422524 331162
rect 422484 328432 422536 328438
rect 422484 328374 422536 328380
rect 422392 318844 422444 318850
rect 422392 318786 422444 318792
rect 422404 311930 422432 318786
rect 422312 311902 422432 311930
rect 422312 311846 422340 311902
rect 422300 311840 422352 311846
rect 422300 311782 422352 311788
rect 422484 311840 422536 311846
rect 422484 311782 422536 311788
rect 422496 309126 422524 311782
rect 422484 309120 422536 309126
rect 422484 309062 422536 309068
rect 422484 299940 422536 299946
rect 422484 299882 422536 299888
rect 422496 282946 422524 299882
rect 422300 282940 422352 282946
rect 422300 282882 422352 282888
rect 422484 282940 422536 282946
rect 422484 282882 422536 282888
rect 422312 282826 422340 282882
rect 422312 282798 422432 282826
rect 422404 273306 422432 282798
rect 422404 273278 422524 273306
rect 422496 263634 422524 273278
rect 422300 263628 422352 263634
rect 422300 263570 422352 263576
rect 422484 263628 422536 263634
rect 422484 263570 422536 263576
rect 422312 263514 422340 263570
rect 422312 263486 422432 263514
rect 422404 253994 422432 263486
rect 422404 253966 422524 253994
rect 422496 244322 422524 253966
rect 422300 244316 422352 244322
rect 422300 244258 422352 244264
rect 422484 244316 422536 244322
rect 422484 244258 422536 244264
rect 422312 244202 422340 244258
rect 422312 244174 422432 244202
rect 422404 234682 422432 244174
rect 422404 234654 422524 234682
rect 422496 225010 422524 234654
rect 422300 225004 422352 225010
rect 422300 224946 422352 224952
rect 422484 225004 422536 225010
rect 422484 224946 422536 224952
rect 422312 224890 422340 224946
rect 422312 224862 422432 224890
rect 422404 215370 422432 224862
rect 422404 215342 422524 215370
rect 422496 205698 422524 215342
rect 422300 205692 422352 205698
rect 422300 205634 422352 205640
rect 422484 205692 422536 205698
rect 422484 205634 422536 205640
rect 422312 205578 422340 205634
rect 422312 205550 422432 205578
rect 422404 196058 422432 205550
rect 422404 196030 422524 196058
rect 422496 186386 422524 196030
rect 422300 186380 422352 186386
rect 422300 186322 422352 186328
rect 422484 186380 422536 186386
rect 422484 186322 422536 186328
rect 422312 186266 422340 186322
rect 422312 186238 422432 186266
rect 422404 183569 422432 186238
rect 422390 183560 422446 183569
rect 422390 183495 422446 183504
rect 422666 183560 422722 183569
rect 422666 183495 422722 183504
rect 422680 173942 422708 183495
rect 422484 173936 422536 173942
rect 422484 173878 422536 173884
rect 422668 173936 422720 173942
rect 422668 173878 422720 173884
rect 422496 167074 422524 173878
rect 422300 167068 422352 167074
rect 422300 167010 422352 167016
rect 422484 167068 422536 167074
rect 422484 167010 422536 167016
rect 422312 166954 422340 167010
rect 422312 166926 422432 166954
rect 422404 164218 422432 166926
rect 422392 164212 422444 164218
rect 422392 164154 422444 164160
rect 422392 157344 422444 157350
rect 422392 157286 422444 157292
rect 422404 154578 422432 157286
rect 422404 154550 422524 154578
rect 422496 147694 422524 154550
rect 422300 147688 422352 147694
rect 422484 147688 422536 147694
rect 422352 147636 422432 147642
rect 422300 147630 422432 147636
rect 422484 147630 422536 147636
rect 422312 147614 422432 147630
rect 422404 144906 422432 147614
rect 422392 144900 422444 144906
rect 422392 144842 422444 144848
rect 422392 137964 422444 137970
rect 422392 137906 422444 137912
rect 422404 135266 422432 137906
rect 422404 135238 422524 135266
rect 422496 128382 422524 135238
rect 422300 128376 422352 128382
rect 422484 128376 422536 128382
rect 422352 128324 422432 128330
rect 422300 128318 422432 128324
rect 422484 128318 422536 128324
rect 422312 128302 422432 128318
rect 422404 118726 422432 128302
rect 422392 118720 422444 118726
rect 422392 118662 422444 118668
rect 422484 118652 422536 118658
rect 422484 118594 422536 118600
rect 422496 109070 422524 118594
rect 422300 109064 422352 109070
rect 422484 109064 422536 109070
rect 422352 109012 422432 109018
rect 422300 109006 422432 109012
rect 422484 109006 422536 109012
rect 422312 108990 422432 109006
rect 422404 106282 422432 108990
rect 422392 106276 422444 106282
rect 422392 106218 422444 106224
rect 422392 99340 422444 99346
rect 422392 99282 422444 99288
rect 422404 96642 422432 99282
rect 422404 96614 422524 96642
rect 422496 89758 422524 96614
rect 422300 89752 422352 89758
rect 422484 89752 422536 89758
rect 422352 89700 422432 89706
rect 422300 89694 422432 89700
rect 422484 89694 422536 89700
rect 422312 89678 422432 89694
rect 422404 86970 422432 89678
rect 422392 86964 422444 86970
rect 422392 86906 422444 86912
rect 422484 77308 422536 77314
rect 422484 77250 422536 77256
rect 422496 67658 422524 77250
rect 422392 67652 422444 67658
rect 422392 67594 422444 67600
rect 422484 67652 422536 67658
rect 422484 67594 422536 67600
rect 422404 60738 422432 67594
rect 422404 60710 422524 60738
rect 422496 48346 422524 60710
rect 422392 48340 422444 48346
rect 422392 48282 422444 48288
rect 422484 48340 422536 48346
rect 422484 48282 422536 48288
rect 422404 41426 422432 48282
rect 422404 41398 422524 41426
rect 422496 27674 422524 41398
rect 422392 27668 422444 27674
rect 422392 27610 422444 27616
rect 422484 27668 422536 27674
rect 422484 27610 422536 27616
rect 422404 22574 422432 27610
rect 422392 22568 422444 22574
rect 422392 22510 422444 22516
rect 422392 9716 422444 9722
rect 422392 9658 422444 9664
rect 422404 5098 422432 9658
rect 422392 5092 422444 5098
rect 422392 5034 422444 5040
rect 423600 4146 423628 337078
rect 424244 336802 424272 340054
rect 424968 337272 425020 337278
rect 424968 337214 425020 337220
rect 424416 337000 424468 337006
rect 424416 336942 424468 336948
rect 424232 336796 424284 336802
rect 424232 336738 424284 336744
rect 424324 336796 424376 336802
rect 424324 336738 424376 336744
rect 420276 4140 420328 4146
rect 420276 4082 420328 4088
rect 420368 4140 420420 4146
rect 420368 4082 420420 4088
rect 420828 4140 420880 4146
rect 420828 4082 420880 4088
rect 421564 4140 421616 4146
rect 421564 4082 421616 4088
rect 422208 4140 422260 4146
rect 422208 4082 422260 4088
rect 422760 4140 422812 4146
rect 422760 4082 422812 4088
rect 423588 4140 423640 4146
rect 423588 4082 423640 4088
rect 420184 2848 420236 2854
rect 420184 2790 420236 2796
rect 420380 480 420408 4082
rect 421576 480 421604 4082
rect 422772 480 422800 4082
rect 424336 3398 424364 336738
rect 424428 4010 424456 336942
rect 424784 87100 424836 87106
rect 424784 87042 424836 87048
rect 424796 86986 424824 87042
rect 424874 87000 424930 87009
rect 424796 86958 424874 86986
rect 424874 86935 424930 86944
rect 424416 4004 424468 4010
rect 424416 3946 424468 3952
rect 424324 3392 424376 3398
rect 424324 3334 424376 3340
rect 424980 3262 425008 337214
rect 425060 204400 425112 204406
rect 425058 204368 425060 204377
rect 425112 204368 425114 204377
rect 425058 204303 425114 204312
rect 425060 180872 425112 180878
rect 425058 180840 425060 180849
rect 425112 180840 425114 180849
rect 425058 180775 425114 180784
rect 425060 169856 425112 169862
rect 425058 169824 425060 169833
rect 425112 169824 425114 169833
rect 425058 169759 425114 169768
rect 425060 122936 425112 122942
rect 425058 122904 425060 122913
rect 425112 122904 425114 122913
rect 425058 122839 425114 122848
rect 425060 110560 425112 110566
rect 425058 110528 425060 110537
rect 425112 110528 425114 110537
rect 425058 110463 425114 110472
rect 425060 87032 425112 87038
rect 425058 87000 425060 87009
rect 425112 87000 425114 87009
rect 425058 86935 425114 86944
rect 425164 6254 425192 340054
rect 425900 336802 425928 340068
rect 426558 340054 426664 340082
rect 425888 336796 425940 336802
rect 425888 336738 425940 336744
rect 425152 6248 425204 6254
rect 425152 6190 425204 6196
rect 426636 3670 426664 340054
rect 426728 340054 427110 340082
rect 426728 5166 426756 340054
rect 427084 336932 427136 336938
rect 427084 336874 427136 336880
rect 426716 5160 426768 5166
rect 426716 5102 426768 5108
rect 426624 3664 426676 3670
rect 426624 3606 426676 3612
rect 426348 3528 426400 3534
rect 426348 3470 426400 3476
rect 425152 3392 425204 3398
rect 425152 3334 425204 3340
rect 423956 3256 424008 3262
rect 423956 3198 424008 3204
rect 424968 3256 425020 3262
rect 424968 3198 425020 3204
rect 423968 480 423996 3198
rect 425164 480 425192 3334
rect 426360 480 426388 3470
rect 427096 2990 427124 336874
rect 427740 336870 427768 340068
rect 428384 337346 428412 340068
rect 428476 340054 428950 340082
rect 428372 337340 428424 337346
rect 428372 337282 428424 337288
rect 427728 336864 427780 336870
rect 427728 336806 427780 336812
rect 428476 334354 428504 340054
rect 429580 337414 429608 340068
rect 429764 340054 430238 340082
rect 430684 340054 430790 340082
rect 431144 340054 431434 340082
rect 429568 337408 429620 337414
rect 429568 337350 429620 337356
rect 428556 337340 428608 337346
rect 428556 337282 428608 337288
rect 428004 334348 428056 334354
rect 428004 334290 428056 334296
rect 428464 334348 428516 334354
rect 428464 334290 428516 334296
rect 428016 328438 428044 334290
rect 428568 334234 428596 337282
rect 429108 336864 429160 336870
rect 429108 336806 429160 336812
rect 428476 334206 428596 334234
rect 428004 328432 428056 328438
rect 428004 328374 428056 328380
rect 427912 318844 427964 318850
rect 427912 318786 427964 318792
rect 427924 311930 427952 318786
rect 427832 311902 427952 311930
rect 427832 311846 427860 311902
rect 427820 311840 427872 311846
rect 427820 311782 427872 311788
rect 428004 311840 428056 311846
rect 428004 311782 428056 311788
rect 428016 309126 428044 311782
rect 428004 309120 428056 309126
rect 428004 309062 428056 309068
rect 428004 299532 428056 299538
rect 428004 299474 428056 299480
rect 428016 282946 428044 299474
rect 427820 282940 427872 282946
rect 427820 282882 427872 282888
rect 428004 282940 428056 282946
rect 428004 282882 428056 282888
rect 427832 282826 427860 282882
rect 427832 282798 427952 282826
rect 427924 273306 427952 282798
rect 427924 273278 428044 273306
rect 428016 263634 428044 273278
rect 427820 263628 427872 263634
rect 427820 263570 427872 263576
rect 428004 263628 428056 263634
rect 428004 263570 428056 263576
rect 427832 263514 427860 263570
rect 427832 263486 427952 263514
rect 427924 253994 427952 263486
rect 427924 253966 428044 253994
rect 428016 244322 428044 253966
rect 427820 244316 427872 244322
rect 427820 244258 427872 244264
rect 428004 244316 428056 244322
rect 428004 244258 428056 244264
rect 427832 244202 427860 244258
rect 427832 244174 427952 244202
rect 427924 234682 427952 244174
rect 427924 234654 428044 234682
rect 428016 225010 428044 234654
rect 427820 225004 427872 225010
rect 427820 224946 427872 224952
rect 428004 225004 428056 225010
rect 428004 224946 428056 224952
rect 427832 224890 427860 224946
rect 427832 224862 427952 224890
rect 427924 215370 427952 224862
rect 427924 215342 428044 215370
rect 428016 205698 428044 215342
rect 427820 205692 427872 205698
rect 427820 205634 427872 205640
rect 428004 205692 428056 205698
rect 428004 205634 428056 205640
rect 427832 205578 427860 205634
rect 427832 205550 428044 205578
rect 428016 186386 428044 205550
rect 427820 186380 427872 186386
rect 427820 186322 427872 186328
rect 428004 186380 428056 186386
rect 428004 186322 428056 186328
rect 427832 186266 427860 186322
rect 427832 186238 427952 186266
rect 427924 167090 427952 186238
rect 427832 167062 427952 167090
rect 427832 166954 427860 167062
rect 427832 166926 427952 166954
rect 427924 147778 427952 166926
rect 427832 147750 427952 147778
rect 427832 147642 427860 147750
rect 427832 147614 428044 147642
rect 428016 144906 428044 147614
rect 427728 144900 427780 144906
rect 427728 144842 427780 144848
rect 428004 144900 428056 144906
rect 428004 144842 428056 144848
rect 427740 135289 427768 144842
rect 427726 135280 427782 135289
rect 427726 135215 427782 135224
rect 427910 135280 427966 135289
rect 427910 135215 427966 135224
rect 427924 128466 427952 135215
rect 427832 128438 427952 128466
rect 427832 128330 427860 128438
rect 427832 128302 427952 128330
rect 427924 109154 427952 128302
rect 427832 109126 427952 109154
rect 427832 109018 427860 109126
rect 427832 108990 427952 109018
rect 427924 106282 427952 108990
rect 427912 106276 427964 106282
rect 427912 106218 427964 106224
rect 427912 99340 427964 99346
rect 427912 99282 427964 99288
rect 427924 96642 427952 99282
rect 427924 96614 428044 96642
rect 428016 89758 428044 96614
rect 427820 89752 427872 89758
rect 428004 89752 428056 89758
rect 427872 89700 427952 89706
rect 427820 89694 427952 89700
rect 428004 89694 428056 89700
rect 427832 89678 427952 89694
rect 427924 76362 427952 89678
rect 427912 76356 427964 76362
rect 427912 76298 427964 76304
rect 428004 67652 428056 67658
rect 428004 67594 428056 67600
rect 428016 51082 428044 67594
rect 427832 51054 428044 51082
rect 427832 50946 427860 51054
rect 427832 50918 427952 50946
rect 427924 31906 427952 50918
rect 427924 31878 428044 31906
rect 428016 29050 428044 31878
rect 427924 29022 428044 29050
rect 427924 28966 427952 29022
rect 427912 28960 427964 28966
rect 427912 28902 427964 28908
rect 427820 19440 427872 19446
rect 427820 19382 427872 19388
rect 427832 19310 427860 19382
rect 427820 19304 427872 19310
rect 427820 19246 427872 19252
rect 427912 9716 427964 9722
rect 427912 9658 427964 9664
rect 427924 5234 427952 9658
rect 427912 5228 427964 5234
rect 427912 5170 427964 5176
rect 427544 4004 427596 4010
rect 427544 3946 427596 3952
rect 427084 2984 427136 2990
rect 427084 2926 427136 2932
rect 427556 480 427584 3946
rect 428476 3534 428504 334206
rect 428464 3528 428516 3534
rect 428464 3470 428516 3476
rect 429120 626 429148 336806
rect 429764 331242 429792 340054
rect 430488 336796 430540 336802
rect 430488 336738 430540 336744
rect 429304 331214 429792 331242
rect 429304 3670 429332 331214
rect 430500 4146 430528 336738
rect 430580 335640 430632 335646
rect 430580 335582 430632 335588
rect 430592 4146 430620 335582
rect 430684 5302 430712 340054
rect 431144 335646 431172 340054
rect 432064 337618 432092 340068
rect 432156 340054 432630 340082
rect 432052 337612 432104 337618
rect 432052 337554 432104 337560
rect 431868 337068 431920 337074
rect 431868 337010 431920 337016
rect 431224 337000 431276 337006
rect 431224 336942 431276 336948
rect 431132 335640 431184 335646
rect 431132 335582 431184 335588
rect 430672 5296 430724 5302
rect 430672 5238 430724 5244
rect 429936 4140 429988 4146
rect 429936 4082 429988 4088
rect 430488 4140 430540 4146
rect 430488 4082 430540 4088
rect 430580 4140 430632 4146
rect 430580 4082 430632 4088
rect 431132 4140 431184 4146
rect 431132 4082 431184 4088
rect 429292 3664 429344 3670
rect 429292 3606 429344 3612
rect 428752 598 429148 626
rect 428752 480 428780 598
rect 429948 480 429976 4082
rect 431144 480 431172 4082
rect 431236 3194 431264 336942
rect 431880 4146 431908 337010
rect 432156 5370 432184 340054
rect 432604 337544 432656 337550
rect 432604 337486 432656 337492
rect 432144 5364 432196 5370
rect 432144 5306 432196 5312
rect 431868 4140 431920 4146
rect 431868 4082 431920 4088
rect 432420 3936 432472 3942
rect 432616 3890 432644 337486
rect 433260 337210 433288 340068
rect 433352 340054 433918 340082
rect 434180 340054 434470 340082
rect 434824 340054 435114 340082
rect 433248 337204 433300 337210
rect 433248 337146 433300 337152
rect 432472 3884 432644 3890
rect 432420 3878 432644 3884
rect 432432 3862 432644 3878
rect 433352 3738 433380 340054
rect 434180 328681 434208 340054
rect 434628 337000 434680 337006
rect 434628 336942 434680 336948
rect 434166 328672 434222 328681
rect 434166 328607 434222 328616
rect 433706 328536 433762 328545
rect 433706 328471 433762 328480
rect 433720 328438 433748 328471
rect 433708 328432 433760 328438
rect 433708 328374 433760 328380
rect 433800 318844 433852 318850
rect 433800 318786 433852 318792
rect 433812 311914 433840 318786
rect 433432 311908 433484 311914
rect 433432 311850 433484 311856
rect 433800 311908 433852 311914
rect 433800 311850 433852 311856
rect 433444 309126 433472 311850
rect 433432 309120 433484 309126
rect 433432 309062 433484 309068
rect 433708 299532 433760 299538
rect 433708 299474 433760 299480
rect 433720 285002 433748 299474
rect 433628 284974 433748 285002
rect 433628 280158 433656 284974
rect 433616 280152 433668 280158
rect 433616 280094 433668 280100
rect 433708 270564 433760 270570
rect 433708 270506 433760 270512
rect 433720 263514 433748 270506
rect 433628 263486 433748 263514
rect 433628 260846 433656 263486
rect 433616 260840 433668 260846
rect 433616 260782 433668 260788
rect 433708 251252 433760 251258
rect 433708 251194 433760 251200
rect 433720 244202 433748 251194
rect 433628 244174 433748 244202
rect 433628 241505 433656 244174
rect 433430 241496 433486 241505
rect 433430 241431 433486 241440
rect 433614 241496 433670 241505
rect 433614 241431 433670 241440
rect 433444 231878 433472 241431
rect 433432 231872 433484 231878
rect 433432 231814 433484 231820
rect 433708 231872 433760 231878
rect 433708 231814 433760 231820
rect 433720 224890 433748 231814
rect 433628 224862 433748 224890
rect 433628 222193 433656 224862
rect 433430 222184 433486 222193
rect 433430 222119 433486 222128
rect 433614 222184 433670 222193
rect 433614 222119 433670 222128
rect 433444 212566 433472 222119
rect 433432 212560 433484 212566
rect 433432 212502 433484 212508
rect 433708 212560 433760 212566
rect 433708 212502 433760 212508
rect 433720 196110 433748 212502
rect 434534 204640 434590 204649
rect 434534 204575 434590 204584
rect 434548 204406 434576 204575
rect 434536 204400 434588 204406
rect 434536 204342 434588 204348
rect 433708 196104 433760 196110
rect 433708 196046 433760 196052
rect 433708 193248 433760 193254
rect 433708 193190 433760 193196
rect 433720 173942 433748 193190
rect 434534 181112 434590 181121
rect 434534 181047 434590 181056
rect 434548 180878 434576 181047
rect 434536 180872 434588 180878
rect 434536 180814 434588 180820
rect 433616 173936 433668 173942
rect 433616 173878 433668 173884
rect 433708 173936 433760 173942
rect 433708 173878 433760 173884
rect 433628 157434 433656 173878
rect 434534 170096 434590 170105
rect 434534 170031 434590 170040
rect 434548 169862 434576 170031
rect 434536 169856 434588 169862
rect 434536 169798 434588 169804
rect 433536 157406 433656 157434
rect 433536 157298 433564 157406
rect 433536 157270 433656 157298
rect 433628 147762 433656 157270
rect 433616 147756 433668 147762
rect 433616 147698 433668 147704
rect 433616 147620 433668 147626
rect 433616 147562 433668 147568
rect 433628 125594 433656 147562
rect 433616 125588 433668 125594
rect 433616 125530 433668 125536
rect 434534 123176 434590 123185
rect 434534 123111 434590 123120
rect 434548 122942 434576 123111
rect 434536 122936 434588 122942
rect 434536 122878 434588 122884
rect 433616 116000 433668 116006
rect 433616 115942 433668 115948
rect 433628 106282 433656 115942
rect 434534 110800 434590 110809
rect 434534 110735 434590 110744
rect 434548 110566 434576 110735
rect 434536 110560 434588 110566
rect 434536 110502 434588 110508
rect 433616 106276 433668 106282
rect 433616 106218 433668 106224
rect 433616 99340 433668 99346
rect 433616 99282 433668 99288
rect 433628 96642 433656 99282
rect 433628 96614 433748 96642
rect 433720 80238 433748 96614
rect 434534 87272 434590 87281
rect 434534 87207 434590 87216
rect 434548 87038 434576 87207
rect 434536 87032 434588 87038
rect 434536 86974 434588 86980
rect 433708 80232 433760 80238
rect 433708 80174 433760 80180
rect 433616 77308 433668 77314
rect 433616 77250 433668 77256
rect 433628 60738 433656 77250
rect 433536 60722 433656 60738
rect 433524 60716 433656 60722
rect 433576 60710 433656 60716
rect 433708 60716 433760 60722
rect 433524 60658 433576 60664
rect 433708 60658 433760 60664
rect 433720 57934 433748 60658
rect 433708 57928 433760 57934
rect 433708 57870 433760 57876
rect 433616 48340 433668 48346
rect 433616 48282 433668 48288
rect 433628 41426 433656 48282
rect 433536 41398 433656 41426
rect 433536 41290 433564 41398
rect 433536 41262 433656 41290
rect 433628 22114 433656 41262
rect 433536 22086 433656 22114
rect 433536 21978 433564 22086
rect 433536 21950 433656 21978
rect 433628 5438 433656 21950
rect 433616 5432 433668 5438
rect 433616 5374 433668 5380
rect 434640 4146 434668 336942
rect 433524 4140 433576 4146
rect 433524 4082 433576 4088
rect 434628 4140 434680 4146
rect 434628 4082 434680 4088
rect 433340 3732 433392 3738
rect 433340 3674 433392 3680
rect 432328 3392 432380 3398
rect 432328 3334 432380 3340
rect 431224 3188 431276 3194
rect 431224 3130 431276 3136
rect 432340 480 432368 3334
rect 433536 480 433564 4082
rect 434824 3806 434852 340054
rect 435744 337550 435772 340068
rect 436204 340054 436310 340082
rect 435732 337544 435784 337550
rect 435732 337486 435784 337492
rect 436008 337068 436060 337074
rect 436008 337010 436060 337016
rect 435364 336864 435416 336870
rect 435364 336806 435416 336812
rect 434812 3800 434864 3806
rect 434812 3742 434864 3748
rect 434536 3732 434588 3738
rect 434536 3674 434588 3680
rect 434548 1850 434576 3674
rect 435376 3194 435404 336806
rect 435364 3188 435416 3194
rect 435364 3130 435416 3136
rect 434548 1822 434668 1850
rect 434640 480 434668 1822
rect 436020 610 436048 337010
rect 436204 5506 436232 340054
rect 436940 337822 436968 340068
rect 437598 340054 437704 340082
rect 436928 337816 436980 337822
rect 436928 337758 436980 337764
rect 437480 337816 437532 337822
rect 437480 337758 437532 337764
rect 437492 336802 437520 337758
rect 437480 336796 437532 336802
rect 437480 336738 437532 336744
rect 436192 5500 436244 5506
rect 436192 5442 436244 5448
rect 437020 4140 437072 4146
rect 437020 4082 437072 4088
rect 435824 604 435876 610
rect 435824 546 435876 552
rect 436008 604 436060 610
rect 436008 546 436060 552
rect 435836 480 435864 546
rect 437032 480 437060 4082
rect 437676 3874 437704 340054
rect 437768 340054 438150 340082
rect 437768 4758 437796 340054
rect 438780 337822 438808 340068
rect 438964 340054 439438 340082
rect 438768 337816 438820 337822
rect 438768 337758 438820 337764
rect 438124 336796 438176 336802
rect 438124 336738 438176 336744
rect 437756 4752 437808 4758
rect 437756 4694 437808 4700
rect 437664 3868 437716 3874
rect 437664 3810 437716 3816
rect 438136 3126 438164 336738
rect 438964 4078 438992 340054
rect 439976 337958 440004 340068
rect 439964 337952 440016 337958
rect 439964 337894 440016 337900
rect 440620 336938 440648 340068
rect 441264 337618 441292 340068
rect 441816 337754 441844 340068
rect 442264 337952 442316 337958
rect 442264 337894 442316 337900
rect 441804 337748 441856 337754
rect 441804 337690 441856 337696
rect 441252 337612 441304 337618
rect 441252 337554 441304 337560
rect 440608 336932 440660 336938
rect 440608 336874 440660 336880
rect 438952 4072 439004 4078
rect 438952 4014 439004 4020
rect 440608 4072 440660 4078
rect 440608 4014 440660 4020
rect 438216 3800 438268 3806
rect 438216 3742 438268 3748
rect 438124 3120 438176 3126
rect 438124 3062 438176 3068
rect 438228 480 438256 3742
rect 439412 3596 439464 3602
rect 439412 3538 439464 3544
rect 439424 480 439452 3538
rect 440620 480 440648 4014
rect 442276 3942 442304 337894
rect 442356 337748 442408 337754
rect 442356 337690 442408 337696
rect 442368 4146 442396 337690
rect 442460 336870 442488 340068
rect 443012 337890 443040 340068
rect 443656 338026 443684 340068
rect 443644 338020 443696 338026
rect 443644 337962 443696 337968
rect 443000 337884 443052 337890
rect 443000 337826 443052 337832
rect 442448 336864 442500 336870
rect 442448 336806 442500 336812
rect 444300 336802 444328 340068
rect 444576 340054 444866 340082
rect 444288 336796 444340 336802
rect 444288 336738 444340 336744
rect 442356 4140 442408 4146
rect 442356 4082 442408 4088
rect 442264 3936 442316 3942
rect 442264 3878 442316 3884
rect 443000 3664 443052 3670
rect 443000 3606 443052 3612
rect 441804 3324 441856 3330
rect 441804 3266 441856 3272
rect 441816 480 441844 3266
rect 443012 480 443040 3606
rect 444576 3466 444604 340054
rect 445496 338094 445524 340068
rect 445484 338088 445536 338094
rect 445484 338030 445536 338036
rect 445024 337816 445076 337822
rect 445024 337758 445076 337764
rect 445036 4078 445064 337758
rect 446140 337686 446168 340068
rect 446416 340054 446706 340082
rect 446128 337680 446180 337686
rect 446128 337622 446180 337628
rect 446416 337482 446444 340054
rect 446404 337476 446456 337482
rect 446404 337418 446456 337424
rect 446496 337476 446548 337482
rect 446496 337418 446548 337424
rect 446404 336796 446456 336802
rect 446404 336738 446456 336744
rect 445024 4072 445076 4078
rect 445024 4014 445076 4020
rect 445392 4072 445444 4078
rect 445392 4014 445444 4020
rect 444564 3460 444616 3466
rect 444564 3402 444616 3408
rect 444196 3120 444248 3126
rect 444196 3062 444248 3068
rect 444208 480 444236 3062
rect 445404 480 445432 4014
rect 446416 3738 446444 336738
rect 446404 3732 446456 3738
rect 446404 3674 446456 3680
rect 446508 3126 446536 337418
rect 447336 337414 447364 340068
rect 447324 337408 447376 337414
rect 447324 337350 447376 337356
rect 447980 337278 448008 340068
rect 447968 337272 448020 337278
rect 447968 337214 448020 337220
rect 448428 337272 448480 337278
rect 448428 337214 448480 337220
rect 447784 336796 447836 336802
rect 447784 336738 447836 336744
rect 447796 3806 447824 336738
rect 447784 3800 447836 3806
rect 447784 3742 447836 3748
rect 446588 3460 446640 3466
rect 446588 3402 446640 3408
rect 446496 3120 446548 3126
rect 446496 3062 446548 3068
rect 446600 480 446628 3402
rect 448440 3330 448468 337214
rect 448532 4010 448560 340068
rect 449176 337210 449204 340068
rect 449820 337958 449848 340068
rect 449808 337952 449860 337958
rect 449808 337894 449860 337900
rect 449256 337884 449308 337890
rect 449256 337826 449308 337832
rect 449164 337204 449216 337210
rect 449164 337146 449216 337152
rect 449268 334506 449296 337826
rect 450372 337346 450400 340068
rect 451016 337550 451044 340068
rect 451004 337544 451056 337550
rect 451004 337486 451056 337492
rect 451188 337544 451240 337550
rect 451188 337486 451240 337492
rect 450360 337340 450412 337346
rect 450360 337282 450412 337288
rect 449176 334478 449296 334506
rect 448520 4004 448572 4010
rect 448520 3946 448572 3952
rect 448980 3868 449032 3874
rect 448980 3810 449032 3816
rect 447784 3324 447836 3330
rect 447784 3266 447836 3272
rect 448428 3324 448480 3330
rect 448428 3266 448480 3272
rect 447796 480 447824 3266
rect 448992 480 449020 3810
rect 449176 3398 449204 334478
rect 451200 3738 451228 337486
rect 451660 337142 451688 340068
rect 451844 340054 452226 340082
rect 451648 337136 451700 337142
rect 451648 337078 451700 337084
rect 451844 335345 451872 340054
rect 451924 338020 451976 338026
rect 451924 337962 451976 337968
rect 451370 335336 451426 335345
rect 451370 335271 451426 335280
rect 451830 335336 451886 335345
rect 451830 335271 451886 335280
rect 451384 325718 451412 335271
rect 451372 325712 451424 325718
rect 451556 325712 451608 325718
rect 451372 325654 451424 325660
rect 451554 325680 451556 325689
rect 451608 325680 451610 325689
rect 451554 325615 451610 325624
rect 451738 325680 451794 325689
rect 451738 325615 451794 325624
rect 451752 316130 451780 325615
rect 451556 316124 451608 316130
rect 451556 316066 451608 316072
rect 451740 316124 451792 316130
rect 451740 316066 451792 316072
rect 451568 315994 451596 316066
rect 451556 315988 451608 315994
rect 451556 315930 451608 315936
rect 451556 302116 451608 302122
rect 451556 302058 451608 302064
rect 451568 292670 451596 302058
rect 451556 292664 451608 292670
rect 451556 292606 451608 292612
rect 451464 292528 451516 292534
rect 451464 292470 451516 292476
rect 451476 288425 451504 292470
rect 451278 288416 451334 288425
rect 451278 288351 451334 288360
rect 451462 288416 451518 288425
rect 451462 288351 451518 288360
rect 451292 278798 451320 288351
rect 451280 278792 451332 278798
rect 451280 278734 451332 278740
rect 451556 278792 451608 278798
rect 451556 278734 451608 278740
rect 451568 273766 451596 278734
rect 451556 273760 451608 273766
rect 451556 273702 451608 273708
rect 451556 263492 451608 263498
rect 451556 263434 451608 263440
rect 451568 259418 451596 263434
rect 451556 259412 451608 259418
rect 451556 259354 451608 259360
rect 451556 244180 451608 244186
rect 451556 244122 451608 244128
rect 451568 234734 451596 244122
rect 451556 234728 451608 234734
rect 451556 234670 451608 234676
rect 451464 234592 451516 234598
rect 451464 234534 451516 234540
rect 451476 231826 451504 234534
rect 451384 231798 451504 231826
rect 451384 225010 451412 231798
rect 451372 225004 451424 225010
rect 451372 224946 451424 224952
rect 451280 222216 451332 222222
rect 451278 222184 451280 222193
rect 451332 222184 451334 222193
rect 451278 222119 451334 222128
rect 451738 222048 451794 222057
rect 451738 221983 451794 221992
rect 451752 205578 451780 221983
rect 451660 205550 451780 205578
rect 451660 196058 451688 205550
rect 451568 196030 451688 196058
rect 451568 195922 451596 196030
rect 451568 195894 451688 195922
rect 451660 186522 451688 195894
rect 451648 186516 451700 186522
rect 451648 186458 451700 186464
rect 451648 186380 451700 186386
rect 451648 186322 451700 186328
rect 451660 182186 451688 186322
rect 451660 182158 451780 182186
rect 451752 172514 451780 182158
rect 451740 172508 451792 172514
rect 451740 172450 451792 172456
rect 451830 162888 451886 162897
rect 451752 162858 451830 162874
rect 451740 162852 451830 162858
rect 451792 162846 451830 162852
rect 451830 162823 451886 162832
rect 451740 162794 451792 162800
rect 451556 147620 451608 147626
rect 451556 147562 451608 147568
rect 451568 138038 451596 147562
rect 451556 138032 451608 138038
rect 451556 137974 451608 137980
rect 451740 137964 451792 137970
rect 451740 137906 451792 137912
rect 451752 128382 451780 137906
rect 451556 128376 451608 128382
rect 451740 128376 451792 128382
rect 451608 128324 451740 128330
rect 451556 128318 451792 128324
rect 451568 128302 451780 128318
rect 451752 118794 451780 128302
rect 451740 118788 451792 118794
rect 451740 118730 451792 118736
rect 451740 118652 451792 118658
rect 451740 118594 451792 118600
rect 451752 115954 451780 118594
rect 451752 115926 451872 115954
rect 451844 109018 451872 115926
rect 451660 108990 451872 109018
rect 451660 99521 451688 108990
rect 451646 99512 451702 99521
rect 451646 99447 451702 99456
rect 451646 96656 451702 96665
rect 451646 96591 451702 96600
rect 451660 46986 451688 96591
rect 451372 46980 451424 46986
rect 451372 46922 451424 46928
rect 451648 46980 451700 46986
rect 451648 46922 451700 46928
rect 451384 41342 451412 46922
rect 451372 41336 451424 41342
rect 451372 41278 451424 41284
rect 451740 41336 451792 41342
rect 451740 41278 451792 41284
rect 451752 31822 451780 41278
rect 451740 31816 451792 31822
rect 451740 31758 451792 31764
rect 451648 31748 451700 31754
rect 451648 31690 451700 31696
rect 451660 22114 451688 31690
rect 451660 22086 451780 22114
rect 451752 12458 451780 22086
rect 451568 12430 451780 12458
rect 451280 4140 451332 4146
rect 451280 4082 451332 4088
rect 450176 3732 450228 3738
rect 450176 3674 450228 3680
rect 451188 3732 451240 3738
rect 451188 3674 451240 3680
rect 449164 3392 449216 3398
rect 449164 3334 449216 3340
rect 450188 480 450216 3674
rect 451292 480 451320 4082
rect 451568 3262 451596 12430
rect 451936 4078 451964 337962
rect 452856 337618 452884 340068
rect 453396 337952 453448 337958
rect 453396 337894 453448 337900
rect 452844 337612 452896 337618
rect 452844 337554 452896 337560
rect 453304 337408 453356 337414
rect 453304 337350 453356 337356
rect 452016 172508 452068 172514
rect 452016 172450 452068 172456
rect 452028 162897 452056 172450
rect 452014 162888 452070 162897
rect 452014 162823 452070 162832
rect 451924 4072 451976 4078
rect 451924 4014 451976 4020
rect 453316 3874 453344 337350
rect 453408 4146 453436 337894
rect 453500 336938 453528 340068
rect 453948 337612 454000 337618
rect 453948 337554 454000 337560
rect 453488 336932 453540 336938
rect 453488 336874 453540 336880
rect 453396 4140 453448 4146
rect 453396 4082 453448 4088
rect 453304 3868 453356 3874
rect 453304 3810 453356 3816
rect 452476 3528 452528 3534
rect 452476 3470 452528 3476
rect 451556 3256 451608 3262
rect 451556 3198 451608 3204
rect 452488 480 452516 3470
rect 453960 610 453988 337554
rect 454052 337074 454080 340068
rect 454696 337754 454724 340068
rect 454684 337748 454736 337754
rect 454684 337690 454736 337696
rect 454040 337068 454092 337074
rect 454040 337010 454092 337016
rect 455340 336802 455368 340068
rect 455616 340054 455906 340082
rect 455328 336796 455380 336802
rect 455328 336738 455380 336744
rect 454040 169992 454092 169998
rect 454038 169960 454040 169969
rect 454092 169960 454094 169969
rect 454038 169895 454094 169904
rect 454040 123072 454092 123078
rect 454038 123040 454040 123049
rect 454092 123040 454094 123049
rect 454038 122975 454094 122984
rect 454868 4072 454920 4078
rect 454868 4014 454920 4020
rect 453672 604 453724 610
rect 453672 546 453724 552
rect 453948 604 454000 610
rect 453948 546 454000 552
rect 453684 480 453712 546
rect 454880 480 454908 4014
rect 455616 3602 455644 340054
rect 456536 337822 456564 340068
rect 457180 337890 457208 340068
rect 457168 337884 457220 337890
rect 457168 337826 457220 337832
rect 456524 337816 456576 337822
rect 456524 337758 456576 337764
rect 456064 337680 456116 337686
rect 456064 337622 456116 337628
rect 456076 4078 456104 337622
rect 457272 331242 457300 340190
rect 458376 337482 458404 340068
rect 459020 338026 459048 340068
rect 459586 340054 459784 340082
rect 459008 338020 459060 338026
rect 459008 337962 459060 337968
rect 458364 337476 458416 337482
rect 458364 337418 458416 337424
rect 456996 331214 457300 331242
rect 456706 157584 456762 157593
rect 456890 157584 456946 157593
rect 456762 157542 456890 157570
rect 456706 157519 456762 157528
rect 456890 157519 456946 157528
rect 456706 134056 456762 134065
rect 456890 134056 456946 134065
rect 456762 134014 456890 134042
rect 456706 133991 456762 134000
rect 456890 133991 456946 134000
rect 456706 76120 456762 76129
rect 456890 76120 456946 76129
rect 456762 76078 456890 76106
rect 456706 76055 456762 76064
rect 456890 76055 456946 76064
rect 456706 63744 456762 63753
rect 456890 63744 456946 63753
rect 456762 63702 456890 63730
rect 456706 63679 456762 63688
rect 456890 63679 456946 63688
rect 456706 40216 456762 40225
rect 456890 40216 456946 40225
rect 456762 40174 456890 40202
rect 456706 40151 456762 40160
rect 456890 40151 456946 40160
rect 456706 16824 456762 16833
rect 456890 16824 456946 16833
rect 456762 16782 456890 16810
rect 456706 16759 456762 16768
rect 456890 16759 456946 16768
rect 456064 4072 456116 4078
rect 456064 4014 456116 4020
rect 456156 4004 456208 4010
rect 456156 3946 456208 3952
rect 455604 3596 455656 3602
rect 455604 3538 455656 3544
rect 456168 1986 456196 3946
rect 456996 3670 457024 331214
rect 458180 169992 458232 169998
rect 458178 169960 458180 169969
rect 458232 169960 458234 169969
rect 458178 169895 458234 169904
rect 458180 123072 458232 123078
rect 458178 123040 458180 123049
rect 458232 123040 458234 123049
rect 458178 122975 458234 122984
rect 459652 3800 459704 3806
rect 459652 3742 459704 3748
rect 456984 3664 457036 3670
rect 456984 3606 457036 3612
rect 458456 3664 458508 3670
rect 458456 3606 458508 3612
rect 457260 3596 457312 3602
rect 457260 3538 457312 3544
rect 456076 1958 456196 1986
rect 456076 480 456104 1958
rect 457272 480 457300 3538
rect 458468 480 458496 3606
rect 459664 480 459692 3742
rect 459756 3466 459784 340054
rect 460216 337278 460244 340068
rect 460768 337414 460796 340068
rect 461412 337550 461440 340068
rect 462056 337958 462084 340068
rect 462044 337952 462096 337958
rect 462044 337894 462096 337900
rect 461400 337544 461452 337550
rect 461400 337486 461452 337492
rect 460756 337408 460808 337414
rect 460756 337350 460808 337356
rect 460848 337408 460900 337414
rect 460848 337350 460900 337356
rect 460204 337272 460256 337278
rect 460204 337214 460256 337220
rect 460204 336796 460256 336802
rect 460204 336738 460256 336744
rect 460216 3534 460244 336738
rect 460204 3528 460256 3534
rect 460204 3470 460256 3476
rect 459744 3460 459796 3466
rect 459744 3402 459796 3408
rect 460860 480 460888 337350
rect 462608 336802 462636 340068
rect 463252 337618 463280 340068
rect 463608 337816 463660 337822
rect 463608 337758 463660 337764
rect 463240 337612 463292 337618
rect 463240 337554 463292 337560
rect 462964 336932 463016 336938
rect 462964 336874 463016 336880
rect 462596 336796 462648 336802
rect 462596 336738 462648 336744
rect 462976 4010 463004 336874
rect 462964 4004 463016 4010
rect 462964 3946 463016 3952
rect 463620 3346 463648 337758
rect 463896 337686 463924 340068
rect 463884 337680 463936 337686
rect 463884 337622 463936 337628
rect 464344 337000 464396 337006
rect 464344 336942 464396 336948
rect 464356 3806 464384 336942
rect 464448 336938 464476 340068
rect 464436 336932 464488 336938
rect 464436 336874 464488 336880
rect 464988 336864 465040 336870
rect 464988 336806 465040 336812
rect 464436 336796 464488 336802
rect 464436 336738 464488 336744
rect 464344 3800 464396 3806
rect 464344 3742 464396 3748
rect 464448 3670 464476 336738
rect 464436 3664 464488 3670
rect 464436 3606 464488 3612
rect 463252 3318 463648 3346
rect 465000 3330 465028 336806
rect 465092 3602 465120 340068
rect 465736 336802 465764 340068
rect 466288 337006 466316 340068
rect 466368 337680 466420 337686
rect 466368 337622 466420 337628
rect 466276 337000 466328 337006
rect 466276 336942 466328 336948
rect 465724 336796 465776 336802
rect 465724 336738 465776 336744
rect 466276 29232 466328 29238
rect 466276 29174 466328 29180
rect 466288 29073 466316 29174
rect 466274 29064 466330 29073
rect 466274 28999 466330 29008
rect 465080 3596 465132 3602
rect 465080 3538 465132 3544
rect 466380 3534 466408 337622
rect 466932 337414 466960 340068
rect 467116 340054 467590 340082
rect 466920 337408 466972 337414
rect 466920 337350 466972 337356
rect 467116 333334 467144 340054
rect 468128 337822 468156 340068
rect 468116 337816 468168 337822
rect 468116 337758 468168 337764
rect 468772 336938 468800 340068
rect 469416 337686 469444 340068
rect 469404 337680 469456 337686
rect 469404 337622 469456 337628
rect 468760 336932 468812 336938
rect 468760 336874 468812 336880
rect 469968 336870 469996 340068
rect 470626 340054 470732 340082
rect 467748 336864 467800 336870
rect 467748 336806 467800 336812
rect 469956 336864 470008 336870
rect 469956 336806 470008 336812
rect 466552 333328 466604 333334
rect 466552 333270 466604 333276
rect 467104 333328 467156 333334
rect 467104 333270 467156 333276
rect 466564 321638 466592 333270
rect 466552 321632 466604 321638
rect 466552 321574 466604 321580
rect 466552 318844 466604 318850
rect 466552 318786 466604 318792
rect 466564 311930 466592 318786
rect 466472 311902 466592 311930
rect 466472 311846 466500 311902
rect 466460 311840 466512 311846
rect 466460 311782 466512 311788
rect 466644 311840 466696 311846
rect 466644 311782 466696 311788
rect 466656 309126 466684 311782
rect 466644 309120 466696 309126
rect 466644 309062 466696 309068
rect 466552 299532 466604 299538
rect 466552 299474 466604 299480
rect 466564 292618 466592 299474
rect 466472 292590 466592 292618
rect 466472 292534 466500 292590
rect 466460 292528 466512 292534
rect 466460 292470 466512 292476
rect 466644 292528 466696 292534
rect 466644 292470 466696 292476
rect 466656 280242 466684 292470
rect 466564 280214 466684 280242
rect 466564 280158 466592 280214
rect 466552 280152 466604 280158
rect 466552 280094 466604 280100
rect 466644 270564 466696 270570
rect 466644 270506 466696 270512
rect 466656 263514 466684 270506
rect 466564 263486 466684 263514
rect 466564 260846 466592 263486
rect 466552 260840 466604 260846
rect 466552 260782 466604 260788
rect 466644 251252 466696 251258
rect 466644 251194 466696 251200
rect 466656 244202 466684 251194
rect 466564 244174 466684 244202
rect 466564 241466 466592 244174
rect 466552 241460 466604 241466
rect 466552 241402 466604 241408
rect 466644 241460 466696 241466
rect 466644 241402 466696 241408
rect 466656 224890 466684 241402
rect 466564 224862 466684 224890
rect 466564 222154 466592 224862
rect 466552 222148 466604 222154
rect 466552 222090 466604 222096
rect 466644 222148 466696 222154
rect 466644 222090 466696 222096
rect 466656 205578 466684 222090
rect 466564 205550 466684 205578
rect 466564 196058 466592 205550
rect 466472 196030 466592 196058
rect 466472 195922 466500 196030
rect 466472 195894 466592 195922
rect 466564 186402 466592 195894
rect 466564 186374 466684 186402
rect 466656 167074 466684 186374
rect 466460 167068 466512 167074
rect 466460 167010 466512 167016
rect 466644 167068 466696 167074
rect 466644 167010 466696 167016
rect 466472 166954 466500 167010
rect 466472 166926 466592 166954
rect 466564 164218 466592 166926
rect 466552 164212 466604 164218
rect 466552 164154 466604 164160
rect 466552 157344 466604 157350
rect 466552 157286 466604 157292
rect 466564 154578 466592 157286
rect 466564 154550 466684 154578
rect 466656 147694 466684 154550
rect 466460 147688 466512 147694
rect 466644 147688 466696 147694
rect 466512 147636 466592 147642
rect 466460 147630 466592 147636
rect 466644 147630 466696 147636
rect 466472 147614 466592 147630
rect 466564 144906 466592 147614
rect 466552 144900 466604 144906
rect 466552 144842 466604 144848
rect 466552 137964 466604 137970
rect 466552 137906 466604 137912
rect 466564 135266 466592 137906
rect 466564 135238 466684 135266
rect 466656 124166 466684 135238
rect 466644 124160 466696 124166
rect 466644 124102 466696 124108
rect 466828 114572 466880 114578
rect 466828 114514 466880 114520
rect 466840 95266 466868 114514
rect 466552 95260 466604 95266
rect 466552 95202 466604 95208
rect 466828 95260 466880 95266
rect 466828 95202 466880 95208
rect 466564 89842 466592 95202
rect 466564 89814 466684 89842
rect 466656 87038 466684 89814
rect 466552 87032 466604 87038
rect 466472 86980 466552 86986
rect 466472 86974 466604 86980
rect 466644 87032 466696 87038
rect 466644 86974 466696 86980
rect 466472 86958 466592 86974
rect 466472 85542 466500 86958
rect 466460 85536 466512 85542
rect 466460 85478 466512 85484
rect 466552 77172 466604 77178
rect 466552 77114 466604 77120
rect 466564 60738 466592 77114
rect 466564 60710 466684 60738
rect 466656 57934 466684 60710
rect 466644 57928 466696 57934
rect 466644 57870 466696 57876
rect 466552 48340 466604 48346
rect 466552 48282 466604 48288
rect 466564 41426 466592 48282
rect 466564 41398 466684 41426
rect 466656 12458 466684 41398
rect 466656 12430 466776 12458
rect 465632 3528 465684 3534
rect 465632 3470 465684 3476
rect 466368 3528 466420 3534
rect 466368 3470 466420 3476
rect 464436 3324 464488 3330
rect 462044 2916 462096 2922
rect 462044 2858 462096 2864
rect 462056 480 462084 2858
rect 463252 480 463280 3318
rect 464436 3266 464488 3272
rect 464988 3324 465040 3330
rect 464988 3266 465040 3272
rect 464448 480 464476 3266
rect 465644 480 465672 3470
rect 466748 2922 466776 12430
rect 467760 3738 467788 336806
rect 469864 336796 469916 336802
rect 469864 336738 469916 336744
rect 469876 4146 469904 336738
rect 469128 4140 469180 4146
rect 469128 4082 469180 4088
rect 469864 4140 469916 4146
rect 469864 4082 469916 4088
rect 470324 4140 470376 4146
rect 470324 4082 470376 4088
rect 467932 3868 467984 3874
rect 467932 3810 467984 3816
rect 466828 3732 466880 3738
rect 466828 3674 466880 3680
rect 467748 3732 467800 3738
rect 467748 3674 467800 3680
rect 466736 2916 466788 2922
rect 466736 2858 466788 2864
rect 466840 480 466868 3674
rect 467944 480 467972 3810
rect 469140 480 469168 4082
rect 470336 480 470364 4082
rect 470704 3874 470732 340054
rect 471256 336802 471284 340068
rect 471348 340054 471822 340082
rect 471992 340054 472466 340082
rect 472544 340054 473110 340082
rect 473372 340054 473662 340082
rect 474306 340054 474688 340082
rect 471244 336796 471296 336802
rect 471244 336738 471296 336744
rect 471348 335730 471376 340054
rect 471992 336784 472020 340054
rect 470796 335702 471376 335730
rect 471900 336756 472020 336784
rect 470796 4146 470824 335702
rect 470784 4140 470836 4146
rect 470784 4082 470836 4088
rect 470692 3868 470744 3874
rect 470692 3810 470744 3816
rect 471900 2854 471928 336756
rect 472544 333282 472572 340054
rect 472176 333254 472572 333282
rect 472176 328438 472204 333254
rect 472164 328432 472216 328438
rect 472164 328374 472216 328380
rect 472072 318844 472124 318850
rect 472072 318786 472124 318792
rect 472084 311930 472112 318786
rect 471992 311902 472112 311930
rect 471992 311846 472020 311902
rect 471980 311840 472032 311846
rect 471980 311782 472032 311788
rect 472164 311840 472216 311846
rect 472164 311782 472216 311788
rect 472176 309126 472204 311782
rect 472164 309120 472216 309126
rect 472164 309062 472216 309068
rect 472072 299532 472124 299538
rect 472072 299474 472124 299480
rect 472084 292618 472112 299474
rect 471992 292590 472112 292618
rect 471992 292534 472020 292590
rect 471980 292528 472032 292534
rect 471980 292470 472032 292476
rect 472164 292528 472216 292534
rect 472164 292470 472216 292476
rect 472176 280242 472204 292470
rect 472084 280214 472204 280242
rect 472084 280158 472112 280214
rect 472072 280152 472124 280158
rect 472072 280094 472124 280100
rect 472164 270564 472216 270570
rect 472164 270506 472216 270512
rect 472176 263514 472204 270506
rect 472084 263486 472204 263514
rect 472084 260846 472112 263486
rect 472072 260840 472124 260846
rect 472072 260782 472124 260788
rect 472164 251252 472216 251258
rect 472164 251194 472216 251200
rect 472176 244202 472204 251194
rect 472084 244174 472204 244202
rect 472084 241505 472112 244174
rect 472070 241496 472126 241505
rect 472070 241431 472126 241440
rect 472346 241496 472402 241505
rect 472346 241431 472402 241440
rect 472360 231878 472388 241431
rect 472164 231872 472216 231878
rect 472164 231814 472216 231820
rect 472348 231872 472400 231878
rect 472348 231814 472400 231820
rect 472176 224890 472204 231814
rect 472084 224862 472204 224890
rect 472084 222193 472112 224862
rect 472070 222184 472126 222193
rect 472070 222119 472126 222128
rect 472346 222184 472402 222193
rect 472346 222119 472402 222128
rect 472360 212566 472388 222119
rect 472164 212560 472216 212566
rect 472164 212502 472216 212508
rect 472348 212560 472400 212566
rect 472348 212502 472400 212508
rect 472176 205578 472204 212502
rect 472084 205550 472204 205578
rect 472084 202881 472112 205550
rect 472070 202872 472126 202881
rect 472070 202807 472126 202816
rect 472346 202872 472402 202881
rect 472346 202807 472402 202816
rect 472360 193254 472388 202807
rect 472164 193248 472216 193254
rect 472164 193190 472216 193196
rect 472348 193248 472400 193254
rect 472348 193190 472400 193196
rect 472176 186266 472204 193190
rect 472084 186238 472204 186266
rect 472084 183569 472112 186238
rect 472070 183560 472126 183569
rect 472070 183495 472126 183504
rect 472346 183560 472402 183569
rect 472346 183495 472402 183504
rect 472360 173942 472388 183495
rect 472164 173936 472216 173942
rect 472164 173878 472216 173884
rect 472348 173936 472400 173942
rect 472348 173878 472400 173884
rect 472176 166954 472204 173878
rect 472084 166926 472204 166954
rect 472084 164218 472112 166926
rect 472072 164212 472124 164218
rect 472072 164154 472124 164160
rect 472348 164212 472400 164218
rect 472348 164154 472400 164160
rect 472360 154601 472388 164154
rect 472162 154592 472218 154601
rect 472162 154527 472218 154536
rect 472346 154592 472402 154601
rect 472346 154527 472402 154536
rect 472176 147642 472204 154527
rect 472084 147614 472204 147642
rect 472084 138038 472112 147614
rect 472072 138032 472124 138038
rect 472072 137974 472124 137980
rect 471980 137964 472032 137970
rect 471980 137906 472032 137912
rect 471992 135289 472020 137906
rect 471978 135280 472034 135289
rect 471978 135215 472034 135224
rect 472162 135280 472218 135289
rect 472162 135215 472218 135224
rect 472176 128330 472204 135215
rect 472084 128302 472204 128330
rect 472084 118726 472112 128302
rect 472072 118720 472124 118726
rect 472072 118662 472124 118668
rect 471980 118652 472032 118658
rect 471980 118594 472032 118600
rect 471992 115977 472020 118594
rect 471978 115968 472034 115977
rect 471978 115903 472034 115912
rect 472162 115968 472218 115977
rect 472162 115903 472218 115912
rect 472176 109018 472204 115903
rect 472084 108990 472204 109018
rect 472084 99414 472112 108990
rect 472072 99408 472124 99414
rect 472072 99350 472124 99356
rect 471980 99340 472032 99346
rect 471980 99282 472032 99288
rect 471992 96665 472020 99282
rect 471978 96656 472034 96665
rect 471978 96591 472034 96600
rect 472162 96656 472218 96665
rect 472162 96591 472218 96600
rect 472176 89706 472204 96591
rect 472084 89678 472204 89706
rect 472084 85542 472112 89678
rect 472072 85536 472124 85542
rect 472072 85478 472124 85484
rect 472072 67652 472124 67658
rect 472072 67594 472124 67600
rect 472084 60738 472112 67594
rect 471992 60722 472112 60738
rect 471980 60716 472112 60722
rect 472032 60710 472112 60716
rect 472164 60716 472216 60722
rect 471980 60658 472032 60664
rect 472164 60658 472216 60664
rect 472176 57934 472204 60658
rect 472164 57928 472216 57934
rect 472164 57870 472216 57876
rect 472072 48340 472124 48346
rect 472072 48282 472124 48288
rect 472084 41426 472112 48282
rect 471992 41410 472112 41426
rect 471980 41404 472112 41410
rect 472032 41398 472112 41404
rect 472164 41404 472216 41410
rect 471980 41346 472032 41352
rect 472164 41346 472216 41352
rect 472176 38622 472204 41346
rect 472164 38616 472216 38622
rect 472164 38558 472216 38564
rect 472164 31204 472216 31210
rect 472164 31146 472216 31152
rect 472176 22302 472204 31146
rect 473266 29336 473322 29345
rect 473266 29271 473322 29280
rect 473280 29238 473308 29271
rect 473268 29232 473320 29238
rect 473268 29174 473320 29180
rect 472164 22296 472216 22302
rect 472164 22238 472216 22244
rect 472164 19372 472216 19378
rect 472164 19314 472216 19320
rect 472176 4146 472204 19314
rect 473372 4146 473400 340054
rect 474660 4146 474688 340054
rect 474936 336802 474964 340068
rect 475488 337686 475516 340068
rect 475476 337680 475528 337686
rect 475476 337622 475528 337628
rect 476132 336802 476160 340068
rect 476776 336938 476804 340068
rect 476764 336932 476816 336938
rect 476764 336874 476816 336880
rect 474924 336796 474976 336802
rect 474924 336738 474976 336744
rect 476028 336796 476080 336802
rect 476028 336738 476080 336744
rect 476120 336796 476172 336802
rect 476120 336738 476172 336744
rect 475934 180976 475990 180985
rect 475934 180911 475936 180920
rect 475988 180911 475990 180920
rect 475936 180882 475988 180888
rect 475934 169960 475990 169969
rect 475934 169895 475936 169904
rect 475988 169895 475990 169904
rect 475936 169866 475988 169872
rect 475934 123040 475990 123049
rect 475934 122975 475936 122984
rect 475988 122975 475990 122984
rect 475936 122946 475988 122952
rect 475934 87136 475990 87145
rect 475934 87071 475936 87080
rect 475988 87071 475990 87080
rect 475936 87042 475988 87048
rect 475934 76120 475990 76129
rect 475934 76055 475936 76064
rect 475988 76055 475990 76064
rect 475936 76026 475988 76032
rect 472164 4140 472216 4146
rect 472164 4082 472216 4088
rect 472716 4140 472768 4146
rect 472716 4082 472768 4088
rect 473360 4140 473412 4146
rect 473360 4082 473412 4088
rect 473912 4140 473964 4146
rect 473912 4082 473964 4088
rect 474648 4140 474700 4146
rect 474648 4082 474700 4088
rect 475108 4140 475160 4146
rect 475108 4082 475160 4088
rect 471520 2848 471572 2854
rect 471520 2790 471572 2796
rect 471888 2848 471940 2854
rect 471888 2790 471940 2796
rect 471532 480 471560 2790
rect 472728 480 472756 4082
rect 473924 480 473952 4082
rect 475120 480 475148 4082
rect 476040 3618 476068 336738
rect 477328 327146 477356 340068
rect 477684 337680 477736 337686
rect 477684 337622 477736 337628
rect 477408 336932 477460 336938
rect 477408 336874 477460 336880
rect 477316 327140 477368 327146
rect 477316 327082 477368 327088
rect 476118 180976 476174 180985
rect 476118 180911 476120 180920
rect 476172 180911 476174 180920
rect 476120 180882 476172 180888
rect 476118 169960 476174 169969
rect 476118 169895 476120 169904
rect 476172 169895 476174 169904
rect 476120 169866 476172 169872
rect 476118 87136 476174 87145
rect 476118 87071 476120 87080
rect 476172 87071 476174 87080
rect 476120 87042 476172 87048
rect 477420 4078 477448 336874
rect 477592 336796 477644 336802
rect 477592 336738 477644 336744
rect 477604 7614 477632 336738
rect 477592 7608 477644 7614
rect 477592 7550 477644 7556
rect 477696 7426 477724 337622
rect 477972 336802 478000 340068
rect 478524 336938 478552 340068
rect 479168 337006 479196 340068
rect 479812 337550 479840 340068
rect 479800 337544 479852 337550
rect 479800 337486 479852 337492
rect 479156 337000 479208 337006
rect 479156 336942 479208 336948
rect 478512 336932 478564 336938
rect 478512 336874 478564 336880
rect 480364 336802 480392 340068
rect 481008 336870 481036 340068
rect 480996 336864 481048 336870
rect 480996 336806 481048 336812
rect 481652 336802 481680 340068
rect 482204 337074 482232 340068
rect 482848 337414 482876 340068
rect 482836 337408 482888 337414
rect 482836 337350 482888 337356
rect 482192 337068 482244 337074
rect 482192 337010 482244 337016
rect 482836 337068 482888 337074
rect 482836 337010 482888 337016
rect 477960 336796 478012 336802
rect 477960 336738 478012 336744
rect 478788 336796 478840 336802
rect 478788 336738 478840 336744
rect 480352 336796 480404 336802
rect 480352 336738 480404 336744
rect 481548 336796 481600 336802
rect 481548 336738 481600 336744
rect 481640 336796 481692 336802
rect 481640 336738 481692 336744
rect 478142 123040 478198 123049
rect 478142 122975 478144 122984
rect 478196 122975 478198 122984
rect 478144 122946 478196 122952
rect 478142 76120 478198 76129
rect 478142 76055 478144 76064
rect 478196 76055 478198 76064
rect 478144 76026 478196 76032
rect 478696 7608 478748 7614
rect 478696 7550 478748 7556
rect 477512 7398 477724 7426
rect 477408 4072 477460 4078
rect 477408 4014 477460 4020
rect 476040 3590 476344 3618
rect 476316 480 476344 3590
rect 477512 480 477540 7398
rect 478708 480 478736 7550
rect 478800 4146 478828 336738
rect 480352 327140 480404 327146
rect 480352 327082 480404 327088
rect 480364 317422 480392 327082
rect 480352 317416 480404 317422
rect 480352 317358 480404 317364
rect 480352 307828 480404 307834
rect 480352 307770 480404 307776
rect 480364 298110 480392 307770
rect 480352 298104 480404 298110
rect 480352 298046 480404 298052
rect 480352 288448 480404 288454
rect 480352 288390 480404 288396
rect 480364 278769 480392 288390
rect 480166 278760 480222 278769
rect 480166 278695 480222 278704
rect 480350 278760 480406 278769
rect 480350 278695 480406 278704
rect 480180 269142 480208 278695
rect 480168 269136 480220 269142
rect 480168 269078 480220 269084
rect 480352 269136 480404 269142
rect 480352 269078 480404 269084
rect 480364 259457 480392 269078
rect 480166 259448 480222 259457
rect 480166 259383 480222 259392
rect 480350 259448 480406 259457
rect 480350 259383 480406 259392
rect 480180 249830 480208 259383
rect 480168 249824 480220 249830
rect 480168 249766 480220 249772
rect 480352 249824 480404 249830
rect 480352 249766 480404 249772
rect 480364 241777 480392 249766
rect 480350 241768 480406 241777
rect 480350 241703 480406 241712
rect 480350 241632 480406 241641
rect 480350 241567 480406 241576
rect 480364 240145 480392 241567
rect 480166 240136 480222 240145
rect 480166 240071 480222 240080
rect 480350 240136 480406 240145
rect 480350 240071 480406 240080
rect 480180 230518 480208 240071
rect 480168 230512 480220 230518
rect 480168 230454 480220 230460
rect 480352 230512 480404 230518
rect 480352 230454 480404 230460
rect 480364 220833 480392 230454
rect 480166 220824 480222 220833
rect 480166 220759 480222 220768
rect 480350 220824 480406 220833
rect 480350 220759 480406 220768
rect 480180 211177 480208 220759
rect 480166 211168 480222 211177
rect 480166 211103 480222 211112
rect 480350 211168 480406 211177
rect 480350 211103 480406 211112
rect 480364 202978 480392 211103
rect 480352 202972 480404 202978
rect 480352 202914 480404 202920
rect 480260 201544 480312 201550
rect 480260 201486 480312 201492
rect 480272 196042 480300 201486
rect 480260 196036 480312 196042
rect 480260 195978 480312 195984
rect 480352 195900 480404 195906
rect 480352 195842 480404 195848
rect 480364 186266 480392 195842
rect 480364 186238 480484 186266
rect 480456 183546 480484 186238
rect 480364 183518 480484 183546
rect 480364 178838 480392 183518
rect 480352 178832 480404 178838
rect 480352 178774 480404 178780
rect 480352 178696 480404 178702
rect 480352 178638 480404 178644
rect 480364 169114 480392 178638
rect 480352 169108 480404 169114
rect 480352 169050 480404 169056
rect 480536 169108 480588 169114
rect 480536 169050 480588 169056
rect 480548 164257 480576 169050
rect 480350 164248 480406 164257
rect 480350 164183 480352 164192
rect 480404 164183 480406 164192
rect 480534 164248 480590 164257
rect 480534 164183 480590 164192
rect 480352 164154 480404 164160
rect 480260 153264 480312 153270
rect 480260 153206 480312 153212
rect 480272 143546 480300 153206
rect 480260 143540 480312 143546
rect 480260 143482 480312 143488
rect 480444 143540 480496 143546
rect 480444 143482 480496 143488
rect 480456 115977 480484 143482
rect 480258 115968 480314 115977
rect 480258 115903 480314 115912
rect 480442 115968 480498 115977
rect 480442 115903 480498 115912
rect 480272 111058 480300 115903
rect 480272 111030 480484 111058
rect 480456 104854 480484 111030
rect 480444 104848 480496 104854
rect 480444 104790 480496 104796
rect 480536 95260 480588 95266
rect 480536 95202 480588 95208
rect 480548 89706 480576 95202
rect 480456 89678 480576 89706
rect 480456 85542 480484 89678
rect 480444 85536 480496 85542
rect 480444 85478 480496 85484
rect 480536 77172 480588 77178
rect 480536 77114 480588 77120
rect 480548 67674 480576 77114
rect 480456 67646 480576 67674
rect 480456 67590 480484 67646
rect 480260 67584 480312 67590
rect 480260 67526 480312 67532
rect 480444 67584 480496 67590
rect 480444 67526 480496 67532
rect 480272 58018 480300 67526
rect 480272 57990 480392 58018
rect 480364 57934 480392 57990
rect 480352 57928 480404 57934
rect 480352 57870 480404 57876
rect 480536 57928 480588 57934
rect 480536 57870 480588 57876
rect 480548 38758 480576 57870
rect 480260 38752 480312 38758
rect 480260 38694 480312 38700
rect 480536 38752 480588 38758
rect 480536 38694 480588 38700
rect 480272 31822 480300 38694
rect 480260 31816 480312 31822
rect 480260 31758 480312 31764
rect 480352 31680 480404 31686
rect 480352 31622 480404 31628
rect 480364 27606 480392 31622
rect 480352 27600 480404 27606
rect 480352 27542 480404 27548
rect 480352 18012 480404 18018
rect 480352 17954 480404 17960
rect 478788 4140 478840 4146
rect 478788 4082 478840 4088
rect 479892 4072 479944 4078
rect 479892 4014 479944 4020
rect 479904 480 479932 4014
rect 480364 1018 480392 17954
rect 481560 3330 481588 336738
rect 482284 4140 482336 4146
rect 482284 4082 482336 4088
rect 481548 3324 481600 3330
rect 481548 3266 481600 3272
rect 480352 1012 480404 1018
rect 480352 954 480404 960
rect 481088 1012 481140 1018
rect 481088 954 481140 960
rect 481100 480 481128 954
rect 482296 480 482324 4082
rect 482848 3874 482876 337010
rect 483204 336932 483256 336938
rect 483204 336874 483256 336880
rect 482928 336796 482980 336802
rect 482928 336738 482980 336744
rect 482836 3868 482888 3874
rect 482836 3810 482888 3816
rect 482940 3398 482968 336738
rect 482928 3392 482980 3398
rect 482928 3334 482980 3340
rect 483216 626 483244 336874
rect 483492 336802 483520 340068
rect 484058 340054 484256 340082
rect 483480 336796 483532 336802
rect 483480 336738 483532 336744
rect 484228 3602 484256 340054
rect 484584 337000 484636 337006
rect 484584 336942 484636 336948
rect 484308 336796 484360 336802
rect 484308 336738 484360 336744
rect 484320 3670 484348 336738
rect 484308 3664 484360 3670
rect 484308 3606 484360 3612
rect 484216 3596 484268 3602
rect 484216 3538 484268 3544
rect 483216 598 483520 626
rect 483492 480 483520 598
rect 484596 480 484624 336942
rect 484688 336802 484716 340068
rect 485332 337482 485360 340068
rect 485884 337686 485912 340068
rect 486542 340054 487108 340082
rect 485872 337680 485924 337686
rect 485872 337622 485924 337628
rect 485964 337544 486016 337550
rect 485964 337486 486016 337492
rect 485320 337476 485372 337482
rect 485320 337418 485372 337424
rect 485044 336864 485096 336870
rect 485044 336806 485096 336812
rect 484676 336796 484728 336802
rect 484676 336738 484728 336744
rect 485056 3262 485084 336806
rect 485688 336796 485740 336802
rect 485688 336738 485740 336744
rect 485700 3738 485728 336738
rect 485688 3732 485740 3738
rect 485688 3674 485740 3680
rect 485044 3256 485096 3262
rect 485044 3198 485096 3204
rect 485976 626 486004 337486
rect 487080 3534 487108 340054
rect 487172 337754 487200 340068
rect 488276 337770 488304 340190
rect 488382 340054 488488 340082
rect 487160 337748 487212 337754
rect 488276 337742 488396 337770
rect 487160 337690 487212 337696
rect 487068 3528 487120 3534
rect 487068 3470 487120 3476
rect 488368 3466 488396 337742
rect 488356 3460 488408 3466
rect 488356 3402 488408 3408
rect 488460 3330 488488 340054
rect 489012 337822 489040 340068
rect 489578 340054 489868 340082
rect 489000 337816 489052 337822
rect 489000 337758 489052 337764
rect 489184 337680 489236 337686
rect 489184 337622 489236 337628
rect 489196 3806 489224 337622
rect 489184 3800 489236 3806
rect 489184 3742 489236 3748
rect 489368 3392 489420 3398
rect 489368 3334 489420 3340
rect 486976 3324 487028 3330
rect 486976 3266 487028 3272
rect 488448 3324 488500 3330
rect 488448 3266 488500 3272
rect 485792 598 486004 626
rect 485792 480 485820 598
rect 486988 480 487016 3266
rect 488172 3256 488224 3262
rect 488172 3198 488224 3204
rect 488184 480 488212 3198
rect 489380 480 489408 3334
rect 489840 3262 489868 340054
rect 490208 337958 490236 340068
rect 490852 338026 490880 340068
rect 490840 338020 490892 338026
rect 490840 337962 490892 337968
rect 490196 337952 490248 337958
rect 490196 337894 490248 337900
rect 491404 337686 491432 340068
rect 492062 340054 492628 340082
rect 491392 337680 491444 337686
rect 491392 337622 491444 337628
rect 492496 337680 492548 337686
rect 492496 337622 492548 337628
rect 491484 337408 491536 337414
rect 491484 337350 491536 337356
rect 490564 3868 490616 3874
rect 490564 3810 490616 3816
rect 489828 3256 489880 3262
rect 489828 3198 489880 3204
rect 490576 480 490604 3810
rect 491496 626 491524 337350
rect 492508 3398 492536 337622
rect 492600 4078 492628 340054
rect 492692 337618 492720 340068
rect 493796 337736 493824 340190
rect 493902 340054 494008 340082
rect 493796 337708 493916 337736
rect 492680 337612 492732 337618
rect 492680 337554 492732 337560
rect 493324 337476 493376 337482
rect 493324 337418 493376 337424
rect 492588 4072 492640 4078
rect 492588 4014 492640 4020
rect 492956 3664 493008 3670
rect 492956 3606 493008 3612
rect 492496 3392 492548 3398
rect 492496 3334 492548 3340
rect 491496 598 491708 626
rect 491680 592 491708 598
rect 491680 564 491800 592
rect 491772 480 491800 564
rect 492968 480 492996 3606
rect 493336 3194 493364 337418
rect 493888 4010 493916 337708
rect 493980 4146 494008 340054
rect 494532 337550 494560 340068
rect 495084 337686 495112 340068
rect 495072 337680 495124 337686
rect 495072 337622 495124 337628
rect 494520 337544 494572 337550
rect 494520 337486 494572 337492
rect 495728 337278 495756 340068
rect 496084 337680 496136 337686
rect 496084 337622 496136 337628
rect 495716 337272 495768 337278
rect 495716 337214 495768 337220
rect 493968 4140 494020 4146
rect 493968 4082 494020 4088
rect 493876 4004 493928 4010
rect 493876 3946 493928 3952
rect 496096 3942 496124 337622
rect 496280 337482 496308 340068
rect 496924 337686 496952 340068
rect 497568 337890 497596 340068
rect 497556 337884 497608 337890
rect 497556 337826 497608 337832
rect 496912 337680 496964 337686
rect 496912 337622 496964 337628
rect 496268 337476 496320 337482
rect 496268 337418 496320 337424
rect 496728 337272 496780 337278
rect 496728 337214 496780 337220
rect 496084 3936 496136 3942
rect 496084 3878 496136 3884
rect 496740 3874 496768 337214
rect 498120 337210 498148 340068
rect 498108 337204 498160 337210
rect 498108 337146 498160 337152
rect 498764 336938 498792 340068
rect 498844 337680 498896 337686
rect 498844 337622 498896 337628
rect 498752 336932 498804 336938
rect 498752 336874 498804 336880
rect 496728 3868 496780 3874
rect 496728 3810 496780 3816
rect 497740 3800 497792 3806
rect 497740 3742 497792 3748
rect 495348 3732 495400 3738
rect 495348 3674 495400 3680
rect 494152 3596 494204 3602
rect 494152 3538 494204 3544
rect 493324 3188 493376 3194
rect 493324 3130 493376 3136
rect 494164 480 494192 3538
rect 495360 480 495388 3674
rect 496544 3188 496596 3194
rect 496544 3130 496596 3136
rect 496556 480 496584 3130
rect 497752 480 497780 3742
rect 498856 3738 498884 337622
rect 498844 3732 498896 3738
rect 498844 3674 498896 3680
rect 499408 3602 499436 340068
rect 499960 337754 499988 340068
rect 500618 340054 500816 340082
rect 499764 337748 499816 337754
rect 499764 337690 499816 337696
rect 499948 337748 500000 337754
rect 499948 337690 500000 337696
rect 499488 336932 499540 336938
rect 499488 336874 499540 336880
rect 499500 3670 499528 336874
rect 499488 3664 499540 3670
rect 499488 3606 499540 3612
rect 499396 3596 499448 3602
rect 499396 3538 499448 3544
rect 498936 3528 498988 3534
rect 498936 3470 498988 3476
rect 498948 480 498976 3470
rect 499776 610 499804 337690
rect 500788 3534 500816 340054
rect 501248 337754 501276 340068
rect 501814 340054 502288 340082
rect 501604 337952 501656 337958
rect 501604 337894 501656 337900
rect 500868 337748 500920 337754
rect 500868 337690 500920 337696
rect 501236 337748 501288 337754
rect 501236 337690 501288 337696
rect 500880 3806 500908 337690
rect 500868 3800 500920 3806
rect 500868 3742 500920 3748
rect 500776 3528 500828 3534
rect 500776 3470 500828 3476
rect 501236 3460 501288 3466
rect 501236 3402 501288 3408
rect 499764 604 499816 610
rect 499764 546 499816 552
rect 500132 604 500184 610
rect 500132 546 500184 552
rect 500144 480 500172 546
rect 501248 480 501276 3402
rect 501616 3126 501644 337894
rect 502260 3466 502288 340054
rect 502444 337618 502472 340068
rect 503102 340054 503576 340082
rect 503444 337952 503496 337958
rect 503444 337894 503496 337900
rect 502616 337816 502668 337822
rect 502616 337758 502668 337764
rect 502432 337612 502484 337618
rect 502432 337554 502484 337560
rect 502248 3460 502300 3466
rect 502248 3402 502300 3408
rect 502628 3346 502656 337758
rect 503456 336802 503484 337894
rect 503548 337770 503576 340054
rect 503640 337958 503668 340068
rect 503628 337952 503680 337958
rect 503628 337894 503680 337900
rect 504284 337822 504312 340068
rect 504272 337816 504324 337822
rect 503548 337742 503668 337770
rect 504272 337758 504324 337764
rect 503536 337612 503588 337618
rect 503536 337554 503588 337560
rect 503444 336796 503496 336802
rect 503444 336738 503496 336744
rect 503548 4962 503576 337554
rect 503536 4956 503588 4962
rect 503536 4898 503588 4904
rect 503640 3584 503668 337742
rect 504928 336938 504956 340068
rect 505008 337816 505060 337822
rect 505008 337758 505060 337764
rect 504916 336932 504968 336938
rect 504916 336874 504968 336880
rect 503640 3556 503760 3584
rect 502432 3324 502484 3330
rect 502628 3318 503668 3346
rect 502432 3266 502484 3272
rect 501604 3120 501656 3126
rect 501604 3062 501656 3068
rect 502444 480 502472 3266
rect 503640 480 503668 3318
rect 503732 2922 503760 3556
rect 504824 3256 504876 3262
rect 504824 3198 504876 3204
rect 503720 2916 503772 2922
rect 503720 2858 503772 2864
rect 504836 480 504864 3198
rect 505020 2990 505048 337758
rect 505480 337754 505508 340068
rect 506138 340054 506336 340082
rect 505468 337748 505520 337754
rect 505468 337690 505520 337696
rect 506308 4826 506336 340054
rect 506388 337748 506440 337754
rect 506388 337690 506440 337696
rect 506296 4820 506348 4826
rect 506296 4762 506348 4768
rect 506020 3120 506072 3126
rect 506020 3062 506072 3068
rect 505008 2984 505060 2990
rect 505008 2926 505060 2932
rect 506032 480 506060 3062
rect 506400 3058 506428 337690
rect 506664 337340 506716 337346
rect 506664 337282 506716 337288
rect 506388 3052 506440 3058
rect 506388 2994 506440 3000
rect 506676 610 506704 337282
rect 506768 337278 506796 340068
rect 506756 337272 506808 337278
rect 506756 337214 506808 337220
rect 507320 337142 507348 340068
rect 507964 337822 507992 340068
rect 507952 337816 508004 337822
rect 507952 337758 508004 337764
rect 508608 337618 508636 340068
rect 509068 340054 509174 340082
rect 508596 337612 508648 337618
rect 508596 337554 508648 337560
rect 507768 337272 507820 337278
rect 507768 337214 507820 337220
rect 507308 337136 507360 337142
rect 507308 337078 507360 337084
rect 507780 3126 507808 337214
rect 509068 337210 509096 340054
rect 509148 337816 509200 337822
rect 509148 337758 509200 337764
rect 509056 337204 509108 337210
rect 509056 337146 509108 337152
rect 509160 4894 509188 337758
rect 509804 337074 509832 340068
rect 510462 340054 510568 340082
rect 509884 337884 509936 337890
rect 509884 337826 509936 337832
rect 509792 337068 509844 337074
rect 509792 337010 509844 337016
rect 509148 4888 509200 4894
rect 509148 4830 509200 4836
rect 509608 4072 509660 4078
rect 509608 4014 509660 4020
rect 508412 3392 508464 3398
rect 508412 3334 508464 3340
rect 507768 3120 507820 3126
rect 507768 3062 507820 3068
rect 506664 604 506716 610
rect 506664 546 506716 552
rect 507216 604 507268 610
rect 507216 546 507268 552
rect 507228 480 507256 546
rect 508424 480 508452 3334
rect 509620 480 509648 4014
rect 509896 3874 509924 337826
rect 510540 4078 510568 340054
rect 510804 337680 510856 337686
rect 510804 337622 510856 337628
rect 510528 4072 510580 4078
rect 510528 4014 510580 4020
rect 509884 3868 509936 3874
rect 509884 3810 509936 3816
rect 510816 480 510844 337622
rect 511000 337482 511028 340068
rect 511658 340054 511948 340082
rect 510988 337476 511040 337482
rect 510988 337418 511040 337424
rect 511816 337476 511868 337482
rect 511816 337418 511868 337424
rect 511828 3262 511856 337418
rect 511816 3256 511868 3262
rect 511816 3198 511868 3204
rect 511920 3194 511948 340054
rect 512288 338094 512316 340068
rect 512276 338088 512328 338094
rect 512276 338030 512328 338036
rect 512840 338026 512868 340068
rect 512828 338020 512880 338026
rect 512828 337962 512880 337968
rect 513484 336870 513512 340068
rect 514588 337668 514616 340190
rect 514680 337890 514708 340068
rect 514668 337884 514720 337890
rect 514668 337826 514720 337832
rect 514588 337640 514708 337668
rect 513564 337544 513616 337550
rect 513564 337486 513616 337492
rect 513472 336864 513524 336870
rect 513472 336806 513524 336812
rect 513196 4140 513248 4146
rect 513196 4082 513248 4088
rect 512000 4004 512052 4010
rect 512000 3946 512052 3952
rect 511908 3188 511960 3194
rect 511908 3130 511960 3136
rect 512012 480 512040 3946
rect 513208 480 513236 4082
rect 513576 610 513604 337486
rect 514574 204504 514630 204513
rect 514574 204439 514630 204448
rect 514588 204105 514616 204439
rect 514574 204096 514630 204105
rect 514574 204031 514630 204040
rect 514574 180976 514630 180985
rect 514574 180911 514630 180920
rect 514588 180577 514616 180911
rect 514574 180568 514630 180577
rect 514574 180503 514630 180512
rect 514576 169992 514628 169998
rect 514574 169960 514576 169969
rect 514628 169960 514630 169969
rect 514574 169895 514630 169904
rect 514574 157584 514630 157593
rect 514574 157519 514630 157528
rect 514588 157185 514616 157519
rect 514574 157176 514630 157185
rect 514574 157111 514630 157120
rect 514574 134056 514630 134065
rect 514574 133991 514630 134000
rect 514588 133657 514616 133991
rect 514574 133648 514630 133657
rect 514574 133583 514630 133592
rect 514576 123072 514628 123078
rect 514574 123040 514576 123049
rect 514628 123040 514630 123049
rect 514574 122975 514630 122984
rect 514574 110664 514630 110673
rect 514574 110599 514630 110608
rect 514588 110265 514616 110599
rect 514574 110256 514630 110265
rect 514574 110191 514630 110200
rect 514576 76152 514628 76158
rect 514574 76120 514576 76129
rect 514628 76120 514630 76129
rect 514574 76055 514630 76064
rect 514574 63744 514630 63753
rect 514574 63679 514630 63688
rect 514588 63345 514616 63679
rect 514574 63336 514630 63345
rect 514574 63271 514630 63280
rect 514574 40216 514630 40225
rect 514574 40151 514630 40160
rect 514588 39817 514616 40151
rect 514574 39808 514630 39817
rect 514574 39743 514630 39752
rect 514574 16824 514630 16833
rect 514574 16759 514576 16768
rect 514628 16759 514630 16768
rect 514576 16730 514628 16736
rect 514680 3398 514708 337640
rect 515324 337482 515352 340068
rect 515876 337822 515904 340068
rect 515864 337816 515916 337822
rect 515864 337758 515916 337764
rect 515312 337476 515364 337482
rect 515312 337418 515364 337424
rect 516520 337006 516548 340068
rect 516784 337680 516836 337686
rect 516784 337622 516836 337628
rect 516508 337000 516560 337006
rect 516508 336942 516560 336948
rect 516046 16824 516102 16833
rect 516046 16759 516048 16768
rect 516100 16759 516102 16768
rect 516048 16730 516100 16736
rect 516796 4876 516824 337622
rect 517164 337278 517192 340068
rect 517612 337408 517664 337414
rect 517612 337350 517664 337356
rect 517152 337272 517204 337278
rect 517152 337214 517204 337220
rect 517428 337000 517480 337006
rect 517428 336942 517480 336948
rect 516876 169992 516928 169998
rect 516874 169960 516876 169969
rect 516928 169960 516930 169969
rect 516874 169895 516930 169904
rect 516876 123072 516928 123078
rect 516874 123040 516876 123049
rect 516928 123040 516930 123049
rect 516874 122975 516930 122984
rect 516876 76152 516928 76158
rect 516874 76120 516876 76129
rect 516928 76120 516930 76129
rect 516874 76055 516930 76064
rect 516704 4848 516824 4876
rect 515588 3936 515640 3942
rect 515588 3878 515640 3884
rect 514668 3392 514720 3398
rect 514668 3334 514720 3340
rect 513564 604 513616 610
rect 513564 546 513616 552
rect 514392 604 514444 610
rect 514392 546 514444 552
rect 514404 480 514432 546
rect 515600 480 515628 3878
rect 516704 2854 516732 4848
rect 517440 4146 517468 336942
rect 517428 4140 517480 4146
rect 517428 4082 517480 4088
rect 516784 3324 516836 3330
rect 516784 3266 516836 3272
rect 516692 2848 516744 2854
rect 516692 2790 516744 2796
rect 516796 480 516824 3266
rect 517624 626 517652 337350
rect 517716 337006 517744 340068
rect 518360 337754 518388 340068
rect 518348 337748 518400 337754
rect 518348 337690 518400 337696
rect 519004 337006 519032 340068
rect 519556 337482 519584 340068
rect 519544 337476 519596 337482
rect 519544 337418 519596 337424
rect 517704 337000 517756 337006
rect 517704 336942 517756 336948
rect 518808 337000 518860 337006
rect 518808 336942 518860 336948
rect 518992 337000 519044 337006
rect 518992 336942 519044 336948
rect 520096 337000 520148 337006
rect 520096 336942 520148 336948
rect 518820 4078 518848 336942
rect 518808 4072 518860 4078
rect 518808 4014 518860 4020
rect 520108 4010 520136 336942
rect 520096 4004 520148 4010
rect 520096 3946 520148 3952
rect 520200 3942 520228 340068
rect 520844 337958 520872 340068
rect 521410 340054 521608 340082
rect 520832 337952 520884 337958
rect 520832 337894 520884 337900
rect 520372 337340 520424 337346
rect 520372 337282 520424 337288
rect 520188 3936 520240 3942
rect 520188 3878 520240 3884
rect 520280 3868 520332 3874
rect 520280 3810 520332 3816
rect 519084 3732 519136 3738
rect 519084 3674 519136 3680
rect 517624 598 517928 626
rect 517900 480 517928 598
rect 519096 480 519124 3674
rect 520292 480 520320 3810
rect 520384 610 520412 337282
rect 521580 3874 521608 340054
rect 522040 337278 522068 340068
rect 522698 340054 522988 340082
rect 522028 337272 522080 337278
rect 522028 337214 522080 337220
rect 521660 204400 521712 204406
rect 521658 204368 521660 204377
rect 521712 204368 521714 204377
rect 521658 204303 521714 204312
rect 521660 180872 521712 180878
rect 521658 180840 521660 180849
rect 521712 180840 521714 180849
rect 521658 180775 521714 180784
rect 521660 157480 521712 157486
rect 521658 157448 521660 157457
rect 521712 157448 521714 157457
rect 521658 157383 521714 157392
rect 521660 133952 521712 133958
rect 521658 133920 521660 133929
rect 521712 133920 521714 133929
rect 521658 133855 521714 133864
rect 521660 110560 521712 110566
rect 521658 110528 521660 110537
rect 521712 110528 521714 110537
rect 521658 110463 521714 110472
rect 521660 63640 521712 63646
rect 521658 63608 521660 63617
rect 521712 63608 521714 63617
rect 521658 63543 521714 63552
rect 521660 40112 521712 40118
rect 521658 40080 521660 40089
rect 521712 40080 521714 40089
rect 521658 40015 521714 40024
rect 521660 29096 521712 29102
rect 521658 29064 521660 29073
rect 521712 29064 521714 29073
rect 521658 28999 521714 29008
rect 521568 3868 521620 3874
rect 521568 3810 521620 3816
rect 522960 3738 522988 340054
rect 523236 337793 523264 340068
rect 523894 340054 524368 340082
rect 523222 337784 523278 337793
rect 523222 337719 523278 337728
rect 524236 169856 524288 169862
rect 524234 169824 524236 169833
rect 524288 169824 524290 169833
rect 524234 169759 524290 169768
rect 524236 122936 524288 122942
rect 524234 122904 524236 122913
rect 524288 122904 524290 122913
rect 524234 122839 524290 122848
rect 524236 76016 524288 76022
rect 524234 75984 524236 75993
rect 524288 75984 524290 75993
rect 524234 75919 524290 75928
rect 524236 16720 524288 16726
rect 524234 16688 524236 16697
rect 524288 16688 524290 16697
rect 524234 16623 524290 16632
rect 522948 3732 523000 3738
rect 522948 3674 523000 3680
rect 524340 3670 524368 340054
rect 524524 336802 524552 340068
rect 525090 340054 525564 340082
rect 524512 336796 524564 336802
rect 524512 336738 524564 336744
rect 525062 87000 525118 87009
rect 525062 86935 525118 86944
rect 525076 86737 525104 86935
rect 525062 86728 525118 86737
rect 525062 86663 525118 86672
rect 525064 3800 525116 3806
rect 525064 3742 525116 3748
rect 522672 3664 522724 3670
rect 522672 3606 522724 3612
rect 524328 3664 524380 3670
rect 524328 3606 524380 3612
rect 520372 604 520424 610
rect 520372 546 520424 552
rect 521476 604 521528 610
rect 521476 546 521528 552
rect 521488 480 521516 546
rect 522684 480 522712 3606
rect 523868 3596 523920 3602
rect 523868 3538 523920 3544
rect 523880 480 523908 3538
rect 525076 480 525104 3742
rect 525536 3602 525564 340054
rect 525616 336796 525668 336802
rect 525616 336738 525668 336744
rect 525628 3806 525656 336738
rect 525616 3800 525668 3806
rect 525616 3742 525668 3748
rect 525524 3596 525576 3602
rect 525524 3538 525576 3544
rect 525720 3369 525748 340068
rect 526364 336802 526392 340068
rect 526916 337686 526944 340068
rect 526904 337680 526956 337686
rect 526904 337622 526956 337628
rect 527560 336802 527588 340068
rect 528204 337385 528232 340068
rect 528190 337376 528246 337385
rect 528190 337311 528246 337320
rect 528756 336802 528784 340068
rect 528940 337606 529244 337634
rect 529400 337618 529428 340068
rect 529478 337784 529534 337793
rect 529478 337719 529534 337728
rect 528940 337550 528968 337606
rect 528928 337544 528980 337550
rect 528928 337486 528980 337492
rect 526352 336796 526404 336802
rect 526352 336738 526404 336744
rect 527548 336796 527600 336802
rect 527548 336738 527600 336744
rect 528468 336796 528520 336802
rect 528468 336738 528520 336744
rect 528744 336796 528796 336802
rect 528744 336738 528796 336744
rect 526442 204504 526498 204513
rect 526442 204439 526498 204448
rect 526456 204406 526484 204439
rect 526444 204400 526496 204406
rect 526444 204342 526496 204348
rect 526442 180976 526498 180985
rect 526442 180911 526498 180920
rect 526456 180878 526484 180911
rect 526444 180872 526496 180878
rect 526444 180814 526496 180820
rect 526442 169960 526498 169969
rect 526442 169895 526498 169904
rect 526456 169862 526484 169895
rect 526444 169856 526496 169862
rect 526444 169798 526496 169804
rect 526442 157584 526498 157593
rect 526442 157519 526498 157528
rect 526456 157486 526484 157519
rect 526444 157480 526496 157486
rect 526444 157422 526496 157428
rect 526442 134056 526498 134065
rect 526442 133991 526498 134000
rect 526456 133958 526484 133991
rect 526444 133952 526496 133958
rect 526444 133894 526496 133900
rect 526442 123040 526498 123049
rect 526442 122975 526498 122984
rect 526456 122942 526484 122975
rect 526444 122936 526496 122942
rect 526444 122878 526496 122884
rect 526442 110664 526498 110673
rect 526442 110599 526498 110608
rect 526456 110566 526484 110599
rect 526444 110560 526496 110566
rect 526444 110502 526496 110508
rect 526442 76120 526498 76129
rect 526442 76055 526498 76064
rect 526456 76022 526484 76055
rect 526444 76016 526496 76022
rect 526444 75958 526496 75964
rect 526442 63744 526498 63753
rect 526442 63679 526498 63688
rect 526456 63646 526484 63679
rect 526444 63640 526496 63646
rect 526444 63582 526496 63588
rect 526442 40216 526498 40225
rect 526442 40151 526498 40160
rect 526456 40118 526484 40151
rect 526444 40112 526496 40118
rect 526444 40054 526496 40060
rect 525890 29200 525946 29209
rect 525890 29135 525946 29144
rect 525904 29102 525932 29135
rect 525892 29096 525944 29102
rect 525892 29038 525944 29044
rect 526442 16824 526498 16833
rect 526442 16759 526498 16768
rect 526456 16726 526484 16759
rect 526444 16720 526496 16726
rect 526444 16662 526496 16668
rect 528480 3534 528508 336738
rect 526260 3528 526312 3534
rect 526260 3470 526312 3476
rect 528468 3528 528520 3534
rect 528468 3470 528520 3476
rect 525706 3360 525762 3369
rect 525706 3295 525762 3304
rect 526272 480 526300 3470
rect 528652 3460 528704 3466
rect 528652 3402 528704 3408
rect 527456 2848 527508 2854
rect 527456 2790 527508 2796
rect 527468 480 527496 2790
rect 528664 480 528692 3402
rect 529216 2854 529244 337606
rect 529388 337612 529440 337618
rect 529388 337554 529440 337560
rect 529492 337482 529520 337719
rect 529480 337476 529532 337482
rect 529480 337418 529532 337424
rect 529848 336796 529900 336802
rect 529848 336738 529900 336744
rect 529756 4956 529808 4962
rect 529756 4898 529808 4904
rect 529768 3346 529796 4898
rect 529860 3466 529888 336738
rect 530596 299470 530624 640766
rect 530674 637936 530730 637945
rect 530674 637871 530730 637880
rect 530688 322930 530716 637871
rect 530780 416770 530808 642806
rect 530860 641028 530912 641034
rect 530860 640970 530912 640976
rect 530872 440230 530900 640970
rect 530950 638344 531006 638353
rect 530950 638279 531006 638288
rect 530964 463690 530992 638279
rect 531056 499526 531084 642874
rect 531136 641096 531188 641102
rect 531136 641038 531188 641044
rect 531148 510610 531176 641038
rect 531240 546446 531268 642942
rect 580172 642796 580224 642802
rect 580172 642738 580224 642744
rect 579804 639736 579856 639742
rect 579804 639678 579856 639684
rect 579816 639441 579844 639678
rect 579802 639432 579858 639441
rect 579802 639367 579858 639376
rect 580080 627904 580132 627910
rect 580080 627846 580132 627852
rect 580092 627745 580120 627846
rect 580078 627736 580134 627745
rect 580078 627671 580134 627680
rect 580080 604444 580132 604450
rect 580080 604386 580132 604392
rect 580092 604217 580120 604386
rect 580078 604208 580134 604217
rect 580078 604143 580134 604152
rect 580080 593360 580132 593366
rect 580080 593302 580132 593308
rect 580092 592521 580120 593302
rect 580078 592512 580134 592521
rect 580078 592447 580134 592456
rect 580080 580984 580132 580990
rect 580080 580926 580132 580932
rect 580092 580825 580120 580926
rect 580078 580816 580134 580825
rect 580078 580751 580134 580760
rect 580080 557524 580132 557530
rect 580080 557466 580132 557472
rect 580092 557297 580120 557466
rect 580078 557288 580134 557297
rect 580078 557223 580134 557232
rect 531228 546440 531280 546446
rect 531228 546382 531280 546388
rect 580080 546440 580132 546446
rect 580080 546382 580132 546388
rect 580092 545601 580120 546382
rect 580078 545592 580134 545601
rect 580078 545527 580134 545536
rect 531136 510604 531188 510610
rect 531136 510546 531188 510552
rect 580080 510604 580132 510610
rect 580080 510546 580132 510552
rect 580092 510377 580120 510546
rect 580078 510368 580134 510377
rect 580078 510303 580134 510312
rect 531044 499520 531096 499526
rect 531044 499462 531096 499468
rect 580080 499520 580132 499526
rect 580080 499462 580132 499468
rect 580092 498681 580120 499462
rect 580078 498672 580134 498681
rect 580078 498607 580134 498616
rect 580184 486849 580212 642738
rect 580448 642728 580500 642734
rect 580448 642670 580500 642676
rect 580356 640756 580408 640762
rect 580356 640698 580408 640704
rect 580264 639328 580316 639334
rect 580264 639270 580316 639276
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 530952 463684 531004 463690
rect 530952 463626 531004 463632
rect 579804 463684 579856 463690
rect 579804 463626 579856 463632
rect 579816 463457 579844 463626
rect 579802 463448 579858 463457
rect 579802 463383 579858 463392
rect 530860 440224 530912 440230
rect 530860 440166 530912 440172
rect 580172 440224 580224 440230
rect 580172 440166 580224 440172
rect 580184 439929 580212 440166
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 530768 416764 530820 416770
rect 530768 416706 530820 416712
rect 580172 416764 580224 416770
rect 580172 416706 580224 416712
rect 580184 416537 580212 416706
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 579620 393304 579672 393310
rect 579620 393246 579672 393252
rect 579632 393009 579660 393246
rect 579618 393000 579674 393009
rect 579618 392935 579674 392944
rect 580172 346384 580224 346390
rect 580172 346326 580224 346332
rect 580184 346089 580212 346326
rect 580170 346080 580226 346089
rect 580170 346015 580226 346024
rect 547144 338088 547196 338094
rect 547144 338030 547196 338036
rect 531320 337408 531372 337414
rect 531320 337350 531372 337356
rect 530676 322924 530728 322930
rect 530676 322866 530728 322872
rect 530584 299464 530636 299470
rect 530584 299406 530636 299412
rect 529848 3460 529900 3466
rect 529848 3402 529900 3408
rect 531332 3346 531360 337350
rect 540244 337204 540296 337210
rect 540244 337146 540296 337152
rect 538220 337136 538272 337142
rect 538220 337078 538272 337084
rect 534080 336932 534132 336938
rect 534080 336874 534132 336880
rect 534092 3346 534120 336874
rect 536102 87408 536158 87417
rect 536102 87343 536158 87352
rect 536116 87009 536144 87343
rect 536102 87000 536158 87009
rect 536102 86935 536158 86944
rect 536932 4820 536984 4826
rect 536932 4762 536984 4768
rect 529768 3318 529888 3346
rect 531332 3318 532280 3346
rect 534092 3318 534580 3346
rect 529204 2848 529256 2854
rect 529204 2790 529256 2796
rect 529860 480 529888 3318
rect 531044 2916 531096 2922
rect 531044 2858 531096 2864
rect 531056 480 531084 2858
rect 532252 480 532280 3318
rect 533436 2984 533488 2990
rect 533436 2926 533488 2932
rect 533448 480 533476 2926
rect 534552 480 534580 3318
rect 535736 3052 535788 3058
rect 535736 2994 535788 3000
rect 535748 480 535776 2994
rect 536944 480 536972 4762
rect 538232 3346 538260 337078
rect 538232 3318 539364 3346
rect 540256 3330 540284 337146
rect 540336 337068 540388 337074
rect 540336 337010 540388 337016
rect 538128 3120 538180 3126
rect 538128 3062 538180 3068
rect 538140 480 538168 3062
rect 539336 480 539364 3318
rect 540244 3324 540296 3330
rect 540244 3266 540296 3272
rect 540348 3262 540376 337010
rect 545764 337000 545816 337006
rect 545764 336942 545816 336948
rect 543004 336864 543056 336870
rect 543004 336806 543056 336812
rect 540886 204776 540942 204785
rect 540886 204711 540942 204720
rect 540900 204377 540928 204711
rect 540886 204368 540942 204377
rect 540886 204303 540942 204312
rect 540886 181248 540942 181257
rect 540886 181183 540942 181192
rect 540900 180849 540928 181183
rect 540886 180840 540942 180849
rect 540886 180775 540942 180784
rect 540886 170232 540942 170241
rect 540886 170167 540942 170176
rect 540900 169833 540928 170167
rect 540886 169824 540942 169833
rect 540886 169759 540942 169768
rect 540886 157856 540942 157865
rect 540886 157791 540942 157800
rect 540900 157457 540928 157791
rect 540886 157448 540942 157457
rect 540886 157383 540942 157392
rect 540886 134328 540942 134337
rect 540886 134263 540942 134272
rect 540900 133929 540928 134263
rect 540886 133920 540942 133929
rect 540886 133855 540942 133864
rect 540886 123312 540942 123321
rect 540886 123247 540942 123256
rect 540900 122913 540928 123247
rect 540886 122904 540942 122913
rect 540886 122839 540942 122848
rect 540886 110936 540942 110945
rect 540886 110871 540942 110880
rect 540900 110537 540928 110871
rect 540886 110528 540942 110537
rect 540886 110463 540942 110472
rect 540886 76392 540942 76401
rect 540886 76327 540942 76336
rect 540900 75993 540928 76327
rect 540886 75984 540942 75993
rect 540886 75919 540942 75928
rect 540886 64016 540942 64025
rect 540886 63951 540942 63960
rect 540900 63617 540928 63951
rect 540886 63608 540942 63617
rect 540886 63543 540942 63552
rect 540886 40488 540942 40497
rect 540886 40423 540942 40432
rect 540900 40089 540928 40423
rect 540886 40080 540942 40089
rect 540886 40015 540942 40024
rect 540794 29472 540850 29481
rect 540794 29407 540850 29416
rect 540808 29050 540836 29407
rect 540886 29064 540942 29073
rect 540808 29022 540886 29050
rect 540886 28999 540942 29008
rect 540886 17096 540942 17105
rect 540886 17031 540942 17040
rect 540900 16697 540928 17031
rect 540886 16688 540942 16697
rect 540886 16623 540942 16632
rect 540520 4888 540572 4894
rect 540520 4830 540572 4836
rect 540336 3256 540388 3262
rect 540336 3198 540388 3204
rect 540532 480 540560 4830
rect 542912 3324 542964 3330
rect 542912 3266 542964 3272
rect 541716 2848 541768 2854
rect 541716 2790 541768 2796
rect 541728 480 541756 2790
rect 542924 480 542952 3266
rect 543016 2922 543044 336806
rect 545672 274984 545724 274990
rect 545670 274952 545672 274961
rect 545724 274952 545726 274961
rect 545670 274887 545726 274896
rect 545776 3262 545804 336942
rect 544108 3256 544160 3262
rect 544108 3198 544160 3204
rect 545764 3256 545816 3262
rect 545764 3198 545816 3204
rect 543004 2916 543056 2922
rect 543004 2858 543056 2864
rect 544120 480 544148 3198
rect 547156 3194 547184 338030
rect 547236 338020 547288 338026
rect 547236 337962 547288 337968
rect 547248 3330 547276 337962
rect 556804 337952 556856 337958
rect 556804 337894 556856 337900
rect 553400 337884 553452 337890
rect 553400 337826 553452 337832
rect 549904 337340 549956 337346
rect 549904 337282 549956 337288
rect 547236 3324 547288 3330
rect 547236 3266 547288 3272
rect 549916 3194 549944 337282
rect 550548 274984 550600 274990
rect 550546 274952 550548 274961
rect 550600 274952 550602 274961
rect 550546 274887 550602 274896
rect 553308 181008 553360 181014
rect 553306 180976 553308 180985
rect 553360 180976 553362 180985
rect 553306 180911 553362 180920
rect 552388 3392 552440 3398
rect 552388 3334 552440 3340
rect 553412 3346 553440 337826
rect 554872 337816 554924 337822
rect 554872 337758 554924 337764
rect 554884 3346 554912 337758
rect 554964 181008 555016 181014
rect 554962 180976 554964 180985
rect 555016 180976 555018 180985
rect 554962 180911 555018 180920
rect 556816 3398 556844 337894
rect 560300 337748 560352 337754
rect 560300 337690 560352 337696
rect 558184 337272 558236 337278
rect 558184 337214 558236 337220
rect 558196 4146 558224 337214
rect 560206 204640 560262 204649
rect 560206 204575 560262 204584
rect 560220 204241 560248 204575
rect 560206 204232 560262 204241
rect 560206 204167 560262 204176
rect 560206 170096 560262 170105
rect 560206 170031 560262 170040
rect 560220 169697 560248 170031
rect 560206 169688 560262 169697
rect 560206 169623 560262 169632
rect 560206 157720 560262 157729
rect 560206 157655 560262 157664
rect 560220 157321 560248 157655
rect 560206 157312 560262 157321
rect 560206 157247 560262 157256
rect 560206 134192 560262 134201
rect 560206 134127 560262 134136
rect 560220 133793 560248 134127
rect 560206 133784 560262 133793
rect 560206 133719 560262 133728
rect 560206 123176 560262 123185
rect 560206 123111 560262 123120
rect 560220 122777 560248 123111
rect 560206 122768 560262 122777
rect 560206 122703 560262 122712
rect 560206 110800 560262 110809
rect 560206 110735 560262 110744
rect 560220 110401 560248 110735
rect 560206 110392 560262 110401
rect 560206 110327 560262 110336
rect 560206 87544 560262 87553
rect 560206 87479 560262 87488
rect 560220 87281 560248 87479
rect 560206 87272 560262 87281
rect 560206 87207 560262 87216
rect 560206 76256 560262 76265
rect 560206 76191 560262 76200
rect 560220 75857 560248 76191
rect 560206 75848 560262 75857
rect 560206 75783 560262 75792
rect 560206 63880 560262 63889
rect 560206 63815 560262 63824
rect 560220 63481 560248 63815
rect 560206 63472 560262 63481
rect 560206 63407 560262 63416
rect 560206 40352 560262 40361
rect 560206 40287 560262 40296
rect 560220 39953 560248 40287
rect 560206 39944 560262 39953
rect 560206 39879 560262 39888
rect 560206 29608 560262 29617
rect 560206 29543 560262 29552
rect 560220 29345 560248 29543
rect 560206 29336 560262 29345
rect 560206 29271 560262 29280
rect 560206 16960 560262 16969
rect 560206 16895 560262 16904
rect 560220 16561 560248 16895
rect 560206 16552 560262 16561
rect 560206 16487 560262 16496
rect 557172 4140 557224 4146
rect 557172 4082 557224 4088
rect 558184 4140 558236 4146
rect 558184 4082 558236 4088
rect 556804 3392 556856 3398
rect 550088 3324 550140 3330
rect 550088 3266 550140 3272
rect 545304 3188 545356 3194
rect 545304 3130 545356 3136
rect 547144 3188 547196 3194
rect 547144 3130 547196 3136
rect 548892 3188 548944 3194
rect 548892 3130 548944 3136
rect 549904 3188 549956 3194
rect 549904 3130 549956 3136
rect 545316 480 545344 3130
rect 547696 3120 547748 3126
rect 547696 3062 547748 3068
rect 546500 3052 546552 3058
rect 546500 2994 546552 3000
rect 546512 480 546540 2994
rect 547708 480 547736 3062
rect 548904 480 548932 3130
rect 550100 480 550128 3266
rect 551192 3120 551244 3126
rect 551192 3062 551244 3068
rect 551204 480 551232 3062
rect 552400 480 552428 3334
rect 553412 3318 553624 3346
rect 554884 3318 556016 3346
rect 556804 3334 556856 3340
rect 553596 480 553624 3318
rect 554780 3256 554832 3262
rect 554780 3198 554832 3204
rect 554792 480 554820 3198
rect 555988 480 556016 3318
rect 557184 480 557212 4082
rect 559564 4072 559616 4078
rect 559564 4014 559616 4020
rect 558368 3324 558420 3330
rect 558368 3266 558420 3272
rect 558380 480 558408 3266
rect 559576 480 559604 4014
rect 560312 3482 560340 337690
rect 563152 337680 563204 337686
rect 563152 337622 563204 337628
rect 563058 274952 563114 274961
rect 563058 274887 563114 274896
rect 563072 274553 563100 274887
rect 563058 274544 563114 274553
rect 563058 274479 563114 274488
rect 561956 4004 562008 4010
rect 561956 3946 562008 3952
rect 560312 3454 560800 3482
rect 560772 480 560800 3454
rect 561968 480 561996 3946
rect 563164 480 563192 337622
rect 573364 337612 573416 337618
rect 573364 337554 573416 337560
rect 567200 337544 567252 337550
rect 567200 337486 567252 337492
rect 565082 337376 565138 337385
rect 565082 337311 565138 337320
rect 565096 3942 565124 337311
rect 564348 3936 564400 3942
rect 564348 3878 564400 3884
rect 565084 3936 565136 3942
rect 565084 3878 565136 3884
rect 564360 480 564388 3878
rect 566740 3868 566792 3874
rect 566740 3810 566792 3816
rect 565544 3392 565596 3398
rect 565544 3334 565596 3340
rect 565556 480 565584 3334
rect 566752 480 566780 3810
rect 567212 3346 567240 337486
rect 569224 337476 569276 337482
rect 569224 337418 569276 337424
rect 569040 3732 569092 3738
rect 569040 3674 569092 3680
rect 567212 3318 567884 3346
rect 567856 480 567884 3318
rect 569052 480 569080 3674
rect 569236 3534 569264 337418
rect 571984 337408 572036 337414
rect 571984 337350 572036 337356
rect 571432 3664 571484 3670
rect 571432 3606 571484 3612
rect 569224 3528 569276 3534
rect 569224 3470 569276 3476
rect 570236 3528 570288 3534
rect 570236 3470 570288 3476
rect 570248 480 570276 3470
rect 571444 480 571472 3606
rect 571996 3058 572024 337350
rect 572626 274816 572682 274825
rect 572682 274774 572760 274802
rect 572626 274751 572682 274760
rect 572732 274689 572760 274774
rect 572718 274680 572774 274689
rect 572718 274615 572774 274624
rect 572626 204504 572682 204513
rect 572626 204439 572682 204448
rect 572640 204354 572668 204439
rect 572718 204368 572774 204377
rect 572640 204326 572718 204354
rect 572718 204303 572774 204312
rect 572626 169960 572682 169969
rect 572626 169895 572682 169904
rect 572640 169810 572668 169895
rect 572718 169824 572774 169833
rect 572640 169782 572718 169810
rect 572718 169759 572774 169768
rect 572626 157584 572682 157593
rect 572626 157519 572682 157528
rect 572640 157434 572668 157519
rect 572718 157448 572774 157457
rect 572640 157406 572718 157434
rect 572718 157383 572774 157392
rect 572626 134056 572682 134065
rect 572626 133991 572682 134000
rect 572640 133906 572668 133991
rect 572718 133920 572774 133929
rect 572640 133878 572718 133906
rect 572718 133855 572774 133864
rect 572626 123040 572682 123049
rect 572626 122975 572682 122984
rect 572640 122890 572668 122975
rect 572718 122904 572774 122913
rect 572640 122862 572718 122890
rect 572718 122839 572774 122848
rect 572626 110664 572682 110673
rect 572626 110599 572682 110608
rect 572640 110514 572668 110599
rect 572718 110528 572774 110537
rect 572640 110486 572718 110514
rect 572718 110463 572774 110472
rect 572626 87136 572682 87145
rect 572626 87071 572628 87080
rect 572680 87071 572682 87080
rect 572628 87042 572680 87048
rect 572626 76120 572682 76129
rect 572626 76055 572682 76064
rect 572640 75970 572668 76055
rect 572718 75984 572774 75993
rect 572640 75942 572718 75970
rect 572718 75919 572774 75928
rect 572626 63744 572682 63753
rect 572626 63679 572682 63688
rect 572640 63594 572668 63679
rect 572718 63608 572774 63617
rect 572640 63566 572718 63594
rect 572718 63543 572774 63552
rect 572626 40216 572682 40225
rect 572626 40151 572682 40160
rect 572640 40066 572668 40151
rect 572718 40080 572774 40089
rect 572640 40038 572718 40066
rect 572718 40015 572774 40024
rect 572628 29232 572680 29238
rect 572626 29200 572628 29209
rect 572680 29200 572682 29209
rect 572626 29135 572682 29144
rect 572626 16824 572682 16833
rect 572626 16759 572682 16768
rect 572640 16674 572668 16759
rect 572718 16688 572774 16697
rect 572640 16646 572718 16674
rect 572718 16623 572774 16632
rect 572628 3800 572680 3806
rect 572628 3742 572680 3748
rect 571984 3052 572036 3058
rect 571984 2994 572036 3000
rect 572640 480 572668 3742
rect 573376 3602 573404 337554
rect 579620 322924 579672 322930
rect 579620 322866 579672 322872
rect 579632 322697 579660 322866
rect 579618 322688 579674 322697
rect 579618 322623 579674 322632
rect 579712 299464 579764 299470
rect 579712 299406 579764 299412
rect 579724 299169 579752 299406
rect 579710 299160 579766 299169
rect 579710 299095 579766 299104
rect 580276 217025 580304 639270
rect 580368 228857 580396 640698
rect 580460 252249 580488 642670
rect 580908 639668 580960 639674
rect 580908 639610 580960 639616
rect 580816 639600 580868 639606
rect 580816 639542 580868 639548
rect 580724 639532 580776 639538
rect 580724 639474 580776 639480
rect 580632 639464 580684 639470
rect 580632 639406 580684 639412
rect 580540 639396 580592 639402
rect 580540 639338 580592 639344
rect 580552 263945 580580 639338
rect 580644 310865 580672 639406
rect 580736 357921 580764 639474
rect 580828 404841 580856 639542
rect 580920 451761 580948 639610
rect 580906 451752 580962 451761
rect 580906 451687 580962 451696
rect 580814 404832 580870 404841
rect 580814 404767 580870 404776
rect 580722 357912 580778 357921
rect 580722 357847 580778 357856
rect 580630 310856 580686 310865
rect 580630 310791 580686 310800
rect 580538 263936 580594 263945
rect 580538 263871 580594 263880
rect 580446 252240 580502 252249
rect 580446 252175 580502 252184
rect 580354 228848 580410 228857
rect 580354 228783 580410 228792
rect 580262 217016 580318 217025
rect 580262 216951 580318 216960
rect 576766 87136 576822 87145
rect 576766 87071 576768 87080
rect 576820 87071 576822 87080
rect 576768 87042 576820 87048
rect 576768 29232 576820 29238
rect 576766 29200 576768 29209
rect 576820 29200 576822 29209
rect 576766 29135 576822 29144
rect 576216 4140 576268 4146
rect 576216 4082 576268 4088
rect 573364 3596 573416 3602
rect 573364 3538 573416 3544
rect 573824 3528 573876 3534
rect 573824 3470 573876 3476
rect 573836 480 573864 3470
rect 575018 3360 575074 3369
rect 575018 3295 575074 3304
rect 575032 480 575060 3295
rect 576228 480 576256 4082
rect 579804 3936 579856 3942
rect 579804 3878 579856 3884
rect 578608 3392 578660 3398
rect 578608 3334 578660 3340
rect 577412 3052 577464 3058
rect 577412 2994 577464 3000
rect 577424 480 577452 2994
rect 578620 480 578648 3334
rect 579816 480 579844 3878
rect 582196 3596 582248 3602
rect 582196 3538 582248 3544
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 3538
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8114 700304 8170 700360
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3514 642912 3570 642968
rect 3146 624824 3202 624880
rect 2778 610408 2834 610464
rect 3146 596028 3148 596048
rect 3148 596028 3200 596048
rect 3200 596028 3202 596048
rect 3146 595992 3202 596028
rect 3146 567296 3202 567352
rect 2778 553052 2780 553072
rect 2780 553052 2832 553072
rect 2832 553052 2834 553072
rect 2778 553016 2834 553052
rect 3238 538600 3294 538656
rect 3238 509904 3294 509960
rect 2778 495488 2834 495544
rect 3238 481072 3294 481128
rect 3146 452412 3148 452432
rect 3148 452412 3200 452432
rect 3200 452412 3202 452432
rect 3146 452376 3202 452412
rect 2778 437996 2780 438016
rect 2780 437996 2832 438016
rect 2832 437996 2834 438016
rect 2778 437960 2834 437996
rect 3238 423680 3294 423736
rect 3422 638152 3478 638208
rect 3330 394984 3386 395040
rect 3238 380604 3240 380624
rect 3240 380604 3292 380624
rect 3292 380604 3294 380624
rect 3238 380568 3294 380604
rect 2778 366152 2834 366208
rect 3330 337492 3332 337512
rect 3332 337492 3384 337512
rect 3384 337492 3386 337512
rect 3330 337456 3386 337492
rect 3146 324264 3202 324320
rect 3146 323040 3202 323096
rect 2778 308796 2780 308816
rect 2780 308796 2832 308816
rect 2832 308796 2834 308816
rect 2778 308760 2834 308796
rect 3330 294344 3386 294400
rect 3146 280100 3148 280120
rect 3148 280100 3200 280120
rect 3200 280100 3202 280120
rect 3146 280064 3202 280100
rect 3146 252456 3202 252512
rect 3146 251232 3202 251288
rect 2778 236952 2834 237008
rect 3330 180648 3386 180704
rect 3330 179424 3386 179480
rect 2778 165008 2834 165064
rect 3330 151680 3386 151736
rect 3330 150728 3386 150784
rect 2962 122032 3018 122088
rect 3330 78920 3386 78976
rect 3698 638288 3754 638344
rect 4066 222536 4122 222592
rect 3974 193840 4030 193896
rect 4894 638424 4950 638480
rect 5078 638560 5134 638616
rect 5262 638696 5318 638752
rect 3882 136312 3938 136368
rect 6918 638424 6974 638480
rect 6918 638016 6974 638072
rect 3790 107616 3846 107672
rect 3698 93200 3754 93256
rect 3606 64504 3662 64560
rect 3514 50088 3570 50144
rect 288898 641960 288954 642016
rect 317786 642776 317842 642832
rect 414018 700304 414074 700360
rect 580170 697992 580226 698048
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 517794 642912 517850 642968
rect 473082 642640 473138 642696
rect 478326 642504 478382 642560
rect 483662 642368 483718 642424
rect 491482 642232 491538 642288
rect 494150 642096 494206 642152
rect 504638 641824 504694 641880
rect 231398 639240 231454 639296
rect 233974 639240 234030 639296
rect 236550 639240 236606 639296
rect 239126 639240 239182 639296
rect 241886 639240 241942 639296
rect 244002 639240 244058 639296
rect 246946 639240 247002 639296
rect 249154 639240 249210 639296
rect 252282 639240 252338 639296
rect 254950 639240 255006 639296
rect 257710 639240 257766 639296
rect 260286 639240 260342 639296
rect 262862 639240 262918 639296
rect 398102 639648 398158 639704
rect 420182 639648 420238 639704
rect 398102 639376 398158 639432
rect 273166 639240 273222 639296
rect 281170 639240 281226 639296
rect 304906 639240 304962 639296
rect 338026 639240 338082 639296
rect 420182 639240 420238 639296
rect 430762 639240 430818 639296
rect 457166 639240 457222 639296
rect 462318 639240 462374 639296
rect 488630 639240 488686 639296
rect 509790 639240 509846 639296
rect 525430 639240 525486 639296
rect 528098 639240 528154 639296
rect 8114 638832 8170 638888
rect 17406 638832 17462 638888
rect 26146 638832 26202 638888
rect 36726 638832 36782 638888
rect 45466 638832 45522 638888
rect 56046 638832 56102 638888
rect 64786 638832 64842 638888
rect 75366 638832 75422 638888
rect 84106 638832 84162 638888
rect 94686 638832 94742 638888
rect 103426 638832 103482 638888
rect 114006 638832 114062 638888
rect 122746 638832 122802 638888
rect 133326 638832 133382 638888
rect 142066 638832 142122 638888
rect 152646 638832 152702 638888
rect 161386 638832 161442 638888
rect 171966 638832 172022 638888
rect 180706 638832 180762 638888
rect 191286 638832 191342 638888
rect 200026 638832 200082 638888
rect 210606 638832 210662 638888
rect 219990 638832 220046 638888
rect 17222 638424 17278 638480
rect 26238 638424 26294 638480
rect 36542 638424 36598 638480
rect 45558 638424 45614 638480
rect 55862 638424 55918 638480
rect 64878 638424 64934 638480
rect 75182 638424 75238 638480
rect 84198 638424 84254 638480
rect 94502 638424 94558 638480
rect 103518 638424 103574 638480
rect 113822 638424 113878 638480
rect 122838 638424 122894 638480
rect 133142 638424 133198 638480
rect 142158 638424 142214 638480
rect 152462 638424 152518 638480
rect 161478 638424 161534 638480
rect 171782 638424 171838 638480
rect 180798 638424 180854 638480
rect 191102 638424 191158 638480
rect 200118 638424 200174 638480
rect 210422 638424 210478 638480
rect 220082 638424 220138 638480
rect 17222 638016 17278 638072
rect 17406 638016 17462 638072
rect 26146 638016 26202 638072
rect 26330 638016 26386 638072
rect 36542 638016 36598 638072
rect 36726 638016 36782 638072
rect 45466 638016 45522 638072
rect 45650 638016 45706 638072
rect 55862 638016 55918 638072
rect 56046 638016 56102 638072
rect 64786 638016 64842 638072
rect 64970 638016 65026 638072
rect 75182 638016 75238 638072
rect 75366 638016 75422 638072
rect 84106 638016 84162 638072
rect 84290 638016 84346 638072
rect 94502 638016 94558 638072
rect 94686 638016 94742 638072
rect 103426 638016 103482 638072
rect 103610 638016 103666 638072
rect 113822 638016 113878 638072
rect 114006 638016 114062 638072
rect 122746 638016 122802 638072
rect 122930 638016 122986 638072
rect 133142 638016 133198 638072
rect 133326 638016 133382 638072
rect 142066 638016 142122 638072
rect 142250 638016 142306 638072
rect 152462 638016 152518 638072
rect 152646 638016 152702 638072
rect 161386 638016 161442 638072
rect 161570 638016 161626 638072
rect 171782 638016 171838 638072
rect 171966 638016 172022 638072
rect 180706 638016 180762 638072
rect 180890 638016 180946 638072
rect 191102 638016 191158 638072
rect 191286 638016 191342 638072
rect 200026 638016 200082 638072
rect 200210 638016 200266 638072
rect 210422 638016 210478 638072
rect 210606 638016 210662 638072
rect 219990 638016 220046 638072
rect 220082 637880 220138 637936
rect 530306 638832 530362 638888
rect 10322 337320 10378 337376
rect 3514 35844 3516 35864
rect 3516 35844 3568 35864
rect 3568 35844 3570 35864
rect 3514 35808 3570 35844
rect 3422 7112 3478 7168
rect 6458 3304 6514 3360
rect 48134 6160 48190 6216
rect 60646 10240 60702 10296
rect 136086 8880 136142 8936
rect 134890 7520 134946 7576
rect 219346 4800 219402 4856
rect 232410 337320 232466 337376
rect 231858 3304 231914 3360
rect 234342 336504 234398 336560
rect 234342 327120 234398 327176
rect 234250 303048 234306 303104
rect 234250 299648 234306 299704
rect 233974 261976 234030 262032
rect 235998 253952 236054 254008
rect 233974 252592 234030 252648
rect 234342 206896 234398 206952
rect 234342 197512 234398 197568
rect 234526 187448 234582 187504
rect 234526 178064 234582 178120
rect 234342 138624 234398 138680
rect 234342 121760 234398 121816
rect 234710 121352 234766 121408
rect 234710 112920 234766 112976
rect 236274 295316 236330 295352
rect 236274 295296 236276 295316
rect 236276 295296 236328 295316
rect 236328 295296 236330 295316
rect 236550 295296 236606 295352
rect 236458 276120 236514 276176
rect 236274 275984 236330 276040
rect 236274 253952 236330 254008
rect 236458 162968 236514 163024
rect 236274 162832 236330 162888
rect 236366 134000 236422 134056
rect 236274 133864 236330 133920
rect 240230 154672 240286 154728
rect 240230 154536 240286 154592
rect 240322 143520 240378 143576
rect 240506 143520 240562 143576
rect 240046 64912 240102 64968
rect 240046 43832 240102 43888
rect 240046 40160 240102 40216
rect 240138 16768 240194 16824
rect 240230 16632 240286 16688
rect 242714 240080 242770 240136
rect 241794 183504 241850 183560
rect 241978 183504 242034 183560
rect 241794 96600 241850 96656
rect 241978 96600 242034 96656
rect 243174 280064 243230 280120
rect 243358 280064 243414 280120
rect 243358 270680 243414 270736
rect 243082 270544 243138 270600
rect 243174 260752 243230 260808
rect 243358 260752 243414 260808
rect 243358 251368 243414 251424
rect 243082 251232 243138 251288
rect 242990 240080 243046 240136
rect 243082 183640 243138 183696
rect 243266 183504 243322 183560
rect 244462 135360 244518 135416
rect 243082 135244 243138 135280
rect 243082 135224 243084 135244
rect 243084 135224 243136 135244
rect 243136 135224 243138 135244
rect 243266 135244 243322 135280
rect 243266 135224 243268 135244
rect 243268 135224 243320 135244
rect 243320 135224 243322 135244
rect 244462 135088 244518 135144
rect 248326 63552 248382 63608
rect 249982 125840 250038 125896
rect 249982 125568 250038 125624
rect 251086 17040 251142 17096
rect 251086 16632 251142 16688
rect 252558 153176 252614 153232
rect 252558 125296 252614 125352
rect 252742 231784 252798 231840
rect 252926 231784 252982 231840
rect 252742 212508 252744 212528
rect 252744 212508 252796 212528
rect 252796 212508 252798 212528
rect 252742 212472 252798 212508
rect 252926 212472 252982 212528
rect 252834 202816 252890 202872
rect 253018 202816 253074 202872
rect 252834 193196 252836 193216
rect 252836 193196 252888 193216
rect 252888 193196 252890 193216
rect 252834 193160 252890 193196
rect 253018 193196 253020 193216
rect 253020 193196 253072 193216
rect 253072 193196 253074 193216
rect 253018 193160 253074 193196
rect 252834 153176 252890 153232
rect 252926 125568 252982 125624
rect 253110 76472 253166 76528
rect 253110 75928 253166 75984
rect 253110 64232 253166 64288
rect 253110 63280 253166 63336
rect 254030 267688 254086 267744
rect 254214 267688 254270 267744
rect 254030 258032 254086 258088
rect 254214 258032 254270 258088
rect 255318 201456 255374 201512
rect 255594 201476 255650 201512
rect 255594 201456 255596 201476
rect 255596 201456 255648 201476
rect 255648 201456 255650 201476
rect 254122 193160 254178 193216
rect 254306 193160 254362 193216
rect 255502 55120 255558 55176
rect 255778 55120 255834 55176
rect 253938 6160 253994 6216
rect 257986 86944 258042 87000
rect 257986 86808 258042 86864
rect 259366 238720 259422 238776
rect 259366 87080 259422 87136
rect 259366 86808 259422 86864
rect 261022 318960 261078 319016
rect 261022 318824 261078 318880
rect 261022 307672 261078 307728
rect 261206 307672 261262 307728
rect 259550 267688 259606 267744
rect 259734 267688 259790 267744
rect 259550 258032 259606 258088
rect 259734 258032 259790 258088
rect 259550 238720 259606 238776
rect 259642 193160 259698 193216
rect 259826 193160 259882 193216
rect 259734 10240 259790 10296
rect 265070 278704 265126 278760
rect 265346 278704 265402 278760
rect 265254 177248 265310 177304
rect 266818 240080 266874 240136
rect 267094 240080 267150 240136
rect 266726 230424 266782 230480
rect 267094 230424 267150 230480
rect 267002 183504 267058 183560
rect 267186 183504 267242 183560
rect 266450 173884 266452 173904
rect 266452 173884 266504 173904
rect 266504 173884 266506 173904
rect 266450 173848 266506 173884
rect 266634 173848 266690 173904
rect 265254 164212 265310 164248
rect 265254 164192 265256 164212
rect 265256 164192 265308 164212
rect 265308 164192 265310 164212
rect 267002 164212 267058 164248
rect 267002 164192 267004 164212
rect 267004 164192 267056 164212
rect 267056 164192 267058 164212
rect 267186 164192 267242 164248
rect 266910 154536 266966 154592
rect 267094 154536 267150 154592
rect 266542 145016 266598 145072
rect 266450 144880 266506 144936
rect 265162 135360 265218 135416
rect 265162 135224 265218 135280
rect 267738 134136 267794 134192
rect 267738 134000 267794 134056
rect 265070 115912 265126 115968
rect 265254 115912 265310 115968
rect 267738 87116 267740 87136
rect 267740 87116 267792 87136
rect 267792 87116 267794 87136
rect 267738 87080 267794 87116
rect 266450 82728 266506 82784
rect 266634 82592 266690 82648
rect 267646 63860 267648 63880
rect 267648 63860 267700 63880
rect 267700 63860 267702 63880
rect 267646 63824 267702 63860
rect 267738 40332 267740 40352
rect 267740 40332 267792 40352
rect 267792 40332 267794 40352
rect 267738 40296 267794 40332
rect 268934 171264 268990 171320
rect 268934 170040 268990 170096
rect 270774 260752 270830 260808
rect 270958 260752 271014 260808
rect 271878 241440 271934 241496
rect 272062 241440 272118 241496
rect 271878 222128 271934 222184
rect 272062 222128 272118 222184
rect 270682 135224 270738 135280
rect 270866 135224 270922 135280
rect 271878 125568 271934 125624
rect 272062 125588 272118 125624
rect 272062 125568 272064 125588
rect 272064 125568 272116 125588
rect 272116 125568 272118 125588
rect 270774 95376 270830 95432
rect 270682 95240 270738 95296
rect 273718 87116 273720 87136
rect 273720 87116 273772 87136
rect 273772 87116 273774 87136
rect 273718 87080 273774 87116
rect 274086 29144 274142 29200
rect 274270 29144 274326 29200
rect 275926 63860 275928 63880
rect 275928 63860 275980 63880
rect 275980 63860 275982 63880
rect 275926 63824 275982 63860
rect 277306 318824 277362 318880
rect 277582 318824 277638 318880
rect 277674 270408 277730 270464
rect 277766 270272 277822 270328
rect 278686 208528 278742 208584
rect 278686 204584 278742 204640
rect 278686 157528 278742 157584
rect 278686 157392 278742 157448
rect 278686 134136 278742 134192
rect 278686 133864 278742 133920
rect 277582 116048 277638 116104
rect 277490 115932 277546 115968
rect 277490 115912 277492 115932
rect 277492 115912 277544 115932
rect 277544 115912 277546 115932
rect 278778 110880 278834 110936
rect 278778 110472 278834 110528
rect 277306 63824 277362 63880
rect 277306 63552 277362 63608
rect 277306 40332 277308 40352
rect 277308 40332 277360 40352
rect 277360 40332 277362 40352
rect 277306 40296 277362 40332
rect 278686 40296 278742 40352
rect 278686 40024 278742 40080
rect 278778 29180 278780 29200
rect 278780 29180 278832 29200
rect 278832 29180 278834 29200
rect 278778 29144 278834 29180
rect 281630 289720 281686 289776
rect 281906 289720 281962 289776
rect 281906 238720 281962 238776
rect 282182 238720 282238 238776
rect 281722 202852 281724 202872
rect 281724 202852 281776 202872
rect 281776 202852 281778 202872
rect 281722 202816 281778 202852
rect 281906 202852 281908 202872
rect 281908 202852 281960 202872
rect 281960 202852 281962 202872
rect 281906 202816 281962 202852
rect 281998 183640 282054 183696
rect 281998 183368 282054 183424
rect 283102 154672 283158 154728
rect 283102 154536 283158 154592
rect 283102 125704 283158 125760
rect 283102 125568 283158 125624
rect 281630 106276 281686 106312
rect 281630 106256 281632 106276
rect 281632 106256 281684 106276
rect 281684 106256 281686 106276
rect 281814 106256 281870 106312
rect 283470 75964 283472 75984
rect 283472 75964 283524 75984
rect 283524 75964 283526 75984
rect 283470 75928 283526 75964
rect 283102 29180 283104 29200
rect 283104 29180 283156 29200
rect 283156 29180 283158 29200
rect 283102 29144 283158 29180
rect 287242 278704 287298 278760
rect 287426 278704 287482 278760
rect 287242 259392 287298 259448
rect 287334 259256 287390 259312
rect 287150 249736 287206 249792
rect 287426 249736 287482 249792
rect 287334 211248 287390 211304
rect 287242 211112 287298 211168
rect 287150 201456 287206 201512
rect 287334 201476 287390 201512
rect 287334 201456 287336 201476
rect 287336 201456 287388 201476
rect 287388 201456 287390 201476
rect 287242 172488 287298 172544
rect 287426 172488 287482 172544
rect 287242 145016 287298 145072
rect 287242 144880 287298 144936
rect 287242 125704 287298 125760
rect 287242 125568 287298 125624
rect 288438 222128 288494 222184
rect 288622 222128 288678 222184
rect 289818 204720 289874 204776
rect 289818 204448 289874 204504
rect 288438 202816 288494 202872
rect 288622 202816 288678 202872
rect 288438 183504 288494 183560
rect 288622 183504 288678 183560
rect 288346 170076 288348 170096
rect 288348 170076 288400 170096
rect 288400 170076 288402 170096
rect 288346 170040 288402 170076
rect 288622 125704 288678 125760
rect 288622 125568 288678 125624
rect 290554 75792 290610 75848
rect 293222 327256 293278 327312
rect 292762 327120 292818 327176
rect 292670 269184 292726 269240
rect 292946 269184 293002 269240
rect 292762 193196 292764 193216
rect 292764 193196 292816 193216
rect 292816 193196 292818 193216
rect 292762 193160 292818 193196
rect 292946 193196 292948 193216
rect 292948 193196 293000 193216
rect 293000 193196 293002 193216
rect 292946 193160 293002 193196
rect 293222 29280 293278 29336
rect 293222 28872 293278 28928
rect 294142 325624 294198 325680
rect 294326 325624 294382 325680
rect 293958 241440 294014 241496
rect 294142 241440 294198 241496
rect 293958 222128 294014 222184
rect 294142 222128 294198 222184
rect 294142 125704 294198 125760
rect 294050 125568 294106 125624
rect 295246 134136 295302 134192
rect 295246 133592 295302 133648
rect 296626 170076 296628 170096
rect 296628 170076 296680 170096
rect 296680 170076 296682 170096
rect 296626 170040 296682 170076
rect 295522 135224 295578 135280
rect 295706 135224 295762 135280
rect 298006 170040 298062 170096
rect 298006 169768 298062 169824
rect 298006 134156 298062 134192
rect 298006 134136 298008 134156
rect 298008 134136 298060 134156
rect 298060 134136 298062 134156
rect 298006 110744 298062 110800
rect 298006 110472 298062 110528
rect 298282 278704 298338 278760
rect 298558 278704 298614 278760
rect 298190 172488 298246 172544
rect 298466 172488 298522 172544
rect 299386 169668 299388 169688
rect 299388 169668 299440 169688
rect 299440 169668 299442 169688
rect 299386 169632 299442 169668
rect 298282 144900 298338 144936
rect 298282 144880 298284 144900
rect 298284 144880 298336 144900
rect 298336 144880 298338 144900
rect 298466 144900 298522 144936
rect 298466 144880 298468 144900
rect 298468 144880 298520 144900
rect 298520 144880 298522 144900
rect 298282 75928 298338 75984
rect 298558 75928 298614 75984
rect 298282 7520 298338 7576
rect 299570 8880 299626 8936
rect 300950 204720 301006 204776
rect 300950 204312 301006 204368
rect 301594 134156 301650 134192
rect 301594 134136 301596 134156
rect 301596 134136 301648 134156
rect 301648 134136 301650 134156
rect 302974 169668 302976 169688
rect 302976 169668 303028 169688
rect 303028 169668 303030 169688
rect 302974 169632 303030 169668
rect 304906 115912 304962 115968
rect 304262 64096 304318 64152
rect 304262 63552 304318 63608
rect 305182 241440 305238 241496
rect 305366 241440 305422 241496
rect 305182 222128 305238 222184
rect 305366 222128 305422 222184
rect 305182 202816 305238 202872
rect 305366 202816 305422 202872
rect 305182 154672 305238 154728
rect 305182 154536 305238 154592
rect 305274 145016 305330 145072
rect 305090 144880 305146 144936
rect 305090 115932 305146 115968
rect 305090 115912 305092 115932
rect 305092 115912 305144 115932
rect 305144 115912 305146 115932
rect 305182 106222 305238 106278
rect 305274 105984 305330 106040
rect 307574 134000 307630 134056
rect 307758 134000 307814 134056
rect 308034 222128 308090 222184
rect 308310 222128 308366 222184
rect 308126 202816 308182 202872
rect 308310 202816 308366 202872
rect 309046 181192 309102 181248
rect 309046 180784 309102 180840
rect 309046 169804 309048 169824
rect 309048 169804 309100 169824
rect 309100 169804 309102 169824
rect 309046 169768 309102 169804
rect 308218 153176 308274 153232
rect 308402 153176 308458 153232
rect 309046 76220 309102 76256
rect 309046 76200 309048 76220
rect 309048 76200 309100 76220
rect 309100 76200 309102 76220
rect 309414 299376 309470 299432
rect 309598 299376 309654 299432
rect 309414 280064 309470 280120
rect 309598 280064 309654 280120
rect 309322 251096 309378 251152
rect 309506 251096 309562 251152
rect 309322 211112 309378 211168
rect 309506 211112 309562 211168
rect 309506 154672 309562 154728
rect 309322 154536 309378 154592
rect 309506 133864 309562 133920
rect 309690 133864 309746 133920
rect 309414 18128 309470 18184
rect 309322 17992 309378 18048
rect 310702 241440 310758 241496
rect 310886 241440 310942 241496
rect 310702 222128 310758 222184
rect 310886 222128 310942 222184
rect 310702 183504 310758 183560
rect 310886 183504 310942 183560
rect 310702 154536 310758 154592
rect 310886 154536 310942 154592
rect 310886 46960 310942 47016
rect 310794 46688 310850 46744
rect 311806 40060 311808 40080
rect 311808 40060 311860 40080
rect 311860 40060 311862 40080
rect 311806 40024 311862 40060
rect 317326 170040 317382 170096
rect 317326 157800 317382 157856
rect 317326 157528 317382 157584
rect 317326 76220 317382 76256
rect 317326 76200 317328 76220
rect 317328 76200 317380 76220
rect 317380 76200 317382 76220
rect 317326 40160 317382 40216
rect 317326 29416 317382 29472
rect 317326 28872 317382 28928
rect 318706 76200 318762 76256
rect 318706 76064 318762 76120
rect 318706 29416 318762 29472
rect 318706 29280 318762 29336
rect 318706 16668 318708 16688
rect 318708 16668 318760 16688
rect 318760 16668 318762 16688
rect 318706 16632 318762 16668
rect 319074 114552 319130 114608
rect 319074 114416 319130 114472
rect 319626 16768 319682 16824
rect 321466 325624 321522 325680
rect 321466 316004 321468 316024
rect 321468 316004 321520 316024
rect 321520 316004 321522 316024
rect 321466 315968 321522 316004
rect 321926 335280 321982 335336
rect 322110 335280 322166 335336
rect 321650 325660 321652 325680
rect 321652 325660 321704 325680
rect 321704 325660 321706 325680
rect 321650 325624 321706 325660
rect 321650 315968 321706 316024
rect 321742 211112 321798 211168
rect 321926 211112 321982 211168
rect 321742 191800 321798 191856
rect 321926 191800 321982 191856
rect 321558 164328 321614 164384
rect 321558 164192 321614 164248
rect 321466 87352 321522 87408
rect 321466 87080 321522 87136
rect 324502 317600 324558 317656
rect 324410 317464 324466 317520
rect 324410 315968 324466 316024
rect 324686 315968 324742 316024
rect 324502 289720 324558 289776
rect 324686 289720 324742 289776
rect 324502 211112 324558 211168
rect 324686 211112 324742 211168
rect 324502 191800 324558 191856
rect 324686 191800 324742 191856
rect 324502 135360 324558 135416
rect 324502 135224 324558 135280
rect 324502 125704 324558 125760
rect 324502 125568 324558 125624
rect 326802 40160 326858 40216
rect 326986 40024 327042 40080
rect 327262 230424 327318 230480
rect 327446 230424 327502 230480
rect 328366 170060 328422 170096
rect 328366 170040 328368 170060
rect 328368 170040 328420 170060
rect 328420 170040 328422 170060
rect 327262 153176 327318 153232
rect 327446 153176 327502 153232
rect 328550 87116 328552 87136
rect 328552 87116 328604 87136
rect 328604 87116 328606 87136
rect 328550 87080 328606 87116
rect 331126 251232 331182 251288
rect 331126 251096 331182 251152
rect 331126 200096 331182 200152
rect 329930 164212 329986 164248
rect 329930 164192 329932 164212
rect 329932 164192 329984 164212
rect 329984 164192 329986 164212
rect 330114 164212 330170 164248
rect 330114 164192 330116 164212
rect 330116 164192 330168 164212
rect 330168 164192 330170 164212
rect 330114 145016 330170 145072
rect 330022 144880 330078 144936
rect 331402 289992 331458 290048
rect 331310 289720 331366 289776
rect 331402 270680 331458 270736
rect 331310 270408 331366 270464
rect 331402 200096 331458 200152
rect 331402 154556 331458 154592
rect 331402 154536 331404 154556
rect 331404 154536 331456 154556
rect 331456 154536 331458 154556
rect 331586 154536 331642 154592
rect 332690 306312 332746 306368
rect 332966 306312 333022 306368
rect 332782 219408 332838 219464
rect 333058 219408 333114 219464
rect 332690 200232 332746 200288
rect 332782 200096 332838 200152
rect 333886 134408 333942 134464
rect 333886 134000 333942 134056
rect 334070 16668 334072 16688
rect 334072 16668 334124 16688
rect 334124 16668 334126 16688
rect 334070 16632 334126 16668
rect 336738 204348 336740 204368
rect 336740 204348 336792 204368
rect 336792 204348 336794 204368
rect 336738 204312 336794 204348
rect 338118 204348 338120 204368
rect 338120 204348 338172 204368
rect 338172 204348 338174 204368
rect 338118 204312 338174 204348
rect 336646 170060 336702 170096
rect 336646 170040 336648 170060
rect 336648 170040 336700 170060
rect 336700 170040 336702 170060
rect 338026 134000 338082 134056
rect 338118 133456 338174 133512
rect 336738 110764 336794 110800
rect 336738 110744 336740 110764
rect 336740 110744 336792 110764
rect 336792 110744 336794 110764
rect 338026 87216 338082 87272
rect 337474 63572 337530 63608
rect 337474 63552 337476 63572
rect 337476 63552 337528 63572
rect 337528 63552 337530 63572
rect 336554 24792 336610 24848
rect 336738 24792 336794 24848
rect 338118 16668 338120 16688
rect 338120 16668 338172 16688
rect 338172 16668 338174 16688
rect 338118 16632 338174 16668
rect 340786 87216 340842 87272
rect 341062 40160 341118 40216
rect 341062 39752 341118 39808
rect 342442 251096 342498 251152
rect 342626 251096 342682 251152
rect 342442 231784 342498 231840
rect 342718 231784 342774 231840
rect 342718 212744 342774 212800
rect 342442 212506 342498 212562
rect 342718 191800 342774 191856
rect 342902 191800 342958 191856
rect 343546 181328 343602 181384
rect 343546 181192 343602 181248
rect 342534 172508 342590 172544
rect 342534 172488 342536 172508
rect 342536 172488 342588 172508
rect 342588 172488 342590 172508
rect 342902 172488 342958 172544
rect 342350 154536 342406 154592
rect 342534 154536 342590 154592
rect 342258 4800 342314 4856
rect 344926 123256 344982 123312
rect 344926 122848 344982 122904
rect 344926 63572 344982 63608
rect 344926 63552 344928 63572
rect 344928 63552 344980 63572
rect 344980 63552 344982 63572
rect 345938 123276 345994 123312
rect 345938 123256 345940 123276
rect 345940 123256 345992 123276
rect 345992 123256 345994 123276
rect 346214 110472 346270 110528
rect 346214 63588 346216 63608
rect 346216 63588 346268 63608
rect 346268 63588 346270 63608
rect 346214 63552 346270 63588
rect 347686 267688 347742 267744
rect 347686 258032 347742 258088
rect 346582 241440 346638 241496
rect 346766 241440 346822 241496
rect 346582 222128 346638 222184
rect 346766 222128 346822 222184
rect 346582 202816 346638 202872
rect 346766 202816 346822 202872
rect 346490 63824 346546 63880
rect 347686 16804 347688 16824
rect 347688 16804 347740 16824
rect 347740 16804 347742 16824
rect 347686 16768 347742 16804
rect 347962 333920 348018 333976
rect 348238 333920 348294 333976
rect 347870 267724 347872 267744
rect 347872 267724 347924 267744
rect 347924 267724 347926 267744
rect 347870 267688 347926 267724
rect 348054 258032 348110 258088
rect 347962 134000 348018 134056
rect 347962 133864 348018 133920
rect 349802 40432 349858 40488
rect 349802 40160 349858 40216
rect 351826 269048 351882 269104
rect 351826 240080 351882 240136
rect 351826 230424 351882 230480
rect 351826 201456 351882 201512
rect 351826 104760 351882 104816
rect 350998 29416 351054 29472
rect 350998 29144 351054 29200
rect 352102 325624 352158 325680
rect 352286 325624 352342 325680
rect 352102 316004 352104 316024
rect 352104 316004 352156 316024
rect 352156 316004 352158 316024
rect 352102 315968 352158 316004
rect 352286 316004 352288 316024
rect 352288 316004 352340 316024
rect 352340 316004 352342 316024
rect 352286 315968 352342 316004
rect 352102 287000 352158 287056
rect 352286 287000 352342 287056
rect 352102 269048 352158 269104
rect 352010 240080 352066 240136
rect 352102 230424 352158 230480
rect 352102 201476 352158 201512
rect 352102 201456 352104 201476
rect 352104 201456 352156 201476
rect 352156 201456 352158 201476
rect 352102 125704 352158 125760
rect 352010 125568 352066 125624
rect 352010 104760 352066 104816
rect 353482 134000 353538 134056
rect 353482 133884 353538 133920
rect 353482 133864 353484 133884
rect 353484 133864 353536 133884
rect 353536 133864 353538 133884
rect 354586 123120 354642 123176
rect 353482 114416 353538 114472
rect 353574 114280 353630 114336
rect 354586 87216 354642 87272
rect 353390 66272 353446 66328
rect 353666 66000 353722 66056
rect 355506 63844 355562 63880
rect 355506 63824 355508 63844
rect 355508 63824 355560 63844
rect 355560 63824 355562 63844
rect 355966 17176 356022 17232
rect 356518 288360 356574 288416
rect 356702 288360 356758 288416
rect 356426 248396 356482 248432
rect 356426 248376 356428 248396
rect 356428 248376 356480 248396
rect 356480 248376 356482 248396
rect 356610 248376 356666 248432
rect 356334 238720 356390 238776
rect 356518 238720 356574 238776
rect 356426 212508 356428 212528
rect 356428 212508 356480 212528
rect 356480 212508 356482 212528
rect 356426 212472 356482 212508
rect 356610 212472 356666 212528
rect 356426 144880 356482 144936
rect 356426 144744 356482 144800
rect 356426 134000 356482 134056
rect 356426 133884 356482 133920
rect 356426 133864 356428 133884
rect 356428 133864 356480 133884
rect 356480 133864 356482 133884
rect 356426 94016 356482 94072
rect 356426 93880 356482 93936
rect 356334 24792 356390 24848
rect 356518 24792 356574 24848
rect 356150 3304 356206 3360
rect 357530 315968 357586 316024
rect 357714 315968 357770 316024
rect 357530 296656 357586 296712
rect 357806 296656 357862 296712
rect 357530 144900 357586 144936
rect 357530 144880 357532 144900
rect 357532 144880 357584 144900
rect 357584 144880 357586 144900
rect 357714 144900 357770 144936
rect 357714 144880 357716 144900
rect 357716 144880 357768 144900
rect 357768 144880 357770 144900
rect 357622 125704 357678 125760
rect 357622 125568 357678 125624
rect 357530 86944 357586 87000
rect 357714 86944 357770 87000
rect 359002 270680 359058 270736
rect 359186 270408 359242 270464
rect 359002 249736 359058 249792
rect 359278 249736 359334 249792
rect 359094 229064 359150 229120
rect 359278 229064 359334 229120
rect 359186 200232 359242 200288
rect 359094 198736 359150 198792
rect 359002 144900 359058 144936
rect 359002 144880 359004 144900
rect 359004 144880 359056 144900
rect 359056 144880 359058 144900
rect 359186 144900 359242 144936
rect 359186 144880 359188 144900
rect 359188 144880 359240 144900
rect 359240 144880 359242 144900
rect 359094 124208 359150 124264
rect 359186 114416 359242 114472
rect 360382 63552 360438 63608
rect 364522 270680 364578 270736
rect 364614 270408 364670 270464
rect 365718 191800 365774 191856
rect 365902 191800 365958 191856
rect 364614 190440 364670 190496
rect 364798 190440 364854 190496
rect 365718 172488 365774 172544
rect 365902 172488 365958 172544
rect 365718 169940 365720 169960
rect 365720 169940 365772 169960
rect 365772 169940 365774 169960
rect 365718 169904 365774 169940
rect 365626 87236 365682 87272
rect 365626 87216 365628 87236
rect 365628 87216 365680 87236
rect 365680 87216 365682 87236
rect 368294 169940 368296 169960
rect 368296 169940 368348 169960
rect 368348 169940 368350 169960
rect 368294 169904 368350 169940
rect 367374 135360 367430 135416
rect 367374 135244 367430 135280
rect 367374 135224 367376 135244
rect 367376 135224 367428 135244
rect 367428 135224 367430 135244
rect 367374 125568 367430 125624
rect 367558 125568 367614 125624
rect 367374 55392 367430 55448
rect 367282 55256 367338 55312
rect 367374 45600 367430 45656
rect 367466 45464 367522 45520
rect 369950 267688 370006 267744
rect 370134 267688 370190 267744
rect 369950 258032 370006 258088
rect 370134 258032 370190 258088
rect 371146 180920 371202 180976
rect 371146 180648 371202 180704
rect 370042 135224 370098 135280
rect 370226 135224 370282 135280
rect 372618 181212 372674 181248
rect 372618 181192 372620 181212
rect 372620 181192 372672 181212
rect 372672 181192 372674 181212
rect 373906 87080 373962 87136
rect 373906 29280 373962 29336
rect 373906 28872 373962 28928
rect 375194 204448 375250 204504
rect 375470 267688 375526 267744
rect 375654 267688 375710 267744
rect 375470 258032 375526 258088
rect 375654 258032 375710 258088
rect 375654 211112 375710 211168
rect 375838 211112 375894 211168
rect 375470 157528 375526 157584
rect 375470 157256 375526 157312
rect 376942 164212 376998 164248
rect 376942 164192 376944 164212
rect 376944 164192 376996 164212
rect 376996 164192 376998 164212
rect 377126 164192 377182 164248
rect 379334 170040 379390 170096
rect 379518 170040 379574 170096
rect 380806 220768 380862 220824
rect 380806 211112 380862 211168
rect 381174 318960 381230 319016
rect 381082 318824 381138 318880
rect 381082 220768 381138 220824
rect 380990 211112 381046 211168
rect 382278 241440 382334 241496
rect 382462 241440 382518 241496
rect 382278 222128 382334 222184
rect 382462 222128 382518 222184
rect 382278 202816 382334 202872
rect 382462 202816 382518 202872
rect 382278 182144 382334 182200
rect 382462 182144 382518 182200
rect 382186 180920 382242 180976
rect 383658 134036 383660 134056
rect 383660 134036 383712 134056
rect 383712 134036 383714 134056
rect 383658 134000 383714 134036
rect 383566 63688 383622 63744
rect 383566 63416 383622 63472
rect 383566 40160 383622 40216
rect 383566 40024 383622 40080
rect 383566 29552 383622 29608
rect 383566 29144 383622 29200
rect 384946 204448 385002 204504
rect 384946 87216 385002 87272
rect 384946 86808 385002 86864
rect 385222 134136 385278 134192
rect 386602 231820 386604 231840
rect 386604 231820 386656 231840
rect 386656 231820 386658 231840
rect 386602 231784 386658 231820
rect 386878 231820 386880 231840
rect 386880 231820 386932 231840
rect 386932 231820 386934 231840
rect 386878 231784 386934 231820
rect 386602 154556 386658 154592
rect 386602 154536 386604 154556
rect 386604 154536 386656 154556
rect 386656 154536 386658 154556
rect 386786 154556 386842 154592
rect 386786 154536 386788 154556
rect 386788 154536 386840 154556
rect 386840 154536 386842 154556
rect 386786 135360 386842 135416
rect 386602 135224 386658 135280
rect 388074 96600 388130 96656
rect 387982 96464 388038 96520
rect 392122 278704 392178 278760
rect 393226 278704 393282 278760
rect 393410 278704 393466 278760
rect 392214 278568 392270 278624
rect 393226 269084 393228 269104
rect 393228 269084 393280 269104
rect 393280 269084 393282 269104
rect 393226 269048 393282 269084
rect 393410 269084 393412 269104
rect 393412 269084 393464 269104
rect 393464 269084 393466 269104
rect 393410 269048 393466 269084
rect 392950 249736 393006 249792
rect 393134 249736 393190 249792
rect 392122 241476 392124 241496
rect 392124 241476 392176 241496
rect 392176 241476 392178 241496
rect 392122 241440 392178 241476
rect 392306 241440 392362 241496
rect 392306 240080 392362 240136
rect 392490 240080 392546 240136
rect 392122 222164 392124 222184
rect 392124 222164 392176 222184
rect 392176 222164 392178 222184
rect 392122 222128 392178 222164
rect 392214 221992 392270 222048
rect 392122 154672 392178 154728
rect 392122 154556 392178 154592
rect 392122 154536 392124 154556
rect 392124 154536 392176 154556
rect 392176 154536 392178 154556
rect 392214 138216 392270 138272
rect 392122 135224 392178 135280
rect 393226 125704 393282 125760
rect 393226 125568 393282 125624
rect 392030 96600 392086 96656
rect 392214 96600 392270 96656
rect 393318 63688 393374 63744
rect 395894 29144 395950 29200
rect 396078 29144 396134 29200
rect 397734 115912 397790 115968
rect 397918 115912 397974 115968
rect 398746 76236 398748 76256
rect 398748 76236 398800 76256
rect 398800 76236 398802 76256
rect 398746 76200 398802 76236
rect 400402 231784 400458 231840
rect 400586 231784 400642 231840
rect 400310 222128 400366 222184
rect 400494 222164 400496 222184
rect 400496 222164 400548 222184
rect 400548 222164 400550 222184
rect 400494 222128 400550 222164
rect 402886 134272 402942 134328
rect 402886 133864 402942 133920
rect 402978 40332 402980 40352
rect 402980 40332 403032 40352
rect 403032 40332 403034 40352
rect 402978 40296 403034 40332
rect 405738 157700 405740 157720
rect 405740 157700 405792 157720
rect 405792 157700 405794 157720
rect 405738 157664 405794 157700
rect 405646 134272 405702 134328
rect 405738 134136 405794 134192
rect 405646 76236 405648 76256
rect 405648 76236 405700 76256
rect 405700 76236 405702 76256
rect 405646 76200 405702 76236
rect 405646 63844 405702 63880
rect 405646 63824 405648 63844
rect 405648 63824 405700 63844
rect 405700 63824 405702 63844
rect 405738 16904 405794 16960
rect 405738 16768 405794 16824
rect 407486 249736 407542 249792
rect 407670 249736 407726 249792
rect 408406 154536 408462 154592
rect 408774 248376 408830 248432
rect 408958 248376 409014 248432
rect 408682 202816 408738 202872
rect 408958 202816 409014 202872
rect 408682 183504 408738 183560
rect 408958 183504 409014 183560
rect 408682 154536 408738 154592
rect 408866 135224 408922 135280
rect 409050 135224 409106 135280
rect 408866 125704 408922 125760
rect 408682 125568 408738 125624
rect 408682 27512 408738 27568
rect 408774 27376 408830 27432
rect 408314 3612 408316 3632
rect 408316 3612 408368 3632
rect 408368 3612 408370 3632
rect 408314 3576 408370 3612
rect 408590 3612 408592 3632
rect 408592 3612 408644 3632
rect 408644 3612 408646 3632
rect 408590 3576 408646 3612
rect 410522 3304 410578 3360
rect 412454 40432 412510 40488
rect 413926 40432 413982 40488
rect 413926 40160 413982 40216
rect 415306 157700 415308 157720
rect 415308 157700 415360 157720
rect 415360 157700 415362 157720
rect 415306 157664 415362 157700
rect 415398 87100 415454 87136
rect 415398 87080 415400 87100
rect 415400 87080 415452 87100
rect 415452 87080 415454 87100
rect 416870 241440 416926 241496
rect 417146 241440 417202 241496
rect 416870 222128 416926 222184
rect 417146 222128 417202 222184
rect 416870 202816 416926 202872
rect 417146 202816 417202 202872
rect 416778 135224 416834 135280
rect 416962 135224 417018 135280
rect 416778 115912 416834 115968
rect 416962 115912 417018 115968
rect 416778 96600 416834 96656
rect 416962 96600 417018 96656
rect 418066 204448 418122 204504
rect 418066 204040 418122 204096
rect 418066 169904 418122 169960
rect 418066 169496 418122 169552
rect 417882 134272 417938 134328
rect 418250 134136 418306 134192
rect 418066 110608 418122 110664
rect 418066 110200 418122 110256
rect 418066 76200 418122 76256
rect 418158 76064 418214 76120
rect 418066 63824 418122 63880
rect 418158 63688 418214 63744
rect 418066 16904 418122 16960
rect 418250 16904 418306 16960
rect 422390 183504 422446 183560
rect 422666 183504 422722 183560
rect 424874 86944 424930 87000
rect 425058 204348 425060 204368
rect 425060 204348 425112 204368
rect 425112 204348 425114 204368
rect 425058 204312 425114 204348
rect 425058 180820 425060 180840
rect 425060 180820 425112 180840
rect 425112 180820 425114 180840
rect 425058 180784 425114 180820
rect 425058 169804 425060 169824
rect 425060 169804 425112 169824
rect 425112 169804 425114 169824
rect 425058 169768 425114 169804
rect 425058 122884 425060 122904
rect 425060 122884 425112 122904
rect 425112 122884 425114 122904
rect 425058 122848 425114 122884
rect 425058 110508 425060 110528
rect 425060 110508 425112 110528
rect 425112 110508 425114 110528
rect 425058 110472 425114 110508
rect 425058 86980 425060 87000
rect 425060 86980 425112 87000
rect 425112 86980 425114 87000
rect 425058 86944 425114 86980
rect 427726 135224 427782 135280
rect 427910 135224 427966 135280
rect 434166 328616 434222 328672
rect 433706 328480 433762 328536
rect 433430 241440 433486 241496
rect 433614 241440 433670 241496
rect 433430 222128 433486 222184
rect 433614 222128 433670 222184
rect 434534 204584 434590 204640
rect 434534 181056 434590 181112
rect 434534 170040 434590 170096
rect 434534 123120 434590 123176
rect 434534 110744 434590 110800
rect 434534 87216 434590 87272
rect 451370 335280 451426 335336
rect 451830 335280 451886 335336
rect 451554 325660 451556 325680
rect 451556 325660 451608 325680
rect 451608 325660 451610 325680
rect 451554 325624 451610 325660
rect 451738 325624 451794 325680
rect 451278 288360 451334 288416
rect 451462 288360 451518 288416
rect 451278 222164 451280 222184
rect 451280 222164 451332 222184
rect 451332 222164 451334 222184
rect 451278 222128 451334 222164
rect 451738 221992 451794 222048
rect 451830 162832 451886 162888
rect 451646 99456 451702 99512
rect 451646 96600 451702 96656
rect 452014 162832 452070 162888
rect 454038 169940 454040 169960
rect 454040 169940 454092 169960
rect 454092 169940 454094 169960
rect 454038 169904 454094 169940
rect 454038 123020 454040 123040
rect 454040 123020 454092 123040
rect 454092 123020 454094 123040
rect 454038 122984 454094 123020
rect 456706 157528 456762 157584
rect 456890 157528 456946 157584
rect 456706 134000 456762 134056
rect 456890 134000 456946 134056
rect 456706 76064 456762 76120
rect 456890 76064 456946 76120
rect 456706 63688 456762 63744
rect 456890 63688 456946 63744
rect 456706 40160 456762 40216
rect 456890 40160 456946 40216
rect 456706 16768 456762 16824
rect 456890 16768 456946 16824
rect 458178 169940 458180 169960
rect 458180 169940 458232 169960
rect 458232 169940 458234 169960
rect 458178 169904 458234 169940
rect 458178 123020 458180 123040
rect 458180 123020 458232 123040
rect 458232 123020 458234 123040
rect 458178 122984 458234 123020
rect 466274 29008 466330 29064
rect 472070 241440 472126 241496
rect 472346 241440 472402 241496
rect 472070 222128 472126 222184
rect 472346 222128 472402 222184
rect 472070 202816 472126 202872
rect 472346 202816 472402 202872
rect 472070 183504 472126 183560
rect 472346 183504 472402 183560
rect 472162 154536 472218 154592
rect 472346 154536 472402 154592
rect 471978 135224 472034 135280
rect 472162 135224 472218 135280
rect 471978 115912 472034 115968
rect 472162 115912 472218 115968
rect 471978 96600 472034 96656
rect 472162 96600 472218 96656
rect 473266 29280 473322 29336
rect 475934 180940 475990 180976
rect 475934 180920 475936 180940
rect 475936 180920 475988 180940
rect 475988 180920 475990 180940
rect 475934 169924 475990 169960
rect 475934 169904 475936 169924
rect 475936 169904 475988 169924
rect 475988 169904 475990 169924
rect 475934 123004 475990 123040
rect 475934 122984 475936 123004
rect 475936 122984 475988 123004
rect 475988 122984 475990 123004
rect 475934 87100 475990 87136
rect 475934 87080 475936 87100
rect 475936 87080 475988 87100
rect 475988 87080 475990 87100
rect 475934 76084 475990 76120
rect 475934 76064 475936 76084
rect 475936 76064 475988 76084
rect 475988 76064 475990 76084
rect 476118 180940 476174 180976
rect 476118 180920 476120 180940
rect 476120 180920 476172 180940
rect 476172 180920 476174 180940
rect 476118 169924 476174 169960
rect 476118 169904 476120 169924
rect 476120 169904 476172 169924
rect 476172 169904 476174 169924
rect 476118 87100 476174 87136
rect 476118 87080 476120 87100
rect 476120 87080 476172 87100
rect 476172 87080 476174 87100
rect 478142 123004 478198 123040
rect 478142 122984 478144 123004
rect 478144 122984 478196 123004
rect 478196 122984 478198 123004
rect 478142 76084 478198 76120
rect 478142 76064 478144 76084
rect 478144 76064 478196 76084
rect 478196 76064 478198 76084
rect 480166 278704 480222 278760
rect 480350 278704 480406 278760
rect 480166 259392 480222 259448
rect 480350 259392 480406 259448
rect 480350 241712 480406 241768
rect 480350 241576 480406 241632
rect 480166 240080 480222 240136
rect 480350 240080 480406 240136
rect 480166 220768 480222 220824
rect 480350 220768 480406 220824
rect 480166 211112 480222 211168
rect 480350 211112 480406 211168
rect 480350 164212 480406 164248
rect 480350 164192 480352 164212
rect 480352 164192 480404 164212
rect 480404 164192 480406 164212
rect 480534 164192 480590 164248
rect 480258 115912 480314 115968
rect 480442 115912 480498 115968
rect 514574 204448 514630 204504
rect 514574 204040 514630 204096
rect 514574 180920 514630 180976
rect 514574 180512 514630 180568
rect 514574 169940 514576 169960
rect 514576 169940 514628 169960
rect 514628 169940 514630 169960
rect 514574 169904 514630 169940
rect 514574 157528 514630 157584
rect 514574 157120 514630 157176
rect 514574 134000 514630 134056
rect 514574 133592 514630 133648
rect 514574 123020 514576 123040
rect 514576 123020 514628 123040
rect 514628 123020 514630 123040
rect 514574 122984 514630 123020
rect 514574 110608 514630 110664
rect 514574 110200 514630 110256
rect 514574 76100 514576 76120
rect 514576 76100 514628 76120
rect 514628 76100 514630 76120
rect 514574 76064 514630 76100
rect 514574 63688 514630 63744
rect 514574 63280 514630 63336
rect 514574 40160 514630 40216
rect 514574 39752 514630 39808
rect 514574 16788 514630 16824
rect 514574 16768 514576 16788
rect 514576 16768 514628 16788
rect 514628 16768 514630 16788
rect 516046 16788 516102 16824
rect 516046 16768 516048 16788
rect 516048 16768 516100 16788
rect 516100 16768 516102 16788
rect 516874 169940 516876 169960
rect 516876 169940 516928 169960
rect 516928 169940 516930 169960
rect 516874 169904 516930 169940
rect 516874 123020 516876 123040
rect 516876 123020 516928 123040
rect 516928 123020 516930 123040
rect 516874 122984 516930 123020
rect 516874 76100 516876 76120
rect 516876 76100 516928 76120
rect 516928 76100 516930 76120
rect 516874 76064 516930 76100
rect 521658 204348 521660 204368
rect 521660 204348 521712 204368
rect 521712 204348 521714 204368
rect 521658 204312 521714 204348
rect 521658 180820 521660 180840
rect 521660 180820 521712 180840
rect 521712 180820 521714 180840
rect 521658 180784 521714 180820
rect 521658 157428 521660 157448
rect 521660 157428 521712 157448
rect 521712 157428 521714 157448
rect 521658 157392 521714 157428
rect 521658 133900 521660 133920
rect 521660 133900 521712 133920
rect 521712 133900 521714 133920
rect 521658 133864 521714 133900
rect 521658 110508 521660 110528
rect 521660 110508 521712 110528
rect 521712 110508 521714 110528
rect 521658 110472 521714 110508
rect 521658 63588 521660 63608
rect 521660 63588 521712 63608
rect 521712 63588 521714 63608
rect 521658 63552 521714 63588
rect 521658 40060 521660 40080
rect 521660 40060 521712 40080
rect 521712 40060 521714 40080
rect 521658 40024 521714 40060
rect 521658 29044 521660 29064
rect 521660 29044 521712 29064
rect 521712 29044 521714 29064
rect 521658 29008 521714 29044
rect 523222 337728 523278 337784
rect 524234 169804 524236 169824
rect 524236 169804 524288 169824
rect 524288 169804 524290 169824
rect 524234 169768 524290 169804
rect 524234 122884 524236 122904
rect 524236 122884 524288 122904
rect 524288 122884 524290 122904
rect 524234 122848 524290 122884
rect 524234 75964 524236 75984
rect 524236 75964 524288 75984
rect 524288 75964 524290 75984
rect 524234 75928 524290 75964
rect 524234 16668 524236 16688
rect 524236 16668 524288 16688
rect 524288 16668 524290 16688
rect 524234 16632 524290 16668
rect 525062 86944 525118 87000
rect 525062 86672 525118 86728
rect 528190 337320 528246 337376
rect 529478 337728 529534 337784
rect 526442 204448 526498 204504
rect 526442 180920 526498 180976
rect 526442 169904 526498 169960
rect 526442 157528 526498 157584
rect 526442 134000 526498 134056
rect 526442 122984 526498 123040
rect 526442 110608 526498 110664
rect 526442 76064 526498 76120
rect 526442 63688 526498 63744
rect 526442 40160 526498 40216
rect 525890 29144 525946 29200
rect 526442 16768 526498 16824
rect 525706 3304 525762 3360
rect 530674 637880 530730 637936
rect 530950 638288 531006 638344
rect 579802 639376 579858 639432
rect 580078 627680 580134 627736
rect 580078 604152 580134 604208
rect 580078 592456 580134 592512
rect 580078 580760 580134 580816
rect 580078 557232 580134 557288
rect 580078 545536 580134 545592
rect 580078 510312 580134 510368
rect 580078 498616 580134 498672
rect 580170 486784 580226 486840
rect 579802 463392 579858 463448
rect 580170 439864 580226 439920
rect 580170 416472 580226 416528
rect 579618 392944 579674 393000
rect 580170 346024 580226 346080
rect 536102 87352 536158 87408
rect 536102 86944 536158 87000
rect 540886 204720 540942 204776
rect 540886 204312 540942 204368
rect 540886 181192 540942 181248
rect 540886 180784 540942 180840
rect 540886 170176 540942 170232
rect 540886 169768 540942 169824
rect 540886 157800 540942 157856
rect 540886 157392 540942 157448
rect 540886 134272 540942 134328
rect 540886 133864 540942 133920
rect 540886 123256 540942 123312
rect 540886 122848 540942 122904
rect 540886 110880 540942 110936
rect 540886 110472 540942 110528
rect 540886 76336 540942 76392
rect 540886 75928 540942 75984
rect 540886 63960 540942 64016
rect 540886 63552 540942 63608
rect 540886 40432 540942 40488
rect 540886 40024 540942 40080
rect 540794 29416 540850 29472
rect 540886 29008 540942 29064
rect 540886 17040 540942 17096
rect 540886 16632 540942 16688
rect 545670 274932 545672 274952
rect 545672 274932 545724 274952
rect 545724 274932 545726 274952
rect 545670 274896 545726 274932
rect 550546 274932 550548 274952
rect 550548 274932 550600 274952
rect 550600 274932 550602 274952
rect 550546 274896 550602 274932
rect 553306 180956 553308 180976
rect 553308 180956 553360 180976
rect 553360 180956 553362 180976
rect 553306 180920 553362 180956
rect 554962 180956 554964 180976
rect 554964 180956 555016 180976
rect 555016 180956 555018 180976
rect 554962 180920 555018 180956
rect 560206 204584 560262 204640
rect 560206 204176 560262 204232
rect 560206 170040 560262 170096
rect 560206 169632 560262 169688
rect 560206 157664 560262 157720
rect 560206 157256 560262 157312
rect 560206 134136 560262 134192
rect 560206 133728 560262 133784
rect 560206 123120 560262 123176
rect 560206 122712 560262 122768
rect 560206 110744 560262 110800
rect 560206 110336 560262 110392
rect 560206 87488 560262 87544
rect 560206 87216 560262 87272
rect 560206 76200 560262 76256
rect 560206 75792 560262 75848
rect 560206 63824 560262 63880
rect 560206 63416 560262 63472
rect 560206 40296 560262 40352
rect 560206 39888 560262 39944
rect 560206 29552 560262 29608
rect 560206 29280 560262 29336
rect 560206 16904 560262 16960
rect 560206 16496 560262 16552
rect 563058 274896 563114 274952
rect 563058 274488 563114 274544
rect 565082 337320 565138 337376
rect 572626 274760 572682 274816
rect 572718 274624 572774 274680
rect 572626 204448 572682 204504
rect 572718 204312 572774 204368
rect 572626 169904 572682 169960
rect 572718 169768 572774 169824
rect 572626 157528 572682 157584
rect 572718 157392 572774 157448
rect 572626 134000 572682 134056
rect 572718 133864 572774 133920
rect 572626 122984 572682 123040
rect 572718 122848 572774 122904
rect 572626 110608 572682 110664
rect 572718 110472 572774 110528
rect 572626 87100 572682 87136
rect 572626 87080 572628 87100
rect 572628 87080 572680 87100
rect 572680 87080 572682 87100
rect 572626 76064 572682 76120
rect 572718 75928 572774 75984
rect 572626 63688 572682 63744
rect 572718 63552 572774 63608
rect 572626 40160 572682 40216
rect 572718 40024 572774 40080
rect 572626 29180 572628 29200
rect 572628 29180 572680 29200
rect 572680 29180 572682 29200
rect 572626 29144 572682 29180
rect 572626 16768 572682 16824
rect 572718 16632 572774 16688
rect 579618 322632 579674 322688
rect 579710 299104 579766 299160
rect 580906 451696 580962 451752
rect 580814 404776 580870 404832
rect 580722 357856 580778 357912
rect 580630 310800 580686 310856
rect 580538 263880 580594 263936
rect 580446 252184 580502 252240
rect 580354 228792 580410 228848
rect 580262 216960 580318 217016
rect 576766 87100 576822 87136
rect 576766 87080 576768 87100
rect 576768 87080 576820 87100
rect 576820 87080 576822 87100
rect 576766 29180 576768 29200
rect 576768 29180 576820 29200
rect 576820 29180 576822 29200
rect 576766 29144 576822 29180
rect 575018 3304 575074 3360
<< metal3 >>
rect 8109 700362 8175 700365
rect 414013 700362 414079 700365
rect 8109 700360 414079 700362
rect 8109 700304 8114 700360
rect 8170 700304 414018 700360
rect 414074 700304 414079 700360
rect 8109 700302 414079 700304
rect 8109 700299 8175 700302
rect 414013 700299 414079 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 494881 686082 494947 686085
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 494237 685883 494303 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 3509 642970 3575 642973
rect 517789 642970 517855 642973
rect 3509 642968 517855 642970
rect 3509 642912 3514 642968
rect 3570 642912 517794 642968
rect 517850 642912 517855 642968
rect 3509 642910 517855 642912
rect 3509 642907 3575 642910
rect 517789 642907 517855 642910
rect 317781 642834 317847 642837
rect 527398 642834 527404 642836
rect 317781 642832 527404 642834
rect 317781 642776 317786 642832
rect 317842 642776 527404 642832
rect 317781 642774 527404 642776
rect 317781 642771 317847 642774
rect 527398 642772 527404 642774
rect 527468 642772 527474 642836
rect 258942 642636 258948 642700
rect 259012 642698 259018 642700
rect 473077 642698 473143 642701
rect 259012 642696 473143 642698
rect 259012 642640 473082 642696
rect 473138 642640 473143 642696
rect 259012 642638 473143 642640
rect 259012 642636 259018 642638
rect 473077 642635 473143 642638
rect 261886 642500 261892 642564
rect 261956 642562 261962 642564
rect 478321 642562 478387 642565
rect 261956 642560 478387 642562
rect 261956 642504 478326 642560
rect 478382 642504 478387 642560
rect 261956 642502 478387 642504
rect 261956 642500 261962 642502
rect 478321 642499 478387 642502
rect 261702 642364 261708 642428
rect 261772 642426 261778 642428
rect 483657 642426 483723 642429
rect 261772 642424 483723 642426
rect 261772 642368 483662 642424
rect 483718 642368 483723 642424
rect 261772 642366 483723 642368
rect 261772 642364 261778 642366
rect 483657 642363 483723 642366
rect 261518 642228 261524 642292
rect 261588 642290 261594 642292
rect 491477 642290 491543 642293
rect 261588 642288 491543 642290
rect 261588 642232 491482 642288
rect 491538 642232 491543 642288
rect 261588 642230 491543 642232
rect 261588 642228 261594 642230
rect 491477 642227 491543 642230
rect 258758 642092 258764 642156
rect 258828 642154 258834 642156
rect 494145 642154 494211 642157
rect 258828 642152 494211 642154
rect 258828 642096 494150 642152
rect 494206 642096 494211 642152
rect 258828 642094 494211 642096
rect 258828 642092 258834 642094
rect 494145 642091 494211 642094
rect 288893 642018 288959 642021
rect 527950 642018 527956 642020
rect 288893 642016 527956 642018
rect 288893 641960 288898 642016
rect 288954 641960 527956 642016
rect 288893 641958 527956 641960
rect 288893 641955 288959 641958
rect 527950 641956 527956 641958
rect 528020 641956 528026 642020
rect 258574 641820 258580 641884
rect 258644 641882 258650 641884
rect 504633 641882 504699 641885
rect 258644 641880 504699 641882
rect 258644 641824 504638 641880
rect 504694 641824 504699 641880
rect 258644 641822 504699 641824
rect 258644 641820 258650 641822
rect 504633 641819 504699 641822
rect 398097 639706 398163 639709
rect 402830 639706 402836 639708
rect 398097 639704 402836 639706
rect 398097 639648 398102 639704
rect 398158 639648 402836 639704
rect 398097 639646 402836 639648
rect 398097 639643 398163 639646
rect 402830 639644 402836 639646
rect 402900 639644 402906 639708
rect 420177 639706 420243 639709
rect 415350 639704 420243 639706
rect 415350 639648 420182 639704
rect 420238 639648 420243 639704
rect 415350 639646 420243 639648
rect 384982 639372 384988 639436
rect 385052 639434 385058 639436
rect 398097 639434 398163 639437
rect 385052 639432 398163 639434
rect 385052 639376 398102 639432
rect 398158 639376 398163 639432
rect 385052 639374 398163 639376
rect 385052 639372 385058 639374
rect 398097 639371 398163 639374
rect 231393 639298 231459 639301
rect 231710 639298 231716 639300
rect 231393 639296 231716 639298
rect -960 639012 480 639252
rect 231393 639240 231398 639296
rect 231454 639240 231716 639296
rect 231393 639238 231716 639240
rect 231393 639235 231459 639238
rect 231710 639236 231716 639238
rect 231780 639236 231786 639300
rect 233969 639298 234035 639301
rect 234470 639298 234476 639300
rect 233969 639296 234476 639298
rect 233969 639240 233974 639296
rect 234030 639240 234476 639296
rect 233969 639238 234476 639240
rect 233969 639235 234035 639238
rect 234470 639236 234476 639238
rect 234540 639236 234546 639300
rect 236545 639298 236611 639301
rect 237230 639298 237236 639300
rect 236545 639296 237236 639298
rect 236545 639240 236550 639296
rect 236606 639240 237236 639296
rect 236545 639238 237236 639240
rect 236545 639235 236611 639238
rect 237230 639236 237236 639238
rect 237300 639236 237306 639300
rect 239121 639298 239187 639301
rect 239990 639298 239996 639300
rect 239121 639296 239996 639298
rect 239121 639240 239126 639296
rect 239182 639240 239996 639296
rect 239121 639238 239996 639240
rect 239121 639235 239187 639238
rect 239990 639236 239996 639238
rect 240060 639236 240066 639300
rect 241881 639298 241947 639301
rect 243997 639300 244063 639301
rect 242750 639298 242756 639300
rect 241881 639296 242756 639298
rect 241881 639240 241886 639296
rect 241942 639240 242756 639296
rect 241881 639238 242756 639240
rect 241881 639235 241947 639238
rect 242750 639236 242756 639238
rect 242820 639236 242826 639300
rect 243997 639296 244044 639300
rect 244108 639298 244114 639300
rect 246941 639298 247007 639301
rect 247534 639298 247540 639300
rect 243997 639240 244002 639296
rect 243997 639236 244044 639240
rect 244108 639238 244154 639298
rect 246941 639296 247540 639298
rect 246941 639240 246946 639296
rect 247002 639240 247540 639296
rect 246941 639238 247540 639240
rect 244108 639236 244114 639238
rect 243997 639235 244063 639236
rect 246941 639235 247007 639238
rect 247534 639236 247540 639238
rect 247604 639236 247610 639300
rect 249006 639236 249012 639300
rect 249076 639298 249082 639300
rect 249149 639298 249215 639301
rect 249076 639296 249215 639298
rect 249076 639240 249154 639296
rect 249210 639240 249215 639296
rect 249076 639238 249215 639240
rect 249076 639236 249082 639238
rect 249149 639235 249215 639238
rect 252277 639300 252343 639301
rect 252277 639296 252324 639300
rect 252388 639298 252394 639300
rect 254945 639298 255011 639301
rect 255078 639298 255084 639300
rect 252277 639240 252282 639296
rect 252277 639236 252324 639240
rect 252388 639238 252434 639298
rect 254945 639296 255084 639298
rect 254945 639240 254950 639296
rect 255006 639240 255084 639296
rect 254945 639238 255084 639240
rect 252388 639236 252394 639238
rect 252277 639235 252343 639236
rect 254945 639235 255011 639238
rect 255078 639236 255084 639238
rect 255148 639236 255154 639300
rect 257705 639298 257771 639301
rect 257838 639298 257844 639300
rect 257705 639296 257844 639298
rect 257705 639240 257710 639296
rect 257766 639240 257844 639296
rect 257705 639238 257844 639240
rect 257705 639235 257771 639238
rect 257838 639236 257844 639238
rect 257908 639236 257914 639300
rect 260281 639298 260347 639301
rect 261334 639298 261340 639300
rect 260281 639296 261340 639298
rect 260281 639240 260286 639296
rect 260342 639240 261340 639296
rect 260281 639238 261340 639240
rect 260281 639235 260347 639238
rect 261334 639236 261340 639238
rect 261404 639236 261410 639300
rect 262857 639298 262923 639301
rect 273161 639300 273227 639301
rect 263358 639298 263364 639300
rect 262857 639296 263364 639298
rect 262857 639240 262862 639296
rect 262918 639240 263364 639296
rect 262857 639238 263364 639240
rect 262857 639235 262923 639238
rect 263358 639236 263364 639238
rect 263428 639236 263434 639300
rect 273110 639298 273116 639300
rect 273070 639238 273116 639298
rect 273180 639296 273227 639300
rect 273222 639240 273227 639296
rect 273110 639236 273116 639238
rect 273180 639236 273227 639240
rect 273161 639235 273227 639236
rect 281165 639300 281231 639301
rect 281165 639296 281212 639300
rect 281276 639298 281282 639300
rect 304901 639298 304967 639301
rect 307518 639298 307524 639300
rect 281165 639240 281170 639296
rect 281165 639236 281212 639240
rect 281276 639238 281322 639298
rect 304901 639296 307524 639298
rect 304901 639240 304906 639296
rect 304962 639240 307524 639296
rect 304901 639238 307524 639240
rect 281276 639236 281282 639238
rect 281165 639235 281231 639236
rect 304901 639235 304967 639238
rect 307518 639236 307524 639238
rect 307588 639236 307594 639300
rect 338021 639298 338087 639301
rect 342662 639298 342668 639300
rect 338021 639296 342668 639298
rect 338021 639240 338026 639296
rect 338082 639240 342668 639296
rect 338021 639238 342668 639240
rect 338021 639235 338087 639238
rect 342662 639236 342668 639238
rect 342732 639236 342738 639300
rect 362166 639236 362172 639300
rect 362236 639298 362242 639300
rect 365110 639298 365116 639300
rect 362236 639238 365116 639298
rect 362236 639236 362242 639238
rect 365110 639236 365116 639238
rect 365180 639236 365186 639300
rect 408534 639298 408540 639300
rect 403022 639238 408540 639298
rect 315982 639100 315988 639164
rect 316052 639162 316058 639164
rect 325550 639162 325556 639164
rect 316052 639102 325556 639162
rect 316052 639100 316058 639102
rect 325550 639100 325556 639102
rect 325620 639100 325626 639164
rect 333278 639100 333284 639164
rect 333348 639162 333354 639164
rect 336406 639162 336412 639164
rect 333348 639102 336412 639162
rect 333348 639100 333354 639102
rect 336406 639100 336412 639102
rect 336476 639100 336482 639164
rect 342478 639100 342484 639164
rect 342548 639162 342554 639164
rect 355542 639162 355548 639164
rect 342548 639102 355548 639162
rect 342548 639100 342554 639102
rect 355542 639100 355548 639102
rect 355612 639100 355618 639164
rect 364190 639100 364196 639164
rect 364260 639162 364266 639164
rect 374862 639162 374868 639164
rect 364260 639102 365546 639162
rect 364260 639100 364266 639102
rect 257654 638964 257660 639028
rect 257724 639026 257730 639028
rect 257724 638966 258090 639026
rect 257724 638964 257730 638966
rect 8109 638890 8175 638893
rect 17401 638890 17467 638893
rect 8109 638888 17467 638890
rect 8109 638832 8114 638888
rect 8170 638832 17406 638888
rect 17462 638832 17467 638888
rect 8109 638830 17467 638832
rect 8109 638827 8175 638830
rect 17401 638827 17467 638830
rect 26141 638890 26207 638893
rect 36721 638890 36787 638893
rect 26141 638888 36787 638890
rect 26141 638832 26146 638888
rect 26202 638832 36726 638888
rect 36782 638832 36787 638888
rect 26141 638830 36787 638832
rect 26141 638827 26207 638830
rect 36721 638827 36787 638830
rect 45461 638890 45527 638893
rect 56041 638890 56107 638893
rect 45461 638888 56107 638890
rect 45461 638832 45466 638888
rect 45522 638832 56046 638888
rect 56102 638832 56107 638888
rect 45461 638830 56107 638832
rect 45461 638827 45527 638830
rect 56041 638827 56107 638830
rect 64781 638890 64847 638893
rect 75361 638890 75427 638893
rect 64781 638888 75427 638890
rect 64781 638832 64786 638888
rect 64842 638832 75366 638888
rect 75422 638832 75427 638888
rect 64781 638830 75427 638832
rect 64781 638827 64847 638830
rect 75361 638827 75427 638830
rect 84101 638890 84167 638893
rect 94681 638890 94747 638893
rect 84101 638888 94747 638890
rect 84101 638832 84106 638888
rect 84162 638832 94686 638888
rect 94742 638832 94747 638888
rect 84101 638830 94747 638832
rect 84101 638827 84167 638830
rect 94681 638827 94747 638830
rect 103421 638890 103487 638893
rect 114001 638890 114067 638893
rect 103421 638888 114067 638890
rect 103421 638832 103426 638888
rect 103482 638832 114006 638888
rect 114062 638832 114067 638888
rect 103421 638830 114067 638832
rect 103421 638827 103487 638830
rect 114001 638827 114067 638830
rect 122741 638890 122807 638893
rect 133321 638890 133387 638893
rect 122741 638888 133387 638890
rect 122741 638832 122746 638888
rect 122802 638832 133326 638888
rect 133382 638832 133387 638888
rect 122741 638830 133387 638832
rect 122741 638827 122807 638830
rect 133321 638827 133387 638830
rect 142061 638890 142127 638893
rect 152641 638890 152707 638893
rect 142061 638888 152707 638890
rect 142061 638832 142066 638888
rect 142122 638832 152646 638888
rect 152702 638832 152707 638888
rect 142061 638830 152707 638832
rect 142061 638827 142127 638830
rect 152641 638827 152707 638830
rect 161381 638890 161447 638893
rect 171961 638890 172027 638893
rect 161381 638888 172027 638890
rect 161381 638832 161386 638888
rect 161442 638832 171966 638888
rect 172022 638832 172027 638888
rect 161381 638830 172027 638832
rect 161381 638827 161447 638830
rect 171961 638827 172027 638830
rect 180701 638890 180767 638893
rect 191281 638890 191347 638893
rect 180701 638888 191347 638890
rect 180701 638832 180706 638888
rect 180762 638832 191286 638888
rect 191342 638832 191347 638888
rect 180701 638830 191347 638832
rect 180701 638827 180767 638830
rect 191281 638827 191347 638830
rect 200021 638890 200087 638893
rect 210601 638890 210667 638893
rect 200021 638888 210667 638890
rect 200021 638832 200026 638888
rect 200082 638832 210606 638888
rect 210662 638832 210667 638888
rect 200021 638830 210667 638832
rect 200021 638827 200087 638830
rect 210601 638827 210667 638830
rect 219985 638890 220051 638893
rect 229870 638890 229876 638892
rect 219985 638888 229876 638890
rect 219985 638832 219990 638888
rect 220046 638832 229876 638888
rect 219985 638830 229876 638832
rect 219985 638827 220051 638830
rect 229870 638828 229876 638830
rect 229940 638828 229946 638892
rect 258030 638890 258090 638966
rect 277158 638964 277164 639028
rect 277228 639026 277234 639028
rect 277228 638966 277410 639026
rect 277228 638964 277234 638966
rect 277350 638892 277410 638966
rect 277526 638964 277532 639028
rect 277596 639026 277602 639028
rect 277596 638966 286794 639026
rect 277596 638964 277602 638966
rect 286734 638892 286794 638966
rect 286910 638964 286916 639028
rect 286980 639026 286986 639028
rect 286980 638966 316050 639026
rect 286980 638964 286986 638966
rect 267774 638890 267780 638892
rect 258030 638830 267780 638890
rect 267774 638828 267780 638830
rect 267844 638828 267850 638892
rect 277342 638828 277348 638892
rect 277412 638828 277418 638892
rect 286726 638828 286732 638892
rect 286796 638828 286802 638892
rect 315990 638890 316050 638966
rect 335302 638964 335308 639028
rect 335372 639026 335378 639028
rect 335372 638966 336290 639026
rect 335372 638964 335378 638966
rect 336230 638890 336290 638966
rect 355174 638964 355180 639028
rect 355244 639026 355250 639028
rect 362350 639026 362356 639028
rect 355244 638966 362356 639026
rect 355244 638964 355250 638966
rect 362350 638964 362356 638966
rect 362420 638964 362426 639028
rect 365486 639026 365546 639102
rect 370086 639102 374868 639162
rect 370086 639026 370146 639102
rect 374862 639100 374868 639102
rect 374932 639100 374938 639164
rect 384062 639100 384068 639164
rect 384132 639162 384138 639164
rect 398598 639162 398604 639164
rect 384132 639102 398604 639162
rect 384132 639100 384138 639102
rect 398598 639100 398604 639102
rect 398668 639100 398674 639164
rect 398966 639100 398972 639164
rect 399036 639162 399042 639164
rect 403022 639162 403082 639238
rect 408534 639236 408540 639238
rect 408604 639236 408610 639300
rect 408718 639236 408724 639300
rect 408788 639298 408794 639300
rect 415350 639298 415410 639646
rect 420177 639643 420243 639646
rect 417734 639508 417740 639572
rect 417804 639570 417810 639572
rect 422702 639570 422708 639572
rect 417804 639510 422708 639570
rect 417804 639508 417810 639510
rect 422702 639508 422708 639510
rect 422772 639508 422778 639572
rect 579797 639434 579863 639437
rect 583520 639434 584960 639524
rect 579797 639432 584960 639434
rect 579797 639376 579802 639432
rect 579858 639376 584960 639432
rect 579797 639374 584960 639376
rect 579797 639371 579863 639374
rect 408788 639238 415410 639298
rect 420177 639298 420243 639301
rect 430757 639298 430823 639301
rect 457161 639298 457227 639301
rect 462313 639300 462379 639301
rect 488625 639300 488691 639301
rect 509785 639300 509851 639301
rect 525425 639300 525491 639301
rect 462262 639298 462268 639300
rect 420177 639296 430823 639298
rect 420177 639240 420182 639296
rect 420238 639240 430762 639296
rect 430818 639240 430823 639296
rect 420177 639238 430823 639240
rect 408788 639236 408794 639238
rect 420177 639235 420243 639238
rect 430757 639235 430823 639238
rect 457118 639296 457227 639298
rect 457118 639240 457166 639296
rect 457222 639240 457227 639296
rect 457118 639235 457227 639240
rect 462222 639238 462268 639298
rect 462332 639296 462379 639300
rect 488574 639298 488580 639300
rect 462374 639240 462379 639296
rect 462262 639236 462268 639238
rect 462332 639236 462379 639240
rect 488534 639238 488580 639298
rect 488644 639296 488691 639300
rect 509734 639298 509740 639300
rect 488686 639240 488691 639296
rect 488574 639236 488580 639238
rect 488644 639236 488691 639240
rect 509694 639238 509740 639298
rect 509804 639296 509851 639300
rect 525374 639298 525380 639300
rect 509846 639240 509851 639296
rect 509734 639236 509740 639238
rect 509804 639236 509851 639240
rect 525334 639238 525380 639298
rect 525444 639296 525491 639300
rect 525486 639240 525491 639296
rect 525374 639236 525380 639238
rect 525444 639236 525491 639240
rect 527214 639236 527220 639300
rect 527284 639298 527290 639300
rect 528093 639298 528159 639301
rect 527284 639296 528159 639298
rect 527284 639240 528098 639296
rect 528154 639240 528159 639296
rect 583520 639284 584960 639374
rect 527284 639238 528159 639240
rect 527284 639236 527290 639238
rect 462313 639235 462379 639236
rect 488625 639235 488691 639236
rect 509785 639235 509851 639236
rect 525425 639235 525491 639236
rect 528093 639235 528159 639238
rect 399036 639102 403082 639162
rect 399036 639100 399042 639102
rect 362542 638966 364994 639026
rect 365486 638966 370146 639026
rect 342478 638890 342484 638892
rect 315990 638830 336106 638890
rect 336230 638830 342484 638890
rect 5257 638754 5323 638757
rect 336046 638754 336106 638830
rect 342478 638828 342484 638830
rect 342548 638828 342554 638892
rect 342662 638828 342668 638892
rect 342732 638890 342738 638892
rect 362542 638890 362602 638966
rect 342732 638830 362602 638890
rect 364934 638890 364994 638966
rect 374494 638964 374500 639028
rect 374564 639026 374570 639028
rect 374564 638966 384682 639026
rect 374564 638964 374570 638966
rect 384430 638890 384436 638892
rect 364934 638830 384436 638890
rect 342732 638828 342738 638830
rect 384430 638828 384436 638830
rect 384500 638828 384506 638892
rect 355174 638754 355180 638756
rect 5257 638752 335738 638754
rect 5257 638696 5262 638752
rect 5318 638696 335738 638752
rect 5257 638694 335738 638696
rect 336046 638694 355180 638754
rect 5257 638691 5323 638694
rect 5073 638618 5139 638621
rect 333278 638618 333284 638620
rect 5073 638616 333284 638618
rect 5073 638560 5078 638616
rect 5134 638560 333284 638616
rect 5073 638558 333284 638560
rect 5073 638555 5139 638558
rect 333278 638556 333284 638558
rect 333348 638556 333354 638620
rect 4889 638482 4955 638485
rect 6913 638482 6979 638485
rect 4889 638480 6979 638482
rect 4889 638424 4894 638480
rect 4950 638424 6918 638480
rect 6974 638424 6979 638480
rect 4889 638422 6979 638424
rect 4889 638419 4955 638422
rect 6913 638419 6979 638422
rect 17217 638482 17283 638485
rect 26233 638482 26299 638485
rect 17217 638480 26299 638482
rect 17217 638424 17222 638480
rect 17278 638424 26238 638480
rect 26294 638424 26299 638480
rect 17217 638422 26299 638424
rect 17217 638419 17283 638422
rect 26233 638419 26299 638422
rect 36537 638482 36603 638485
rect 45553 638482 45619 638485
rect 36537 638480 45619 638482
rect 36537 638424 36542 638480
rect 36598 638424 45558 638480
rect 45614 638424 45619 638480
rect 36537 638422 45619 638424
rect 36537 638419 36603 638422
rect 45553 638419 45619 638422
rect 55857 638482 55923 638485
rect 64873 638482 64939 638485
rect 55857 638480 64939 638482
rect 55857 638424 55862 638480
rect 55918 638424 64878 638480
rect 64934 638424 64939 638480
rect 55857 638422 64939 638424
rect 55857 638419 55923 638422
rect 64873 638419 64939 638422
rect 75177 638482 75243 638485
rect 84193 638482 84259 638485
rect 75177 638480 84259 638482
rect 75177 638424 75182 638480
rect 75238 638424 84198 638480
rect 84254 638424 84259 638480
rect 75177 638422 84259 638424
rect 75177 638419 75243 638422
rect 84193 638419 84259 638422
rect 94497 638482 94563 638485
rect 103513 638482 103579 638485
rect 94497 638480 103579 638482
rect 94497 638424 94502 638480
rect 94558 638424 103518 638480
rect 103574 638424 103579 638480
rect 94497 638422 103579 638424
rect 94497 638419 94563 638422
rect 103513 638419 103579 638422
rect 113817 638482 113883 638485
rect 122833 638482 122899 638485
rect 113817 638480 122899 638482
rect 113817 638424 113822 638480
rect 113878 638424 122838 638480
rect 122894 638424 122899 638480
rect 113817 638422 122899 638424
rect 113817 638419 113883 638422
rect 122833 638419 122899 638422
rect 133137 638482 133203 638485
rect 142153 638482 142219 638485
rect 133137 638480 142219 638482
rect 133137 638424 133142 638480
rect 133198 638424 142158 638480
rect 142214 638424 142219 638480
rect 133137 638422 142219 638424
rect 133137 638419 133203 638422
rect 142153 638419 142219 638422
rect 152457 638482 152523 638485
rect 161473 638482 161539 638485
rect 152457 638480 161539 638482
rect 152457 638424 152462 638480
rect 152518 638424 161478 638480
rect 161534 638424 161539 638480
rect 152457 638422 161539 638424
rect 152457 638419 152523 638422
rect 161473 638419 161539 638422
rect 171777 638482 171843 638485
rect 180793 638482 180859 638485
rect 171777 638480 180859 638482
rect 171777 638424 171782 638480
rect 171838 638424 180798 638480
rect 180854 638424 180859 638480
rect 171777 638422 180859 638424
rect 171777 638419 171843 638422
rect 180793 638419 180859 638422
rect 191097 638482 191163 638485
rect 200113 638482 200179 638485
rect 191097 638480 200179 638482
rect 191097 638424 191102 638480
rect 191158 638424 200118 638480
rect 200174 638424 200179 638480
rect 191097 638422 200179 638424
rect 191097 638419 191163 638422
rect 200113 638419 200179 638422
rect 210417 638482 210483 638485
rect 220077 638482 220143 638485
rect 210417 638480 220143 638482
rect 210417 638424 210422 638480
rect 210478 638424 220082 638480
rect 220138 638424 220143 638480
rect 210417 638422 220143 638424
rect 210417 638419 210483 638422
rect 220077 638419 220143 638422
rect 234286 638420 234292 638484
rect 234356 638482 234362 638484
rect 239438 638482 239444 638484
rect 234356 638422 239444 638482
rect 234356 638420 234362 638422
rect 239438 638420 239444 638422
rect 239508 638420 239514 638484
rect 244222 638420 244228 638484
rect 244292 638482 244298 638484
rect 258022 638482 258028 638484
rect 244292 638422 258028 638482
rect 244292 638420 244298 638422
rect 258022 638420 258028 638422
rect 258092 638420 258098 638484
rect 267590 638420 267596 638484
rect 267660 638482 267666 638484
rect 277526 638482 277532 638484
rect 267660 638422 277532 638482
rect 267660 638420 267666 638422
rect 277526 638420 277532 638422
rect 277596 638420 277602 638484
rect 286726 638420 286732 638484
rect 286796 638482 286802 638484
rect 296662 638482 296668 638484
rect 286796 638422 296668 638482
rect 286796 638420 286802 638422
rect 296662 638420 296668 638422
rect 296732 638420 296738 638484
rect 306598 638420 306604 638484
rect 306668 638482 306674 638484
rect 315982 638482 315988 638484
rect 306668 638422 315988 638482
rect 306668 638420 306674 638422
rect 315982 638420 315988 638422
rect 316052 638420 316058 638484
rect 325550 638420 325556 638484
rect 325620 638482 325626 638484
rect 335302 638482 335308 638484
rect 325620 638422 335308 638482
rect 325620 638420 325626 638422
rect 335302 638420 335308 638422
rect 335372 638420 335378 638484
rect 335678 638482 335738 638694
rect 355174 638692 355180 638694
rect 355244 638692 355250 638756
rect 355358 638692 355364 638756
rect 355428 638754 355434 638756
rect 362166 638754 362172 638756
rect 355428 638694 362172 638754
rect 355428 638692 355434 638694
rect 362166 638692 362172 638694
rect 362236 638692 362242 638756
rect 362350 638692 362356 638756
rect 362420 638754 362426 638756
rect 374494 638754 374500 638756
rect 362420 638694 374500 638754
rect 362420 638692 362426 638694
rect 374494 638692 374500 638694
rect 374564 638692 374570 638756
rect 374678 638692 374684 638756
rect 374748 638754 374754 638756
rect 384246 638754 384252 638756
rect 374748 638694 384252 638754
rect 374748 638692 374754 638694
rect 384246 638692 384252 638694
rect 384316 638692 384322 638756
rect 384622 638754 384682 638966
rect 402830 638964 402836 639028
rect 402900 639026 402906 639028
rect 402900 638966 403082 639026
rect 402900 638964 402906 638966
rect 384798 638828 384804 638892
rect 384868 638890 384874 638892
rect 384982 638890 384988 638892
rect 384868 638830 384988 638890
rect 384868 638828 384874 638830
rect 384982 638828 384988 638830
rect 385052 638828 385058 638892
rect 403022 638890 403082 638966
rect 408534 638964 408540 639028
rect 408604 639026 408610 639028
rect 408604 638966 409154 639026
rect 408604 638964 408610 638966
rect 408350 638890 408356 638892
rect 403022 638830 408356 638890
rect 408350 638828 408356 638830
rect 408420 638828 408426 638892
rect 408534 638828 408540 638892
rect 408604 638890 408610 638892
rect 409094 638890 409154 638966
rect 437238 638964 437244 639028
rect 437308 639026 437314 639028
rect 437308 638966 437674 639026
rect 437308 638964 437314 638966
rect 417918 638890 417924 638892
rect 408604 638830 408970 638890
rect 409094 638830 417924 638890
rect 408604 638828 408610 638830
rect 408718 638754 408724 638756
rect 384622 638694 408724 638754
rect 408718 638692 408724 638694
rect 408788 638692 408794 638756
rect 408910 638754 408970 638830
rect 417918 638828 417924 638830
rect 417988 638828 417994 638892
rect 437422 638890 437428 638892
rect 421974 638830 437428 638890
rect 421974 638754 422034 638830
rect 437422 638828 437428 638830
rect 437492 638828 437498 638892
rect 408910 638694 422034 638754
rect 422702 638692 422708 638756
rect 422772 638754 422778 638756
rect 437238 638754 437244 638756
rect 422772 638694 437244 638754
rect 422772 638692 422778 638694
rect 437238 638692 437244 638694
rect 437308 638692 437314 638756
rect 437614 638754 437674 638966
rect 456558 638964 456564 639028
rect 456628 639026 456634 639028
rect 457118 639026 457178 639235
rect 456628 638966 457178 639026
rect 456628 638964 456634 638966
rect 437790 638828 437796 638892
rect 437860 638890 437866 638892
rect 530301 638890 530367 638893
rect 437860 638888 530367 638890
rect 437860 638832 530306 638888
rect 530362 638832 530367 638888
rect 437860 638830 530367 638832
rect 437860 638828 437866 638830
rect 530301 638827 530367 638830
rect 456558 638754 456564 638756
rect 437614 638694 456564 638754
rect 456558 638692 456564 638694
rect 456628 638692 456634 638756
rect 336406 638556 336412 638620
rect 336476 638618 336482 638620
rect 462262 638618 462268 638620
rect 336476 638558 364442 638618
rect 336476 638556 336482 638558
rect 355358 638482 355364 638484
rect 335678 638422 355364 638482
rect 355358 638420 355364 638422
rect 355428 638420 355434 638484
rect 355542 638420 355548 638484
rect 355612 638482 355618 638484
rect 364190 638482 364196 638484
rect 355612 638422 364196 638482
rect 355612 638420 355618 638422
rect 364190 638420 364196 638422
rect 364260 638420 364266 638484
rect 364382 638482 364442 638558
rect 364750 638558 462268 638618
rect 364750 638482 364810 638558
rect 462262 638556 462268 638558
rect 462332 638556 462338 638620
rect 364382 638422 364810 638482
rect 365110 638420 365116 638484
rect 365180 638482 365186 638484
rect 374678 638482 374684 638484
rect 365180 638422 374684 638482
rect 365180 638420 365186 638422
rect 374678 638420 374684 638422
rect 374748 638420 374754 638484
rect 374862 638420 374868 638484
rect 374932 638482 374938 638484
rect 384062 638482 384068 638484
rect 374932 638422 384068 638482
rect 374932 638420 374938 638422
rect 384062 638420 384068 638422
rect 384132 638420 384138 638484
rect 384246 638420 384252 638484
rect 384316 638482 384322 638484
rect 417734 638482 417740 638484
rect 384316 638422 417740 638482
rect 384316 638420 384322 638422
rect 417734 638420 417740 638422
rect 417804 638420 417810 638484
rect 417918 638420 417924 638484
rect 417988 638482 417994 638484
rect 488574 638482 488580 638484
rect 417988 638422 488580 638482
rect 417988 638420 417994 638422
rect 488574 638420 488580 638422
rect 488644 638420 488650 638484
rect 525190 638420 525196 638484
rect 525260 638482 525266 638484
rect 529054 638482 529060 638484
rect 525260 638422 529060 638482
rect 525260 638420 525266 638422
rect 529054 638420 529060 638422
rect 529124 638420 529130 638484
rect 3693 638346 3759 638349
rect 509734 638346 509740 638348
rect 3693 638344 509740 638346
rect 3693 638288 3698 638344
rect 3754 638288 509740 638344
rect 3693 638286 509740 638288
rect 3693 638283 3759 638286
rect 509734 638284 509740 638286
rect 509804 638284 509810 638348
rect 525558 638284 525564 638348
rect 525628 638346 525634 638348
rect 530945 638346 531011 638349
rect 525628 638344 531011 638346
rect 525628 638288 530950 638344
rect 531006 638288 531011 638344
rect 525628 638286 531011 638288
rect 525628 638284 525634 638286
rect 530945 638283 531011 638286
rect 3417 638210 3483 638213
rect 525374 638210 525380 638212
rect 3417 638208 525380 638210
rect 3417 638152 3422 638208
rect 3478 638152 525380 638208
rect 3417 638150 525380 638152
rect 3417 638147 3483 638150
rect 525374 638148 525380 638150
rect 525444 638148 525450 638212
rect 6913 638074 6979 638077
rect 17217 638074 17283 638077
rect 6913 638072 17283 638074
rect 6913 638016 6918 638072
rect 6974 638016 17222 638072
rect 17278 638016 17283 638072
rect 6913 638014 17283 638016
rect 6913 638011 6979 638014
rect 17217 638011 17283 638014
rect 17401 638074 17467 638077
rect 26141 638074 26207 638077
rect 17401 638072 26207 638074
rect 17401 638016 17406 638072
rect 17462 638016 26146 638072
rect 26202 638016 26207 638072
rect 17401 638014 26207 638016
rect 17401 638011 17467 638014
rect 26141 638011 26207 638014
rect 26325 638074 26391 638077
rect 36537 638074 36603 638077
rect 26325 638072 36603 638074
rect 26325 638016 26330 638072
rect 26386 638016 36542 638072
rect 36598 638016 36603 638072
rect 26325 638014 36603 638016
rect 26325 638011 26391 638014
rect 36537 638011 36603 638014
rect 36721 638074 36787 638077
rect 45461 638074 45527 638077
rect 36721 638072 45527 638074
rect 36721 638016 36726 638072
rect 36782 638016 45466 638072
rect 45522 638016 45527 638072
rect 36721 638014 45527 638016
rect 36721 638011 36787 638014
rect 45461 638011 45527 638014
rect 45645 638074 45711 638077
rect 55857 638074 55923 638077
rect 45645 638072 55923 638074
rect 45645 638016 45650 638072
rect 45706 638016 55862 638072
rect 55918 638016 55923 638072
rect 45645 638014 55923 638016
rect 45645 638011 45711 638014
rect 55857 638011 55923 638014
rect 56041 638074 56107 638077
rect 64781 638074 64847 638077
rect 56041 638072 64847 638074
rect 56041 638016 56046 638072
rect 56102 638016 64786 638072
rect 64842 638016 64847 638072
rect 56041 638014 64847 638016
rect 56041 638011 56107 638014
rect 64781 638011 64847 638014
rect 64965 638074 65031 638077
rect 75177 638074 75243 638077
rect 64965 638072 75243 638074
rect 64965 638016 64970 638072
rect 65026 638016 75182 638072
rect 75238 638016 75243 638072
rect 64965 638014 75243 638016
rect 64965 638011 65031 638014
rect 75177 638011 75243 638014
rect 75361 638074 75427 638077
rect 84101 638074 84167 638077
rect 75361 638072 84167 638074
rect 75361 638016 75366 638072
rect 75422 638016 84106 638072
rect 84162 638016 84167 638072
rect 75361 638014 84167 638016
rect 75361 638011 75427 638014
rect 84101 638011 84167 638014
rect 84285 638074 84351 638077
rect 94497 638074 94563 638077
rect 84285 638072 94563 638074
rect 84285 638016 84290 638072
rect 84346 638016 94502 638072
rect 94558 638016 94563 638072
rect 84285 638014 94563 638016
rect 84285 638011 84351 638014
rect 94497 638011 94563 638014
rect 94681 638074 94747 638077
rect 103421 638074 103487 638077
rect 94681 638072 103487 638074
rect 94681 638016 94686 638072
rect 94742 638016 103426 638072
rect 103482 638016 103487 638072
rect 94681 638014 103487 638016
rect 94681 638011 94747 638014
rect 103421 638011 103487 638014
rect 103605 638074 103671 638077
rect 113817 638074 113883 638077
rect 103605 638072 113883 638074
rect 103605 638016 103610 638072
rect 103666 638016 113822 638072
rect 113878 638016 113883 638072
rect 103605 638014 113883 638016
rect 103605 638011 103671 638014
rect 113817 638011 113883 638014
rect 114001 638074 114067 638077
rect 122741 638074 122807 638077
rect 114001 638072 122807 638074
rect 114001 638016 114006 638072
rect 114062 638016 122746 638072
rect 122802 638016 122807 638072
rect 114001 638014 122807 638016
rect 114001 638011 114067 638014
rect 122741 638011 122807 638014
rect 122925 638074 122991 638077
rect 133137 638074 133203 638077
rect 122925 638072 133203 638074
rect 122925 638016 122930 638072
rect 122986 638016 133142 638072
rect 133198 638016 133203 638072
rect 122925 638014 133203 638016
rect 122925 638011 122991 638014
rect 133137 638011 133203 638014
rect 133321 638074 133387 638077
rect 142061 638074 142127 638077
rect 133321 638072 142127 638074
rect 133321 638016 133326 638072
rect 133382 638016 142066 638072
rect 142122 638016 142127 638072
rect 133321 638014 142127 638016
rect 133321 638011 133387 638014
rect 142061 638011 142127 638014
rect 142245 638074 142311 638077
rect 152457 638074 152523 638077
rect 142245 638072 152523 638074
rect 142245 638016 142250 638072
rect 142306 638016 152462 638072
rect 152518 638016 152523 638072
rect 142245 638014 152523 638016
rect 142245 638011 142311 638014
rect 152457 638011 152523 638014
rect 152641 638074 152707 638077
rect 161381 638074 161447 638077
rect 152641 638072 161447 638074
rect 152641 638016 152646 638072
rect 152702 638016 161386 638072
rect 161442 638016 161447 638072
rect 152641 638014 161447 638016
rect 152641 638011 152707 638014
rect 161381 638011 161447 638014
rect 161565 638074 161631 638077
rect 171777 638074 171843 638077
rect 161565 638072 171843 638074
rect 161565 638016 161570 638072
rect 161626 638016 171782 638072
rect 171838 638016 171843 638072
rect 161565 638014 171843 638016
rect 161565 638011 161631 638014
rect 171777 638011 171843 638014
rect 171961 638074 172027 638077
rect 180701 638074 180767 638077
rect 171961 638072 180767 638074
rect 171961 638016 171966 638072
rect 172022 638016 180706 638072
rect 180762 638016 180767 638072
rect 171961 638014 180767 638016
rect 171961 638011 172027 638014
rect 180701 638011 180767 638014
rect 180885 638074 180951 638077
rect 191097 638074 191163 638077
rect 180885 638072 191163 638074
rect 180885 638016 180890 638072
rect 180946 638016 191102 638072
rect 191158 638016 191163 638072
rect 180885 638014 191163 638016
rect 180885 638011 180951 638014
rect 191097 638011 191163 638014
rect 191281 638074 191347 638077
rect 200021 638074 200087 638077
rect 191281 638072 200087 638074
rect 191281 638016 191286 638072
rect 191342 638016 200026 638072
rect 200082 638016 200087 638072
rect 191281 638014 200087 638016
rect 191281 638011 191347 638014
rect 200021 638011 200087 638014
rect 200205 638074 200271 638077
rect 210417 638074 210483 638077
rect 200205 638072 210483 638074
rect 200205 638016 200210 638072
rect 200266 638016 210422 638072
rect 210478 638016 210483 638072
rect 200205 638014 210483 638016
rect 200205 638011 200271 638014
rect 210417 638011 210483 638014
rect 210601 638074 210667 638077
rect 219985 638074 220051 638077
rect 210601 638072 220051 638074
rect 210601 638016 210606 638072
rect 210662 638016 219990 638072
rect 220046 638016 220051 638072
rect 210601 638014 220051 638016
rect 210601 638011 210667 638014
rect 219985 638011 220051 638014
rect 229870 638012 229876 638076
rect 229940 638074 229946 638076
rect 257654 638074 257660 638076
rect 229940 638014 257660 638074
rect 229940 638012 229946 638014
rect 257654 638012 257660 638014
rect 257724 638012 257730 638076
rect 258022 638012 258028 638076
rect 258092 638074 258098 638076
rect 267590 638074 267596 638076
rect 258092 638014 267596 638074
rect 258092 638012 258098 638014
rect 267590 638012 267596 638014
rect 267660 638012 267666 638076
rect 273110 638012 273116 638076
rect 273180 638074 273186 638076
rect 525190 638074 525196 638076
rect 273180 638014 525196 638074
rect 273180 638012 273186 638014
rect 525190 638012 525196 638014
rect 525260 638012 525266 638076
rect 220077 637938 220143 637941
rect 234286 637938 234292 637940
rect 220077 637936 234292 637938
rect 220077 637880 220082 637936
rect 220138 637880 234292 637936
rect 220077 637878 234292 637880
rect 220077 637875 220143 637878
rect 234286 637876 234292 637878
rect 234356 637876 234362 637940
rect 239438 637876 239444 637940
rect 239508 637938 239514 637940
rect 244222 637938 244228 637940
rect 239508 637878 244228 637938
rect 239508 637876 239514 637878
rect 244222 637876 244228 637878
rect 244292 637876 244298 637940
rect 267774 637876 267780 637940
rect 267844 637938 267850 637940
rect 277158 637938 277164 637940
rect 267844 637878 277164 637938
rect 267844 637876 267850 637878
rect 277158 637876 277164 637878
rect 277228 637876 277234 637940
rect 281206 637876 281212 637940
rect 281276 637938 281282 637940
rect 530669 637938 530735 637941
rect 281276 637936 530735 637938
rect 281276 637880 530674 637936
rect 530730 637880 530735 637936
rect 281276 637878 530735 637880
rect 281276 637876 281282 637878
rect 530669 637875 530735 637878
rect 277342 637740 277348 637804
rect 277412 637802 277418 637804
rect 286910 637802 286916 637804
rect 277412 637742 286916 637802
rect 277412 637740 277418 637742
rect 286910 637740 286916 637742
rect 286980 637740 286986 637804
rect 296662 637740 296668 637804
rect 296732 637802 296738 637804
rect 306598 637802 306604 637804
rect 296732 637742 306604 637802
rect 296732 637740 296738 637742
rect 306598 637740 306604 637742
rect 306668 637740 306674 637804
rect 307518 637740 307524 637804
rect 307588 637802 307594 637804
rect 525558 637802 525564 637804
rect 307588 637742 525564 637802
rect 307588 637740 307594 637742
rect 525558 637740 525564 637742
rect 525628 637740 525634 637804
rect 527582 637468 527588 637532
rect 527652 637468 527658 637532
rect 527590 637394 527650 637468
rect 528134 637394 528140 637396
rect 527590 637334 528140 637394
rect 528134 637332 528140 637334
rect 528204 637332 528210 637396
rect 528134 628146 528140 628148
rect 527406 628086 528140 628146
rect 527406 628012 527466 628086
rect 528134 628084 528140 628086
rect 528204 628084 528210 628148
rect 527398 627948 527404 628012
rect 527468 627948 527474 628012
rect 580073 627738 580139 627741
rect 583520 627738 584960 627828
rect 580073 627736 584960 627738
rect 580073 627680 580078 627736
rect 580134 627680 584960 627736
rect 580073 627678 584960 627680
rect 580073 627675 580139 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3141 624882 3207 624885
rect -960 624880 3207 624882
rect -960 624824 3146 624880
rect 3202 624824 3207 624880
rect -960 624822 3207 624824
rect -960 624732 480 624822
rect 3141 624819 3207 624822
rect 527398 621012 527404 621076
rect 527468 621074 527474 621076
rect 528318 621074 528324 621076
rect 527468 621014 528324 621074
rect 527468 621012 527474 621014
rect 528318 621012 528324 621014
rect 528388 621012 528394 621076
rect 528318 618156 528324 618220
rect 528388 618156 528394 618220
rect 528326 618082 528386 618156
rect 528870 618082 528876 618084
rect 528326 618022 528876 618082
rect 528870 618020 528876 618022
rect 528940 618020 528946 618084
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 2773 610466 2839 610469
rect -960 610464 2839 610466
rect -960 610408 2778 610464
rect 2834 610408 2839 610464
rect -960 610406 2839 610408
rect -960 610316 480 610406
rect 2773 610403 2839 610406
rect 528502 608636 528508 608700
rect 528572 608698 528578 608700
rect 528870 608698 528876 608700
rect 528572 608638 528876 608698
rect 528572 608636 528578 608638
rect 528870 608636 528876 608638
rect 528940 608636 528946 608700
rect 580073 604210 580139 604213
rect 583520 604210 584960 604300
rect 580073 604208 584960 604210
rect 580073 604152 580078 604208
rect 580134 604152 584960 604208
rect 580073 604150 584960 604152
rect 580073 604147 580139 604150
rect 583520 604060 584960 604150
rect 527582 601700 527588 601764
rect 527652 601762 527658 601764
rect 528502 601762 528508 601764
rect 527652 601702 528508 601762
rect 527652 601700 527658 601702
rect 528502 601700 528508 601702
rect 528572 601700 528578 601764
rect -960 596050 480 596140
rect 3141 596050 3207 596053
rect -960 596048 3207 596050
rect -960 595992 3146 596048
rect 3202 595992 3207 596048
rect -960 595990 3207 595992
rect -960 595900 480 595990
rect 3141 595987 3207 595990
rect 580073 592514 580139 592517
rect 583520 592514 584960 592604
rect 580073 592512 584960 592514
rect 580073 592456 580078 592512
rect 580134 592456 584960 592512
rect 580073 592454 584960 592456
rect 580073 592451 580139 592454
rect 583520 592364 584960 592454
rect 527582 592180 527588 592244
rect 527652 592180 527658 592244
rect 527590 591972 527650 592180
rect 527582 591908 527588 591972
rect 527652 591908 527658 591972
rect 527398 589460 527404 589524
rect 527468 589522 527474 589524
rect 527582 589522 527588 589524
rect 527468 589462 527588 589522
rect 527468 589460 527474 589462
rect 527582 589460 527588 589462
rect 527652 589460 527658 589524
rect -960 581620 480 581860
rect 580073 580818 580139 580821
rect 583520 580818 584960 580908
rect 580073 580816 584960 580818
rect 580073 580760 580078 580816
rect 580134 580760 584960 580816
rect 580073 580758 584960 580760
rect 580073 580755 580139 580758
rect 583520 580668 584960 580758
rect 527214 570482 527220 570484
rect 527038 570422 527220 570482
rect 527038 570074 527098 570422
rect 527214 570420 527220 570422
rect 527284 570420 527290 570484
rect 527582 570210 527588 570212
rect 527406 570150 527588 570210
rect 527406 570076 527466 570150
rect 527582 570148 527588 570150
rect 527652 570148 527658 570212
rect 527214 570074 527220 570076
rect 527038 570014 527220 570074
rect 527214 570012 527220 570014
rect 527284 570012 527290 570076
rect 527398 570012 527404 570076
rect 527468 570012 527474 570076
rect 583520 568836 584960 569076
rect 527398 568516 527404 568580
rect 527468 568578 527474 568580
rect 528134 568578 528140 568580
rect 527468 568518 528140 568578
rect 527468 568516 527474 568518
rect 528134 568516 528140 568518
rect 528204 568516 528210 568580
rect -960 567354 480 567444
rect 3141 567354 3207 567357
rect -960 567352 3207 567354
rect -960 567296 3146 567352
rect 3202 567296 3207 567352
rect -960 567294 3207 567296
rect -960 567204 480 567294
rect 3141 567291 3207 567294
rect 528134 559194 528140 559196
rect 527590 559134 528140 559194
rect 527590 559060 527650 559134
rect 528134 559132 528140 559134
rect 528204 559132 528210 559196
rect 527582 558996 527588 559060
rect 527652 558996 527658 559060
rect 580073 557290 580139 557293
rect 583520 557290 584960 557380
rect 580073 557288 584960 557290
rect 580073 557232 580078 557288
rect 580134 557232 584960 557288
rect 580073 557230 584960 557232
rect 580073 557227 580139 557230
rect 583520 557140 584960 557230
rect 527582 553964 527588 554028
rect 527652 553964 527658 554028
rect 527590 553754 527650 553964
rect 527950 553754 527956 553756
rect 527590 553694 527956 553754
rect 527950 553692 527956 553694
rect 528020 553692 528026 553756
rect 527950 553346 527956 553348
rect 527590 553286 527956 553346
rect -960 553074 480 553164
rect 2773 553074 2839 553077
rect 527590 553076 527650 553286
rect 527950 553284 527956 553286
rect 528020 553284 528026 553348
rect -960 553072 2839 553074
rect -960 553016 2778 553072
rect 2834 553016 2839 553072
rect -960 553014 2839 553016
rect -960 552924 480 553014
rect 2773 553011 2839 553014
rect 527582 553012 527588 553076
rect 527652 553012 527658 553076
rect 580073 545594 580139 545597
rect 583520 545594 584960 545684
rect 580073 545592 584960 545594
rect 580073 545536 580078 545592
rect 580134 545536 584960 545592
rect 580073 545534 584960 545536
rect 580073 545531 580139 545534
rect 583520 545444 584960 545534
rect -960 538658 480 538748
rect 3233 538658 3299 538661
rect -960 538656 3299 538658
rect -960 538600 3238 538656
rect 3294 538600 3299 538656
rect -960 538598 3299 538600
rect -960 538508 480 538598
rect 3233 538595 3299 538598
rect 583520 533898 584960 533988
rect 583342 533838 584960 533898
rect 527582 533700 527588 533764
rect 527652 533700 527658 533764
rect 527590 532810 527650 533700
rect 538262 533022 547890 533082
rect 538262 532810 538322 533022
rect 547830 532946 547890 533022
rect 557582 533022 567210 533082
rect 547830 532886 557458 532946
rect 527590 532750 538322 532810
rect 557398 532810 557458 532886
rect 557582 532810 557642 533022
rect 567150 532946 567210 533022
rect 567150 532886 576778 532946
rect 557398 532750 557642 532810
rect 576718 532810 576778 532886
rect 583342 532810 583402 533838
rect 583520 533748 584960 533838
rect 576718 532750 583402 532810
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 527582 514796 527588 514860
rect 527652 514796 527658 514860
rect 527590 514724 527650 514796
rect 527582 514660 527588 514724
rect 527652 514660 527658 514724
rect 527582 512212 527588 512276
rect 527652 512274 527658 512276
rect 527652 512214 527834 512274
rect 527652 512212 527658 512214
rect 527774 512140 527834 512214
rect 527766 512076 527772 512140
rect 527836 512076 527842 512140
rect 580073 510370 580139 510373
rect 583520 510370 584960 510460
rect 580073 510368 584960 510370
rect 580073 510312 580078 510368
rect 580134 510312 584960 510368
rect 580073 510310 584960 510312
rect 580073 510307 580139 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3233 509962 3299 509965
rect -960 509960 3299 509962
rect -960 509904 3238 509960
rect 3294 509904 3299 509960
rect -960 509902 3299 509904
rect -960 509812 480 509902
rect 3233 509899 3299 509902
rect 527766 505202 527772 505204
rect 527406 505142 527772 505202
rect 527406 504932 527466 505142
rect 527766 505140 527772 505142
rect 527836 505140 527842 505204
rect 527398 504868 527404 504932
rect 527468 504868 527474 504932
rect 580073 498674 580139 498677
rect 583520 498674 584960 498764
rect 580073 498672 584960 498674
rect 580073 498616 580078 498672
rect 580134 498616 584960 498672
rect 580073 498614 584960 498616
rect 580073 498611 580139 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 2773 495546 2839 495549
rect -960 495544 2839 495546
rect -960 495488 2778 495544
rect 2834 495488 2839 495544
rect -960 495486 2839 495488
rect -960 495396 480 495486
rect 2773 495483 2839 495486
rect 527766 492492 527772 492556
rect 527836 492492 527842 492556
rect 527774 492418 527834 492492
rect 528134 492418 528140 492420
rect 527774 492358 528140 492418
rect 528134 492356 528140 492358
rect 528204 492356 528210 492420
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 527582 482972 527588 483036
rect 527652 483034 527658 483036
rect 528134 483034 528140 483036
rect 527652 482974 528140 483034
rect 527652 482972 527658 482974
rect 528134 482972 528140 482974
rect 528204 482972 528210 483036
rect -960 481130 480 481220
rect 3233 481130 3299 481133
rect -960 481128 3299 481130
rect -960 481072 3238 481128
rect 3294 481072 3299 481128
rect -960 481070 3299 481072
rect -960 480980 480 481070
rect 3233 481067 3299 481070
rect 583520 474996 584960 475236
rect 527582 471820 527588 471884
rect 527652 471820 527658 471884
rect 527590 471746 527650 471820
rect 527950 471746 527956 471748
rect 527590 471686 527956 471746
rect 527950 471684 527956 471686
rect 528020 471684 528026 471748
rect -960 466700 480 466940
rect 579797 463450 579863 463453
rect 583520 463450 584960 463540
rect 579797 463448 584960 463450
rect 579797 463392 579802 463448
rect 579858 463392 584960 463448
rect 579797 463390 584960 463392
rect 579797 463387 579863 463390
rect 583520 463300 584960 463390
rect 527950 462300 527956 462364
rect 528020 462362 528026 462364
rect 528134 462362 528140 462364
rect 528020 462302 528140 462362
rect 528020 462300 528026 462302
rect 528134 462300 528140 462302
rect 528204 462300 528210 462364
rect 527766 454004 527772 454068
rect 527836 454066 527842 454068
rect 528134 454066 528140 454068
rect 527836 454006 528140 454066
rect 527836 454004 527842 454006
rect 528134 454004 528140 454006
rect 528204 454004 528210 454068
rect -960 452434 480 452524
rect 3141 452434 3207 452437
rect -960 452432 3207 452434
rect -960 452376 3146 452432
rect 3202 452376 3207 452432
rect -960 452374 3207 452376
rect -960 452284 480 452374
rect 3141 452371 3207 452374
rect 580901 451754 580967 451757
rect 583520 451754 584960 451844
rect 580901 451752 584960 451754
rect 580901 451696 580906 451752
rect 580962 451696 584960 451752
rect 580901 451694 584960 451696
rect 580901 451691 580967 451694
rect 583520 451604 584960 451694
rect 527766 447266 527772 447268
rect 527590 447206 527772 447266
rect 527590 446996 527650 447206
rect 527766 447204 527772 447206
rect 527836 447204 527842 447268
rect 527582 446932 527588 446996
rect 527652 446932 527658 446996
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 2773 438018 2839 438021
rect -960 438016 2839 438018
rect -960 437960 2778 438016
rect 2834 437960 2839 438016
rect -960 437958 2839 437960
rect -960 437868 480 437958
rect 2773 437955 2839 437958
rect 527214 428300 527220 428364
rect 527284 428362 527290 428364
rect 527766 428362 527772 428364
rect 527284 428302 527772 428362
rect 527284 428300 527290 428302
rect 527766 428300 527772 428302
rect 527836 428300 527842 428364
rect 583520 428076 584960 428316
rect 527582 425098 527588 425100
rect 527038 425038 527588 425098
rect 527038 424962 527098 425038
rect 527582 425036 527588 425038
rect 527652 425036 527658 425100
rect 527582 424962 527588 424964
rect 527038 424902 527588 424962
rect 527582 424900 527588 424902
rect 527652 424900 527658 424964
rect -960 423738 480 423828
rect 3233 423738 3299 423741
rect -960 423736 3299 423738
rect -960 423680 3238 423736
rect 3294 423680 3299 423736
rect -960 423678 3299 423680
rect -960 423588 480 423678
rect 3233 423675 3299 423678
rect 527214 421636 527220 421700
rect 527284 421698 527290 421700
rect 527766 421698 527772 421700
rect 527284 421638 527772 421698
rect 527284 421636 527290 421638
rect 527766 421636 527772 421638
rect 527836 421636 527842 421700
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 580809 404834 580875 404837
rect 583520 404834 584960 404924
rect 580809 404832 584960 404834
rect 580809 404776 580814 404832
rect 580870 404776 584960 404832
rect 580809 404774 584960 404776
rect 580809 404771 580875 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 3325 395042 3391 395045
rect -960 395040 3391 395042
rect -960 394984 3330 395040
rect 3386 394984 3391 395040
rect -960 394982 3391 394984
rect -960 394892 480 394982
rect 3325 394979 3391 394982
rect 579613 393002 579679 393005
rect 583520 393002 584960 393092
rect 579613 393000 584960 393002
rect 579613 392944 579618 393000
rect 579674 392944 584960 393000
rect 579613 392942 584960 392944
rect 579613 392939 579679 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3233 380626 3299 380629
rect -960 380624 3299 380626
rect -960 380568 3238 380624
rect 3294 380568 3299 380624
rect -960 380566 3299 380568
rect -960 380476 480 380566
rect 3233 380563 3299 380566
rect 583520 369610 584960 369700
rect 583342 369550 584960 369610
rect 527582 368732 527588 368796
rect 527652 368794 527658 368796
rect 527652 368734 528570 368794
rect 527652 368732 527658 368734
rect 528510 368658 528570 368734
rect 538262 368734 547890 368794
rect 528510 368598 538138 368658
rect 538078 368522 538138 368598
rect 538262 368522 538322 368734
rect 547830 368658 547890 368734
rect 557582 368734 567210 368794
rect 547830 368598 557458 368658
rect 538078 368462 538322 368522
rect 557398 368522 557458 368598
rect 557582 368522 557642 368734
rect 567150 368658 567210 368734
rect 583342 368658 583402 369550
rect 583520 369460 584960 369550
rect 567150 368598 576778 368658
rect 557398 368462 557642 368522
rect 576718 368522 576778 368598
rect 576902 368598 583402 368658
rect 576902 368522 576962 368598
rect 576718 368462 576962 368522
rect -960 366210 480 366300
rect 2773 366210 2839 366213
rect -960 366208 2839 366210
rect -960 366152 2778 366208
rect 2834 366152 2839 366208
rect -960 366150 2839 366152
rect -960 366060 480 366150
rect 2773 366147 2839 366150
rect 580717 357914 580783 357917
rect 583520 357914 584960 358004
rect 580717 357912 584960 357914
rect 580717 357856 580722 357912
rect 580778 357856 584960 357912
rect 580717 357854 584960 357856
rect 580717 357851 580783 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 580165 346082 580231 346085
rect 583520 346082 584960 346172
rect 580165 346080 584960 346082
rect 580165 346024 580170 346080
rect 580226 346024 584960 346080
rect 580165 346022 584960 346024
rect 580165 346019 580231 346022
rect 583520 345932 584960 346022
rect 523217 337786 523283 337789
rect 529473 337786 529539 337789
rect 523217 337784 529539 337786
rect 523217 337728 523222 337784
rect 523278 337728 529478 337784
rect 529534 337728 529539 337784
rect 523217 337726 529539 337728
rect 523217 337723 523283 337726
rect 529473 337723 529539 337726
rect -960 337514 480 337604
rect 3325 337514 3391 337517
rect -960 337512 3391 337514
rect -960 337456 3330 337512
rect 3386 337456 3391 337512
rect -960 337454 3391 337456
rect -960 337364 480 337454
rect 3325 337451 3391 337454
rect 10317 337378 10383 337381
rect 232405 337378 232471 337381
rect 10317 337376 232471 337378
rect 10317 337320 10322 337376
rect 10378 337320 232410 337376
rect 232466 337320 232471 337376
rect 10317 337318 232471 337320
rect 10317 337315 10383 337318
rect 232405 337315 232471 337318
rect 528185 337378 528251 337381
rect 565077 337378 565143 337381
rect 528185 337376 565143 337378
rect 528185 337320 528190 337376
rect 528246 337320 565082 337376
rect 565138 337320 565143 337376
rect 528185 337318 565143 337320
rect 528185 337315 528251 337318
rect 565077 337315 565143 337318
rect 234286 336636 234292 336700
rect 234356 336636 234362 336700
rect 234294 336565 234354 336636
rect 234294 336560 234403 336565
rect 234294 336504 234342 336560
rect 234398 336504 234403 336560
rect 234294 336502 234403 336504
rect 234337 336499 234403 336502
rect 321921 335338 321987 335341
rect 322105 335338 322171 335341
rect 321921 335336 322171 335338
rect 321921 335280 321926 335336
rect 321982 335280 322110 335336
rect 322166 335280 322171 335336
rect 321921 335278 322171 335280
rect 321921 335275 321987 335278
rect 322105 335275 322171 335278
rect 451365 335338 451431 335341
rect 451825 335338 451891 335341
rect 451365 335336 451891 335338
rect 451365 335280 451370 335336
rect 451426 335280 451830 335336
rect 451886 335280 451891 335336
rect 451365 335278 451891 335280
rect 451365 335275 451431 335278
rect 451825 335275 451891 335278
rect 583520 334236 584960 334476
rect 347957 333978 348023 333981
rect 348233 333978 348299 333981
rect 347957 333976 348299 333978
rect 347957 333920 347962 333976
rect 348018 333920 348238 333976
rect 348294 333920 348299 333976
rect 347957 333918 348299 333920
rect 347957 333915 348023 333918
rect 348233 333915 348299 333918
rect 434161 328674 434227 328677
rect 433566 328672 434227 328674
rect 433566 328616 434166 328672
rect 434222 328616 434227 328672
rect 433566 328614 434227 328616
rect 433566 328538 433626 328614
rect 434161 328611 434227 328614
rect 433701 328538 433767 328541
rect 433566 328536 433767 328538
rect 433566 328480 433706 328536
rect 433762 328480 433767 328536
rect 433566 328478 433767 328480
rect 433701 328475 433767 328478
rect 293217 327314 293283 327317
rect 292622 327312 293283 327314
rect 292622 327256 293222 327312
rect 293278 327256 293283 327312
rect 292622 327254 293283 327256
rect 234337 327178 234403 327181
rect 234654 327178 234660 327180
rect 234337 327176 234660 327178
rect 234337 327120 234342 327176
rect 234398 327120 234660 327176
rect 234337 327118 234660 327120
rect 234337 327115 234403 327118
rect 234654 327116 234660 327118
rect 234724 327116 234730 327180
rect 292622 327178 292682 327254
rect 293217 327251 293283 327254
rect 292757 327178 292823 327181
rect 292622 327176 292823 327178
rect 292622 327120 292762 327176
rect 292818 327120 292823 327176
rect 292622 327118 292823 327120
rect 292757 327115 292823 327118
rect 294137 325682 294203 325685
rect 294321 325682 294387 325685
rect 294137 325680 294387 325682
rect 294137 325624 294142 325680
rect 294198 325624 294326 325680
rect 294382 325624 294387 325680
rect 294137 325622 294387 325624
rect 294137 325619 294203 325622
rect 294321 325619 294387 325622
rect 321461 325682 321527 325685
rect 321645 325682 321711 325685
rect 321461 325680 321711 325682
rect 321461 325624 321466 325680
rect 321522 325624 321650 325680
rect 321706 325624 321711 325680
rect 321461 325622 321711 325624
rect 321461 325619 321527 325622
rect 321645 325619 321711 325622
rect 352097 325682 352163 325685
rect 352281 325682 352347 325685
rect 352097 325680 352347 325682
rect 352097 325624 352102 325680
rect 352158 325624 352286 325680
rect 352342 325624 352347 325680
rect 352097 325622 352347 325624
rect 352097 325619 352163 325622
rect 352281 325619 352347 325622
rect 451549 325682 451615 325685
rect 451733 325682 451799 325685
rect 451549 325680 451799 325682
rect 451549 325624 451554 325680
rect 451610 325624 451738 325680
rect 451794 325624 451799 325680
rect 451549 325622 451799 325624
rect 451549 325619 451615 325622
rect 451733 325619 451799 325622
rect 3141 324322 3207 324325
rect 258942 324322 258948 324324
rect 3141 324320 258948 324322
rect 3141 324264 3146 324320
rect 3202 324264 258948 324320
rect 3141 324262 258948 324264
rect 3141 324259 3207 324262
rect 258942 324260 258948 324262
rect 259012 324260 259018 324324
rect -960 323098 480 323188
rect 3141 323098 3207 323101
rect -960 323096 3207 323098
rect -960 323040 3146 323096
rect 3202 323040 3207 323096
rect -960 323038 3207 323040
rect -960 322948 480 323038
rect 3141 323035 3207 323038
rect 579613 322690 579679 322693
rect 583520 322690 584960 322780
rect 579613 322688 584960 322690
rect 579613 322632 579618 322688
rect 579674 322632 584960 322688
rect 579613 322630 584960 322632
rect 579613 322627 579679 322630
rect 583520 322540 584960 322630
rect 234654 319018 234660 319020
rect 234294 318958 234660 319018
rect 234294 318884 234354 318958
rect 234654 318956 234660 318958
rect 234724 318956 234730 319020
rect 261017 319018 261083 319021
rect 381169 319018 381235 319021
rect 260974 319016 261083 319018
rect 260974 318960 261022 319016
rect 261078 318960 261083 319016
rect 260974 318955 261083 318960
rect 380942 319016 381235 319018
rect 380942 318960 381174 319016
rect 381230 318960 381235 319016
rect 380942 318958 381235 318960
rect 260974 318885 261034 318955
rect 234286 318820 234292 318884
rect 234356 318820 234362 318884
rect 260974 318880 261083 318885
rect 260974 318824 261022 318880
rect 261078 318824 261083 318880
rect 260974 318822 261083 318824
rect 261017 318819 261083 318822
rect 277301 318882 277367 318885
rect 277577 318882 277643 318885
rect 277301 318880 277643 318882
rect 277301 318824 277306 318880
rect 277362 318824 277582 318880
rect 277638 318824 277643 318880
rect 277301 318822 277643 318824
rect 380942 318882 381002 318958
rect 381169 318955 381235 318958
rect 381077 318882 381143 318885
rect 380942 318880 381143 318882
rect 380942 318824 381082 318880
rect 381138 318824 381143 318880
rect 380942 318822 381143 318824
rect 277301 318819 277367 318822
rect 277577 318819 277643 318822
rect 381077 318819 381143 318822
rect 324497 317658 324563 317661
rect 324270 317656 324563 317658
rect 324270 317600 324502 317656
rect 324558 317600 324563 317656
rect 324270 317598 324563 317600
rect 324270 317522 324330 317598
rect 324497 317595 324563 317598
rect 324405 317522 324471 317525
rect 324270 317520 324471 317522
rect 324270 317464 324410 317520
rect 324466 317464 324471 317520
rect 324270 317462 324471 317464
rect 324405 317459 324471 317462
rect 321461 316026 321527 316029
rect 321645 316026 321711 316029
rect 321461 316024 321711 316026
rect 321461 315968 321466 316024
rect 321522 315968 321650 316024
rect 321706 315968 321711 316024
rect 321461 315966 321711 315968
rect 321461 315963 321527 315966
rect 321645 315963 321711 315966
rect 324405 316026 324471 316029
rect 324681 316026 324747 316029
rect 324405 316024 324747 316026
rect 324405 315968 324410 316024
rect 324466 315968 324686 316024
rect 324742 315968 324747 316024
rect 324405 315966 324747 315968
rect 324405 315963 324471 315966
rect 324681 315963 324747 315966
rect 352097 316026 352163 316029
rect 352281 316026 352347 316029
rect 352097 316024 352347 316026
rect 352097 315968 352102 316024
rect 352158 315968 352286 316024
rect 352342 315968 352347 316024
rect 352097 315966 352347 315968
rect 352097 315963 352163 315966
rect 352281 315963 352347 315966
rect 357525 316026 357591 316029
rect 357709 316026 357775 316029
rect 357525 316024 357775 316026
rect 357525 315968 357530 316024
rect 357586 315968 357714 316024
rect 357770 315968 357775 316024
rect 357525 315966 357775 315968
rect 357525 315963 357591 315966
rect 357709 315963 357775 315966
rect 580625 310858 580691 310861
rect 583520 310858 584960 310948
rect 580625 310856 584960 310858
rect 580625 310800 580630 310856
rect 580686 310800 584960 310856
rect 580625 310798 584960 310800
rect 580625 310795 580691 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 2773 308818 2839 308821
rect -960 308816 2839 308818
rect -960 308760 2778 308816
rect 2834 308760 2839 308816
rect -960 308758 2839 308760
rect -960 308668 480 308758
rect 2773 308755 2839 308758
rect 261017 307730 261083 307733
rect 261201 307730 261267 307733
rect 261017 307728 261267 307730
rect 261017 307672 261022 307728
rect 261078 307672 261206 307728
rect 261262 307672 261267 307728
rect 261017 307670 261267 307672
rect 261017 307667 261083 307670
rect 261201 307667 261267 307670
rect 332685 306370 332751 306373
rect 332961 306370 333027 306373
rect 332685 306368 333027 306370
rect 332685 306312 332690 306368
rect 332746 306312 332966 306368
rect 333022 306312 333027 306368
rect 332685 306310 333027 306312
rect 332685 306307 332751 306310
rect 332961 306307 333027 306310
rect 234245 303108 234311 303109
rect 234245 303106 234292 303108
rect 234200 303104 234292 303106
rect 234200 303048 234250 303104
rect 234200 303046 234292 303048
rect 234245 303044 234292 303046
rect 234356 303044 234362 303108
rect 234245 303043 234311 303044
rect 234245 299706 234311 299709
rect 234245 299704 234354 299706
rect 234245 299648 234250 299704
rect 234306 299648 234354 299704
rect 234245 299643 234354 299648
rect 234294 299572 234354 299643
rect 234286 299508 234292 299572
rect 234356 299508 234362 299572
rect 309409 299434 309475 299437
rect 309593 299434 309659 299437
rect 309409 299432 309659 299434
rect 309409 299376 309414 299432
rect 309470 299376 309598 299432
rect 309654 299376 309659 299432
rect 309409 299374 309659 299376
rect 309409 299371 309475 299374
rect 309593 299371 309659 299374
rect 579705 299162 579771 299165
rect 583520 299162 584960 299252
rect 579705 299160 584960 299162
rect 579705 299104 579710 299160
rect 579766 299104 584960 299160
rect 579705 299102 584960 299104
rect 579705 299099 579771 299102
rect 583520 299012 584960 299102
rect 357525 296714 357591 296717
rect 357801 296714 357867 296717
rect 357525 296712 357867 296714
rect 357525 296656 357530 296712
rect 357586 296656 357806 296712
rect 357862 296656 357867 296712
rect 357525 296654 357867 296656
rect 357525 296651 357591 296654
rect 357801 296651 357867 296654
rect 236269 295354 236335 295357
rect 236545 295354 236611 295357
rect 236269 295352 236611 295354
rect 236269 295296 236274 295352
rect 236330 295296 236550 295352
rect 236606 295296 236611 295352
rect 236269 295294 236611 295296
rect 236269 295291 236335 295294
rect 236545 295291 236611 295294
rect -960 294402 480 294492
rect 3325 294402 3391 294405
rect -960 294400 3391 294402
rect -960 294344 3330 294400
rect 3386 294344 3391 294400
rect -960 294342 3391 294344
rect -960 294252 480 294342
rect 3325 294339 3391 294342
rect 234286 290396 234292 290460
rect 234356 290458 234362 290460
rect 234654 290458 234660 290460
rect 234356 290398 234660 290458
rect 234356 290396 234362 290398
rect 234654 290396 234660 290398
rect 234724 290396 234730 290460
rect 331397 290050 331463 290053
rect 331262 290048 331463 290050
rect 331262 289992 331402 290048
rect 331458 289992 331463 290048
rect 331262 289990 331463 289992
rect 331262 289781 331322 289990
rect 331397 289987 331463 289990
rect 281625 289778 281691 289781
rect 281901 289778 281967 289781
rect 281625 289776 281967 289778
rect 281625 289720 281630 289776
rect 281686 289720 281906 289776
rect 281962 289720 281967 289776
rect 281625 289718 281967 289720
rect 281625 289715 281691 289718
rect 281901 289715 281967 289718
rect 324497 289778 324563 289781
rect 324681 289778 324747 289781
rect 324497 289776 324747 289778
rect 324497 289720 324502 289776
rect 324558 289720 324686 289776
rect 324742 289720 324747 289776
rect 324497 289718 324747 289720
rect 331262 289776 331371 289781
rect 331262 289720 331310 289776
rect 331366 289720 331371 289776
rect 331262 289718 331371 289720
rect 324497 289715 324563 289718
rect 324681 289715 324747 289718
rect 331305 289715 331371 289718
rect 356513 288418 356579 288421
rect 356697 288418 356763 288421
rect 356513 288416 356763 288418
rect 356513 288360 356518 288416
rect 356574 288360 356702 288416
rect 356758 288360 356763 288416
rect 356513 288358 356763 288360
rect 356513 288355 356579 288358
rect 356697 288355 356763 288358
rect 451273 288418 451339 288421
rect 451457 288418 451523 288421
rect 451273 288416 451523 288418
rect 451273 288360 451278 288416
rect 451334 288360 451462 288416
rect 451518 288360 451523 288416
rect 451273 288358 451523 288360
rect 451273 288355 451339 288358
rect 451457 288355 451523 288358
rect 583520 287316 584960 287556
rect 352097 287058 352163 287061
rect 352281 287058 352347 287061
rect 352097 287056 352347 287058
rect 352097 287000 352102 287056
rect 352158 287000 352286 287056
rect 352342 287000 352347 287056
rect 352097 286998 352347 287000
rect 352097 286995 352163 286998
rect 352281 286995 352347 286998
rect -960 280122 480 280212
rect 3141 280122 3207 280125
rect -960 280120 3207 280122
rect -960 280064 3146 280120
rect 3202 280064 3207 280120
rect -960 280062 3207 280064
rect -960 279972 480 280062
rect 3141 280059 3207 280062
rect 243169 280122 243235 280125
rect 243353 280122 243419 280125
rect 243169 280120 243419 280122
rect 243169 280064 243174 280120
rect 243230 280064 243358 280120
rect 243414 280064 243419 280120
rect 243169 280062 243419 280064
rect 243169 280059 243235 280062
rect 243353 280059 243419 280062
rect 309409 280122 309475 280125
rect 309593 280122 309659 280125
rect 309409 280120 309659 280122
rect 309409 280064 309414 280120
rect 309470 280064 309598 280120
rect 309654 280064 309659 280120
rect 309409 280062 309659 280064
rect 309409 280059 309475 280062
rect 309593 280059 309659 280062
rect 265065 278762 265131 278765
rect 265341 278762 265407 278765
rect 265065 278760 265407 278762
rect 265065 278704 265070 278760
rect 265126 278704 265346 278760
rect 265402 278704 265407 278760
rect 265065 278702 265407 278704
rect 265065 278699 265131 278702
rect 265341 278699 265407 278702
rect 287237 278762 287303 278765
rect 287421 278762 287487 278765
rect 287237 278760 287487 278762
rect 287237 278704 287242 278760
rect 287298 278704 287426 278760
rect 287482 278704 287487 278760
rect 287237 278702 287487 278704
rect 287237 278699 287303 278702
rect 287421 278699 287487 278702
rect 298277 278762 298343 278765
rect 298553 278762 298619 278765
rect 392117 278762 392183 278765
rect 298277 278760 298619 278762
rect 298277 278704 298282 278760
rect 298338 278704 298558 278760
rect 298614 278704 298619 278760
rect 298277 278702 298619 278704
rect 298277 278699 298343 278702
rect 298553 278699 298619 278702
rect 391982 278760 392183 278762
rect 391982 278704 392122 278760
rect 392178 278704 392183 278760
rect 391982 278702 392183 278704
rect 391982 278626 392042 278702
rect 392117 278699 392183 278702
rect 393221 278762 393287 278765
rect 393405 278762 393471 278765
rect 393221 278760 393471 278762
rect 393221 278704 393226 278760
rect 393282 278704 393410 278760
rect 393466 278704 393471 278760
rect 393221 278702 393471 278704
rect 393221 278699 393287 278702
rect 393405 278699 393471 278702
rect 480161 278762 480227 278765
rect 480345 278762 480411 278765
rect 480161 278760 480411 278762
rect 480161 278704 480166 278760
rect 480222 278704 480350 278760
rect 480406 278704 480411 278760
rect 480161 278702 480411 278704
rect 480161 278699 480227 278702
rect 480345 278699 480411 278702
rect 392209 278626 392275 278629
rect 391982 278624 392275 278626
rect 391982 278568 392214 278624
rect 392270 278568 392275 278624
rect 391982 278566 392275 278568
rect 392209 278563 392275 278566
rect 236453 276178 236519 276181
rect 236134 276176 236519 276178
rect 236134 276120 236458 276176
rect 236514 276120 236519 276176
rect 236134 276118 236519 276120
rect 236134 276042 236194 276118
rect 236453 276115 236519 276118
rect 236269 276042 236335 276045
rect 236134 276040 236335 276042
rect 236134 275984 236274 276040
rect 236330 275984 236335 276040
rect 236134 275982 236335 275984
rect 236269 275979 236335 275982
rect 583520 275770 584960 275860
rect 583342 275710 584960 275770
rect 545665 274954 545731 274957
rect 534030 274952 545731 274954
rect 534030 274896 545670 274952
rect 545726 274896 545731 274952
rect 534030 274894 545731 274896
rect 529054 274620 529060 274684
rect 529124 274682 529130 274684
rect 534030 274682 534090 274894
rect 545665 274891 545731 274894
rect 550541 274954 550607 274957
rect 563053 274954 563119 274957
rect 550541 274952 563119 274954
rect 550541 274896 550546 274952
rect 550602 274896 563058 274952
rect 563114 274896 563119 274952
rect 550541 274894 563119 274896
rect 550541 274891 550607 274894
rect 563053 274891 563119 274894
rect 572621 274818 572687 274821
rect 569910 274816 572687 274818
rect 569910 274760 572626 274816
rect 572682 274760 572687 274816
rect 569910 274758 572687 274760
rect 569910 274682 569970 274758
rect 572621 274755 572687 274758
rect 529124 274622 534090 274682
rect 563286 274622 569970 274682
rect 572713 274682 572779 274685
rect 583342 274682 583402 275710
rect 583520 275620 584960 275710
rect 572713 274680 583402 274682
rect 572713 274624 572718 274680
rect 572774 274624 583402 274680
rect 572713 274622 583402 274624
rect 529124 274620 529130 274622
rect 563053 274546 563119 274549
rect 563286 274546 563346 274622
rect 572713 274619 572779 274622
rect 563053 274544 563346 274546
rect 563053 274488 563058 274544
rect 563114 274488 563346 274544
rect 563053 274486 563346 274488
rect 563053 274483 563119 274486
rect 234470 273458 234476 273460
rect 234110 273398 234476 273458
rect 234110 273324 234170 273398
rect 234470 273396 234476 273398
rect 234540 273396 234546 273460
rect 234102 273260 234108 273324
rect 234172 273260 234178 273324
rect 243353 270738 243419 270741
rect 331397 270738 331463 270741
rect 358997 270738 359063 270741
rect 364517 270738 364583 270741
rect 242942 270736 243419 270738
rect 242942 270680 243358 270736
rect 243414 270680 243419 270736
rect 242942 270678 243419 270680
rect 242942 270602 243002 270678
rect 243353 270675 243419 270678
rect 331262 270736 331463 270738
rect 331262 270680 331402 270736
rect 331458 270680 331463 270736
rect 331262 270678 331463 270680
rect 243077 270602 243143 270605
rect 242942 270600 243143 270602
rect 242942 270544 243082 270600
rect 243138 270544 243143 270600
rect 242942 270542 243143 270544
rect 243077 270539 243143 270542
rect 331262 270469 331322 270678
rect 331397 270675 331463 270678
rect 358862 270736 359063 270738
rect 358862 270680 359002 270736
rect 359058 270680 359063 270736
rect 358862 270678 359063 270680
rect 277669 270466 277735 270469
rect 277534 270464 277735 270466
rect 277534 270408 277674 270464
rect 277730 270408 277735 270464
rect 277534 270406 277735 270408
rect 331262 270464 331371 270469
rect 331262 270408 331310 270464
rect 331366 270408 331371 270464
rect 331262 270406 331371 270408
rect 358862 270466 358922 270678
rect 358997 270675 359063 270678
rect 364382 270736 364583 270738
rect 364382 270680 364522 270736
rect 364578 270680 364583 270736
rect 364382 270678 364583 270680
rect 359181 270466 359247 270469
rect 358862 270464 359247 270466
rect 358862 270408 359186 270464
rect 359242 270408 359247 270464
rect 358862 270406 359247 270408
rect 364382 270466 364442 270678
rect 364517 270675 364583 270678
rect 364609 270466 364675 270469
rect 364382 270464 364675 270466
rect 364382 270408 364614 270464
rect 364670 270408 364675 270464
rect 364382 270406 364675 270408
rect 277534 270330 277594 270406
rect 277669 270403 277735 270406
rect 331305 270403 331371 270406
rect 359181 270403 359247 270406
rect 364609 270403 364675 270406
rect 277761 270330 277827 270333
rect 277534 270328 277827 270330
rect 277534 270272 277766 270328
rect 277822 270272 277827 270328
rect 277534 270270 277827 270272
rect 277761 270267 277827 270270
rect 292665 269242 292731 269245
rect 292941 269242 293007 269245
rect 292665 269240 293007 269242
rect 292665 269184 292670 269240
rect 292726 269184 292946 269240
rect 293002 269184 293007 269240
rect 292665 269182 293007 269184
rect 292665 269179 292731 269182
rect 292941 269179 293007 269182
rect 351821 269106 351887 269109
rect 352097 269106 352163 269109
rect 351821 269104 352163 269106
rect 351821 269048 351826 269104
rect 351882 269048 352102 269104
rect 352158 269048 352163 269104
rect 351821 269046 352163 269048
rect 351821 269043 351887 269046
rect 352097 269043 352163 269046
rect 393221 269106 393287 269109
rect 393405 269106 393471 269109
rect 393221 269104 393471 269106
rect 393221 269048 393226 269104
rect 393282 269048 393410 269104
rect 393466 269048 393471 269104
rect 393221 269046 393471 269048
rect 393221 269043 393287 269046
rect 393405 269043 393471 269046
rect 254025 267746 254091 267749
rect 254209 267746 254275 267749
rect 254025 267744 254275 267746
rect 254025 267688 254030 267744
rect 254086 267688 254214 267744
rect 254270 267688 254275 267744
rect 254025 267686 254275 267688
rect 254025 267683 254091 267686
rect 254209 267683 254275 267686
rect 259545 267746 259611 267749
rect 259729 267746 259795 267749
rect 259545 267744 259795 267746
rect 259545 267688 259550 267744
rect 259606 267688 259734 267744
rect 259790 267688 259795 267744
rect 259545 267686 259795 267688
rect 259545 267683 259611 267686
rect 259729 267683 259795 267686
rect 347681 267746 347747 267749
rect 347865 267746 347931 267749
rect 347681 267744 347931 267746
rect 347681 267688 347686 267744
rect 347742 267688 347870 267744
rect 347926 267688 347931 267744
rect 347681 267686 347931 267688
rect 347681 267683 347747 267686
rect 347865 267683 347931 267686
rect 369945 267746 370011 267749
rect 370129 267746 370195 267749
rect 369945 267744 370195 267746
rect 369945 267688 369950 267744
rect 370006 267688 370134 267744
rect 370190 267688 370195 267744
rect 369945 267686 370195 267688
rect 369945 267683 370011 267686
rect 370129 267683 370195 267686
rect 375465 267746 375531 267749
rect 375649 267746 375715 267749
rect 375465 267744 375715 267746
rect 375465 267688 375470 267744
rect 375526 267688 375654 267744
rect 375710 267688 375715 267744
rect 375465 267686 375715 267688
rect 375465 267683 375531 267686
rect 375649 267683 375715 267686
rect 261886 266250 261892 266252
rect 614 266190 261892 266250
rect -960 265706 480 265796
rect 614 265706 674 266190
rect 261886 266188 261892 266190
rect 261956 266188 261962 266252
rect -960 265646 674 265706
rect -960 265556 480 265646
rect 580533 263938 580599 263941
rect 583520 263938 584960 264028
rect 580533 263936 584960 263938
rect 580533 263880 580538 263936
rect 580594 263880 584960 263936
rect 580533 263878 584960 263880
rect 580533 263875 580599 263878
rect 234102 263802 234108 263804
rect 233926 263742 234108 263802
rect 233926 263532 233986 263742
rect 234102 263740 234108 263742
rect 234172 263740 234178 263804
rect 583520 263788 584960 263878
rect 233918 263468 233924 263532
rect 233988 263468 233994 263532
rect 233918 262108 233924 262172
rect 233988 262108 233994 262172
rect 233926 262037 233986 262108
rect 233926 262032 234035 262037
rect 233926 261976 233974 262032
rect 234030 261976 234035 262032
rect 233926 261974 234035 261976
rect 233969 261971 234035 261974
rect 243169 260810 243235 260813
rect 243353 260810 243419 260813
rect 243169 260808 243419 260810
rect 243169 260752 243174 260808
rect 243230 260752 243358 260808
rect 243414 260752 243419 260808
rect 243169 260750 243419 260752
rect 243169 260747 243235 260750
rect 243353 260747 243419 260750
rect 270769 260810 270835 260813
rect 270953 260810 271019 260813
rect 270769 260808 271019 260810
rect 270769 260752 270774 260808
rect 270830 260752 270958 260808
rect 271014 260752 271019 260808
rect 270769 260750 271019 260752
rect 270769 260747 270835 260750
rect 270953 260747 271019 260750
rect 287237 259450 287303 259453
rect 480161 259450 480227 259453
rect 480345 259450 480411 259453
rect 287237 259448 287346 259450
rect 287237 259392 287242 259448
rect 287298 259392 287346 259448
rect 287237 259387 287346 259392
rect 480161 259448 480411 259450
rect 480161 259392 480166 259448
rect 480222 259392 480350 259448
rect 480406 259392 480411 259448
rect 480161 259390 480411 259392
rect 480161 259387 480227 259390
rect 480345 259387 480411 259390
rect 287286 259317 287346 259387
rect 287286 259312 287395 259317
rect 287286 259256 287334 259312
rect 287390 259256 287395 259312
rect 287286 259254 287395 259256
rect 287329 259251 287395 259254
rect 254025 258090 254091 258093
rect 254209 258090 254275 258093
rect 254025 258088 254275 258090
rect 254025 258032 254030 258088
rect 254086 258032 254214 258088
rect 254270 258032 254275 258088
rect 254025 258030 254275 258032
rect 254025 258027 254091 258030
rect 254209 258027 254275 258030
rect 259545 258090 259611 258093
rect 259729 258090 259795 258093
rect 259545 258088 259795 258090
rect 259545 258032 259550 258088
rect 259606 258032 259734 258088
rect 259790 258032 259795 258088
rect 259545 258030 259795 258032
rect 259545 258027 259611 258030
rect 259729 258027 259795 258030
rect 347681 258090 347747 258093
rect 348049 258090 348115 258093
rect 347681 258088 348115 258090
rect 347681 258032 347686 258088
rect 347742 258032 348054 258088
rect 348110 258032 348115 258088
rect 347681 258030 348115 258032
rect 347681 258027 347747 258030
rect 348049 258027 348115 258030
rect 369945 258090 370011 258093
rect 370129 258090 370195 258093
rect 369945 258088 370195 258090
rect 369945 258032 369950 258088
rect 370006 258032 370134 258088
rect 370190 258032 370195 258088
rect 369945 258030 370195 258032
rect 369945 258027 370011 258030
rect 370129 258027 370195 258030
rect 375465 258090 375531 258093
rect 375649 258090 375715 258093
rect 375465 258088 375715 258090
rect 375465 258032 375470 258088
rect 375526 258032 375654 258088
rect 375710 258032 375715 258088
rect 375465 258030 375715 258032
rect 375465 258027 375531 258030
rect 375649 258027 375715 258030
rect 235993 254010 236059 254013
rect 236269 254010 236335 254013
rect 235993 254008 236335 254010
rect 235993 253952 235998 254008
rect 236054 253952 236274 254008
rect 236330 253952 236335 254008
rect 235993 253950 236335 253952
rect 235993 253947 236059 253950
rect 236269 253947 236335 253950
rect 233969 252650 234035 252653
rect 234102 252650 234108 252652
rect 233969 252648 234108 252650
rect 233969 252592 233974 252648
rect 234030 252592 234108 252648
rect 233969 252590 234108 252592
rect 233969 252587 234035 252590
rect 234102 252588 234108 252590
rect 234172 252588 234178 252652
rect 3141 252514 3207 252517
rect 261702 252514 261708 252516
rect 3141 252512 233986 252514
rect 3141 252456 3146 252512
rect 3202 252456 233986 252512
rect 3141 252454 233986 252456
rect 3141 252451 3207 252454
rect 233926 252378 233986 252454
rect 234478 252454 261708 252514
rect 234478 252378 234538 252454
rect 261702 252452 261708 252454
rect 261772 252452 261778 252516
rect 233926 252318 234538 252378
rect 580441 252242 580507 252245
rect 583520 252242 584960 252332
rect 580441 252240 584960 252242
rect 580441 252184 580446 252240
rect 580502 252184 584960 252240
rect 580441 252182 584960 252184
rect 580441 252179 580507 252182
rect 583520 252092 584960 252182
rect 243353 251426 243419 251429
rect 242942 251424 243419 251426
rect -960 251290 480 251380
rect 242942 251368 243358 251424
rect 243414 251368 243419 251424
rect 242942 251366 243419 251368
rect 3141 251290 3207 251293
rect -960 251288 3207 251290
rect -960 251232 3146 251288
rect 3202 251232 3207 251288
rect -960 251230 3207 251232
rect 242942 251290 243002 251366
rect 243353 251363 243419 251366
rect 243077 251290 243143 251293
rect 242942 251288 243143 251290
rect 242942 251232 243082 251288
rect 243138 251232 243143 251288
rect 242942 251230 243143 251232
rect -960 251140 480 251230
rect 3141 251227 3207 251230
rect 243077 251227 243143 251230
rect 331121 251290 331187 251293
rect 331121 251288 331322 251290
rect 331121 251232 331126 251288
rect 331182 251232 331322 251288
rect 331121 251230 331322 251232
rect 331121 251227 331187 251230
rect 309317 251154 309383 251157
rect 309501 251154 309567 251157
rect 309317 251152 309567 251154
rect 309317 251096 309322 251152
rect 309378 251096 309506 251152
rect 309562 251096 309567 251152
rect 309317 251094 309567 251096
rect 309317 251091 309383 251094
rect 309501 251091 309567 251094
rect 331121 251154 331187 251157
rect 331262 251154 331322 251230
rect 331121 251152 331322 251154
rect 331121 251096 331126 251152
rect 331182 251096 331322 251152
rect 331121 251094 331322 251096
rect 342437 251154 342503 251157
rect 342621 251154 342687 251157
rect 342437 251152 342687 251154
rect 342437 251096 342442 251152
rect 342498 251096 342626 251152
rect 342682 251096 342687 251152
rect 342437 251094 342687 251096
rect 331121 251091 331187 251094
rect 342437 251091 342503 251094
rect 342621 251091 342687 251094
rect 287145 249794 287211 249797
rect 287421 249794 287487 249797
rect 287145 249792 287487 249794
rect 287145 249736 287150 249792
rect 287206 249736 287426 249792
rect 287482 249736 287487 249792
rect 287145 249734 287487 249736
rect 287145 249731 287211 249734
rect 287421 249731 287487 249734
rect 358997 249794 359063 249797
rect 359273 249794 359339 249797
rect 358997 249792 359339 249794
rect 358997 249736 359002 249792
rect 359058 249736 359278 249792
rect 359334 249736 359339 249792
rect 358997 249734 359339 249736
rect 358997 249731 359063 249734
rect 359273 249731 359339 249734
rect 392945 249794 393011 249797
rect 393129 249794 393195 249797
rect 392945 249792 393195 249794
rect 392945 249736 392950 249792
rect 393006 249736 393134 249792
rect 393190 249736 393195 249792
rect 392945 249734 393195 249736
rect 392945 249731 393011 249734
rect 393129 249731 393195 249734
rect 407481 249794 407547 249797
rect 407665 249794 407731 249797
rect 407481 249792 407731 249794
rect 407481 249736 407486 249792
rect 407542 249736 407670 249792
rect 407726 249736 407731 249792
rect 407481 249734 407731 249736
rect 407481 249731 407547 249734
rect 407665 249731 407731 249734
rect 356421 248434 356487 248437
rect 356605 248434 356671 248437
rect 356421 248432 356671 248434
rect 356421 248376 356426 248432
rect 356482 248376 356610 248432
rect 356666 248376 356671 248432
rect 356421 248374 356671 248376
rect 356421 248371 356487 248374
rect 356605 248371 356671 248374
rect 408769 248434 408835 248437
rect 408953 248434 409019 248437
rect 408769 248432 409019 248434
rect 408769 248376 408774 248432
rect 408830 248376 408958 248432
rect 409014 248376 409019 248432
rect 408769 248374 409019 248376
rect 408769 248371 408835 248374
rect 408953 248371 409019 248374
rect 234102 247692 234108 247756
rect 234172 247754 234178 247756
rect 234470 247754 234476 247756
rect 234172 247694 234476 247754
rect 234172 247692 234178 247694
rect 234470 247692 234476 247694
rect 234540 247692 234546 247756
rect 480345 241770 480411 241773
rect 480345 241768 480546 241770
rect 480345 241712 480350 241768
rect 480406 241712 480546 241768
rect 480345 241710 480546 241712
rect 480345 241707 480411 241710
rect 480345 241634 480411 241637
rect 480486 241634 480546 241710
rect 480345 241632 480546 241634
rect 480345 241576 480350 241632
rect 480406 241576 480546 241632
rect 480345 241574 480546 241576
rect 480345 241571 480411 241574
rect 271873 241498 271939 241501
rect 272057 241498 272123 241501
rect 271873 241496 272123 241498
rect 271873 241440 271878 241496
rect 271934 241440 272062 241496
rect 272118 241440 272123 241496
rect 271873 241438 272123 241440
rect 271873 241435 271939 241438
rect 272057 241435 272123 241438
rect 293953 241498 294019 241501
rect 294137 241498 294203 241501
rect 293953 241496 294203 241498
rect 293953 241440 293958 241496
rect 294014 241440 294142 241496
rect 294198 241440 294203 241496
rect 293953 241438 294203 241440
rect 293953 241435 294019 241438
rect 294137 241435 294203 241438
rect 305177 241498 305243 241501
rect 305361 241498 305427 241501
rect 305177 241496 305427 241498
rect 305177 241440 305182 241496
rect 305238 241440 305366 241496
rect 305422 241440 305427 241496
rect 305177 241438 305427 241440
rect 305177 241435 305243 241438
rect 305361 241435 305427 241438
rect 310697 241498 310763 241501
rect 310881 241498 310947 241501
rect 310697 241496 310947 241498
rect 310697 241440 310702 241496
rect 310758 241440 310886 241496
rect 310942 241440 310947 241496
rect 310697 241438 310947 241440
rect 310697 241435 310763 241438
rect 310881 241435 310947 241438
rect 346577 241498 346643 241501
rect 346761 241498 346827 241501
rect 346577 241496 346827 241498
rect 346577 241440 346582 241496
rect 346638 241440 346766 241496
rect 346822 241440 346827 241496
rect 346577 241438 346827 241440
rect 346577 241435 346643 241438
rect 346761 241435 346827 241438
rect 382273 241498 382339 241501
rect 382457 241498 382523 241501
rect 382273 241496 382523 241498
rect 382273 241440 382278 241496
rect 382334 241440 382462 241496
rect 382518 241440 382523 241496
rect 382273 241438 382523 241440
rect 382273 241435 382339 241438
rect 382457 241435 382523 241438
rect 392117 241498 392183 241501
rect 392301 241498 392367 241501
rect 392117 241496 392367 241498
rect 392117 241440 392122 241496
rect 392178 241440 392306 241496
rect 392362 241440 392367 241496
rect 392117 241438 392367 241440
rect 392117 241435 392183 241438
rect 392301 241435 392367 241438
rect 416865 241498 416931 241501
rect 417141 241498 417207 241501
rect 416865 241496 417207 241498
rect 416865 241440 416870 241496
rect 416926 241440 417146 241496
rect 417202 241440 417207 241496
rect 416865 241438 417207 241440
rect 416865 241435 416931 241438
rect 417141 241435 417207 241438
rect 433425 241498 433491 241501
rect 433609 241498 433675 241501
rect 433425 241496 433675 241498
rect 433425 241440 433430 241496
rect 433486 241440 433614 241496
rect 433670 241440 433675 241496
rect 433425 241438 433675 241440
rect 433425 241435 433491 241438
rect 433609 241435 433675 241438
rect 472065 241498 472131 241501
rect 472341 241498 472407 241501
rect 472065 241496 472407 241498
rect 472065 241440 472070 241496
rect 472126 241440 472346 241496
rect 472402 241440 472407 241496
rect 472065 241438 472407 241440
rect 472065 241435 472131 241438
rect 472341 241435 472407 241438
rect 583520 240396 584960 240636
rect 242709 240138 242775 240141
rect 242985 240138 243051 240141
rect 242709 240136 243051 240138
rect 242709 240080 242714 240136
rect 242770 240080 242990 240136
rect 243046 240080 243051 240136
rect 242709 240078 243051 240080
rect 242709 240075 242775 240078
rect 242985 240075 243051 240078
rect 266813 240138 266879 240141
rect 267089 240138 267155 240141
rect 266813 240136 267155 240138
rect 266813 240080 266818 240136
rect 266874 240080 267094 240136
rect 267150 240080 267155 240136
rect 266813 240078 267155 240080
rect 266813 240075 266879 240078
rect 267089 240075 267155 240078
rect 351821 240138 351887 240141
rect 352005 240138 352071 240141
rect 351821 240136 352071 240138
rect 351821 240080 351826 240136
rect 351882 240080 352010 240136
rect 352066 240080 352071 240136
rect 351821 240078 352071 240080
rect 351821 240075 351887 240078
rect 352005 240075 352071 240078
rect 392301 240138 392367 240141
rect 392485 240138 392551 240141
rect 392301 240136 392551 240138
rect 392301 240080 392306 240136
rect 392362 240080 392490 240136
rect 392546 240080 392551 240136
rect 392301 240078 392551 240080
rect 392301 240075 392367 240078
rect 392485 240075 392551 240078
rect 480161 240138 480227 240141
rect 480345 240138 480411 240141
rect 480161 240136 480411 240138
rect 480161 240080 480166 240136
rect 480222 240080 480350 240136
rect 480406 240080 480411 240136
rect 480161 240078 480411 240080
rect 480161 240075 480227 240078
rect 480345 240075 480411 240078
rect 259361 238778 259427 238781
rect 259545 238778 259611 238781
rect 259361 238776 259611 238778
rect 259361 238720 259366 238776
rect 259422 238720 259550 238776
rect 259606 238720 259611 238776
rect 259361 238718 259611 238720
rect 259361 238715 259427 238718
rect 259545 238715 259611 238718
rect 281901 238778 281967 238781
rect 282177 238778 282243 238781
rect 281901 238776 282243 238778
rect 281901 238720 281906 238776
rect 281962 238720 282182 238776
rect 282238 238720 282243 238776
rect 281901 238718 282243 238720
rect 281901 238715 281967 238718
rect 282177 238715 282243 238718
rect 356329 238778 356395 238781
rect 356513 238778 356579 238781
rect 356329 238776 356579 238778
rect 356329 238720 356334 238776
rect 356390 238720 356518 238776
rect 356574 238720 356579 238776
rect 356329 238718 356579 238720
rect 356329 238715 356395 238718
rect 356513 238715 356579 238718
rect -960 237010 480 237100
rect 2773 237010 2839 237013
rect -960 237008 2839 237010
rect -960 236952 2778 237008
rect 2834 236952 2839 237008
rect -960 236950 2839 236952
rect -960 236860 480 236950
rect 2773 236947 2839 236950
rect 252737 231842 252803 231845
rect 252921 231842 252987 231845
rect 252737 231840 252987 231842
rect 252737 231784 252742 231840
rect 252798 231784 252926 231840
rect 252982 231784 252987 231840
rect 252737 231782 252987 231784
rect 252737 231779 252803 231782
rect 252921 231779 252987 231782
rect 342437 231842 342503 231845
rect 342713 231842 342779 231845
rect 342437 231840 342779 231842
rect 342437 231784 342442 231840
rect 342498 231784 342718 231840
rect 342774 231784 342779 231840
rect 342437 231782 342779 231784
rect 342437 231779 342503 231782
rect 342713 231779 342779 231782
rect 386597 231842 386663 231845
rect 386873 231842 386939 231845
rect 386597 231840 386939 231842
rect 386597 231784 386602 231840
rect 386658 231784 386878 231840
rect 386934 231784 386939 231840
rect 386597 231782 386939 231784
rect 386597 231779 386663 231782
rect 386873 231779 386939 231782
rect 400397 231842 400463 231845
rect 400581 231842 400647 231845
rect 400397 231840 400647 231842
rect 400397 231784 400402 231840
rect 400458 231784 400586 231840
rect 400642 231784 400647 231840
rect 400397 231782 400647 231784
rect 400397 231779 400463 231782
rect 400581 231779 400647 231782
rect 266721 230482 266787 230485
rect 267089 230482 267155 230485
rect 266721 230480 267155 230482
rect 266721 230424 266726 230480
rect 266782 230424 267094 230480
rect 267150 230424 267155 230480
rect 266721 230422 267155 230424
rect 266721 230419 266787 230422
rect 267089 230419 267155 230422
rect 327257 230482 327323 230485
rect 327441 230482 327507 230485
rect 327257 230480 327507 230482
rect 327257 230424 327262 230480
rect 327318 230424 327446 230480
rect 327502 230424 327507 230480
rect 327257 230422 327507 230424
rect 327257 230419 327323 230422
rect 327441 230419 327507 230422
rect 351821 230482 351887 230485
rect 352097 230482 352163 230485
rect 351821 230480 352163 230482
rect 351821 230424 351826 230480
rect 351882 230424 352102 230480
rect 352158 230424 352163 230480
rect 351821 230422 352163 230424
rect 351821 230419 351887 230422
rect 352097 230419 352163 230422
rect 359089 229122 359155 229125
rect 359273 229122 359339 229125
rect 359089 229120 359339 229122
rect 359089 229064 359094 229120
rect 359150 229064 359278 229120
rect 359334 229064 359339 229120
rect 359089 229062 359339 229064
rect 359089 229059 359155 229062
rect 359273 229059 359339 229062
rect 580349 228850 580415 228853
rect 583520 228850 584960 228940
rect 580349 228848 584960 228850
rect 580349 228792 580354 228848
rect 580410 228792 584960 228848
rect 580349 228790 584960 228792
rect 580349 228787 580415 228790
rect 583520 228700 584960 228790
rect 234470 225178 234476 225180
rect 234294 225118 234476 225178
rect 234294 224908 234354 225118
rect 234470 225116 234476 225118
rect 234540 225116 234546 225180
rect 234286 224844 234292 224908
rect 234356 224844 234362 224908
rect -960 222594 480 222684
rect 4061 222594 4127 222597
rect -960 222592 4127 222594
rect -960 222536 4066 222592
rect 4122 222536 4127 222592
rect -960 222534 4127 222536
rect -960 222444 480 222534
rect 4061 222531 4127 222534
rect 271873 222186 271939 222189
rect 272057 222186 272123 222189
rect 271873 222184 272123 222186
rect 271873 222128 271878 222184
rect 271934 222128 272062 222184
rect 272118 222128 272123 222184
rect 271873 222126 272123 222128
rect 271873 222123 271939 222126
rect 272057 222123 272123 222126
rect 288433 222186 288499 222189
rect 288617 222186 288683 222189
rect 288433 222184 288683 222186
rect 288433 222128 288438 222184
rect 288494 222128 288622 222184
rect 288678 222128 288683 222184
rect 288433 222126 288683 222128
rect 288433 222123 288499 222126
rect 288617 222123 288683 222126
rect 293953 222186 294019 222189
rect 294137 222186 294203 222189
rect 293953 222184 294203 222186
rect 293953 222128 293958 222184
rect 294014 222128 294142 222184
rect 294198 222128 294203 222184
rect 293953 222126 294203 222128
rect 293953 222123 294019 222126
rect 294137 222123 294203 222126
rect 305177 222186 305243 222189
rect 305361 222186 305427 222189
rect 305177 222184 305427 222186
rect 305177 222128 305182 222184
rect 305238 222128 305366 222184
rect 305422 222128 305427 222184
rect 305177 222126 305427 222128
rect 305177 222123 305243 222126
rect 305361 222123 305427 222126
rect 308029 222186 308095 222189
rect 308305 222186 308371 222189
rect 308029 222184 308371 222186
rect 308029 222128 308034 222184
rect 308090 222128 308310 222184
rect 308366 222128 308371 222184
rect 308029 222126 308371 222128
rect 308029 222123 308095 222126
rect 308305 222123 308371 222126
rect 310697 222186 310763 222189
rect 310881 222186 310947 222189
rect 310697 222184 310947 222186
rect 310697 222128 310702 222184
rect 310758 222128 310886 222184
rect 310942 222128 310947 222184
rect 310697 222126 310947 222128
rect 310697 222123 310763 222126
rect 310881 222123 310947 222126
rect 346577 222186 346643 222189
rect 346761 222186 346827 222189
rect 346577 222184 346827 222186
rect 346577 222128 346582 222184
rect 346638 222128 346766 222184
rect 346822 222128 346827 222184
rect 346577 222126 346827 222128
rect 346577 222123 346643 222126
rect 346761 222123 346827 222126
rect 382273 222186 382339 222189
rect 382457 222186 382523 222189
rect 382273 222184 382523 222186
rect 382273 222128 382278 222184
rect 382334 222128 382462 222184
rect 382518 222128 382523 222184
rect 382273 222126 382523 222128
rect 382273 222123 382339 222126
rect 382457 222123 382523 222126
rect 392117 222186 392183 222189
rect 400305 222186 400371 222189
rect 400489 222186 400555 222189
rect 392117 222184 392226 222186
rect 392117 222128 392122 222184
rect 392178 222128 392226 222184
rect 392117 222123 392226 222128
rect 400305 222184 400555 222186
rect 400305 222128 400310 222184
rect 400366 222128 400494 222184
rect 400550 222128 400555 222184
rect 400305 222126 400555 222128
rect 400305 222123 400371 222126
rect 400489 222123 400555 222126
rect 416865 222186 416931 222189
rect 417141 222186 417207 222189
rect 416865 222184 417207 222186
rect 416865 222128 416870 222184
rect 416926 222128 417146 222184
rect 417202 222128 417207 222184
rect 416865 222126 417207 222128
rect 416865 222123 416931 222126
rect 417141 222123 417207 222126
rect 433425 222186 433491 222189
rect 433609 222186 433675 222189
rect 451273 222186 451339 222189
rect 433425 222184 433675 222186
rect 433425 222128 433430 222184
rect 433486 222128 433614 222184
rect 433670 222128 433675 222184
rect 433425 222126 433675 222128
rect 433425 222123 433491 222126
rect 433609 222123 433675 222126
rect 451230 222184 451339 222186
rect 451230 222128 451278 222184
rect 451334 222128 451339 222184
rect 451230 222123 451339 222128
rect 472065 222186 472131 222189
rect 472341 222186 472407 222189
rect 472065 222184 472407 222186
rect 472065 222128 472070 222184
rect 472126 222128 472346 222184
rect 472402 222128 472407 222184
rect 472065 222126 472407 222128
rect 472065 222123 472131 222126
rect 472341 222123 472407 222126
rect 392166 222053 392226 222123
rect 392166 222048 392275 222053
rect 392166 221992 392214 222048
rect 392270 221992 392275 222048
rect 392166 221990 392275 221992
rect 451230 222050 451290 222123
rect 451733 222050 451799 222053
rect 451230 222048 451799 222050
rect 451230 221992 451738 222048
rect 451794 221992 451799 222048
rect 451230 221990 451799 221992
rect 392209 221987 392275 221990
rect 451733 221987 451799 221990
rect 380801 220826 380867 220829
rect 381077 220826 381143 220829
rect 380801 220824 381143 220826
rect 380801 220768 380806 220824
rect 380862 220768 381082 220824
rect 381138 220768 381143 220824
rect 380801 220766 381143 220768
rect 380801 220763 380867 220766
rect 381077 220763 381143 220766
rect 480161 220826 480227 220829
rect 480345 220826 480411 220829
rect 480161 220824 480411 220826
rect 480161 220768 480166 220824
rect 480222 220768 480350 220824
rect 480406 220768 480411 220824
rect 480161 220766 480411 220768
rect 480161 220763 480227 220766
rect 480345 220763 480411 220766
rect 332777 219466 332843 219469
rect 333053 219466 333119 219469
rect 332777 219464 333119 219466
rect 332777 219408 332782 219464
rect 332838 219408 333058 219464
rect 333114 219408 333119 219464
rect 332777 219406 333119 219408
rect 332777 219403 332843 219406
rect 333053 219403 333119 219406
rect 580257 217018 580323 217021
rect 583520 217018 584960 217108
rect 580257 217016 584960 217018
rect 580257 216960 580262 217016
rect 580318 216960 584960 217016
rect 580257 216958 584960 216960
rect 580257 216955 580323 216958
rect 583520 216868 584960 216958
rect 342713 212802 342779 212805
rect 342302 212800 342779 212802
rect 342302 212744 342718 212800
rect 342774 212744 342779 212800
rect 342302 212742 342779 212744
rect 342302 212564 342362 212742
rect 342713 212739 342779 212742
rect 342437 212564 342503 212567
rect 342302 212562 342503 212564
rect 252737 212530 252803 212533
rect 252921 212530 252987 212533
rect 252737 212528 252987 212530
rect 252737 212472 252742 212528
rect 252798 212472 252926 212528
rect 252982 212472 252987 212528
rect 342302 212506 342442 212562
rect 342498 212506 342503 212562
rect 342302 212504 342503 212506
rect 342437 212501 342503 212504
rect 356421 212530 356487 212533
rect 356605 212530 356671 212533
rect 356421 212528 356671 212530
rect 252737 212470 252987 212472
rect 252737 212467 252803 212470
rect 252921 212467 252987 212470
rect 356421 212472 356426 212528
rect 356482 212472 356610 212528
rect 356666 212472 356671 212528
rect 356421 212470 356671 212472
rect 356421 212467 356487 212470
rect 356605 212467 356671 212470
rect 287329 211306 287395 211309
rect 287286 211304 287395 211306
rect 287286 211248 287334 211304
rect 287390 211248 287395 211304
rect 287286 211243 287395 211248
rect 287286 211173 287346 211243
rect 287237 211168 287346 211173
rect 287237 211112 287242 211168
rect 287298 211112 287346 211168
rect 287237 211110 287346 211112
rect 309317 211170 309383 211173
rect 309501 211170 309567 211173
rect 309317 211168 309567 211170
rect 309317 211112 309322 211168
rect 309378 211112 309506 211168
rect 309562 211112 309567 211168
rect 309317 211110 309567 211112
rect 287237 211107 287303 211110
rect 309317 211107 309383 211110
rect 309501 211107 309567 211110
rect 321737 211170 321803 211173
rect 321921 211170 321987 211173
rect 321737 211168 321987 211170
rect 321737 211112 321742 211168
rect 321798 211112 321926 211168
rect 321982 211112 321987 211168
rect 321737 211110 321987 211112
rect 321737 211107 321803 211110
rect 321921 211107 321987 211110
rect 324497 211170 324563 211173
rect 324681 211170 324747 211173
rect 324497 211168 324747 211170
rect 324497 211112 324502 211168
rect 324558 211112 324686 211168
rect 324742 211112 324747 211168
rect 324497 211110 324747 211112
rect 324497 211107 324563 211110
rect 324681 211107 324747 211110
rect 375649 211170 375715 211173
rect 375833 211170 375899 211173
rect 375649 211168 375899 211170
rect 375649 211112 375654 211168
rect 375710 211112 375838 211168
rect 375894 211112 375899 211168
rect 375649 211110 375899 211112
rect 375649 211107 375715 211110
rect 375833 211107 375899 211110
rect 380801 211170 380867 211173
rect 380985 211170 381051 211173
rect 380801 211168 381051 211170
rect 380801 211112 380806 211168
rect 380862 211112 380990 211168
rect 381046 211112 381051 211168
rect 380801 211110 381051 211112
rect 380801 211107 380867 211110
rect 380985 211107 381051 211110
rect 480161 211170 480227 211173
rect 480345 211170 480411 211173
rect 480161 211168 480411 211170
rect 480161 211112 480166 211168
rect 480222 211112 480350 211168
rect 480406 211112 480411 211168
rect 480161 211110 480411 211112
rect 480161 211107 480227 211110
rect 480345 211107 480411 211110
rect 263358 208524 263364 208588
rect 263428 208586 263434 208588
rect 278681 208586 278747 208589
rect 263428 208584 278747 208586
rect 263428 208528 278686 208584
rect 278742 208528 278747 208584
rect 263428 208526 278747 208528
rect 263428 208524 263434 208526
rect 278681 208523 278747 208526
rect 261518 208314 261524 208316
rect -960 208178 480 208268
rect 614 208254 261524 208314
rect 614 208178 674 208254
rect 261518 208252 261524 208254
rect 261588 208252 261594 208316
rect -960 208118 674 208178
rect -960 208028 480 208118
rect 234337 206954 234403 206957
rect 234470 206954 234476 206956
rect 234337 206952 234476 206954
rect 234337 206896 234342 206952
rect 234398 206896 234476 206952
rect 234337 206894 234476 206896
rect 234337 206891 234403 206894
rect 234470 206892 234476 206894
rect 234540 206892 234546 206956
rect 583520 205322 584960 205412
rect 583342 205262 584960 205322
rect 289813 204778 289879 204781
rect 300945 204778 301011 204781
rect 289813 204776 301011 204778
rect 289813 204720 289818 204776
rect 289874 204720 300950 204776
rect 301006 204720 301011 204776
rect 289813 204718 301011 204720
rect 289813 204715 289879 204718
rect 300945 204715 301011 204718
rect 362902 204716 362908 204780
rect 362972 204778 362978 204780
rect 372470 204778 372476 204780
rect 362972 204718 372476 204778
rect 362972 204716 362978 204718
rect 372470 204716 372476 204718
rect 372540 204716 372546 204780
rect 463366 204778 463372 204780
rect 456566 204718 463372 204778
rect 278681 204642 278747 204645
rect 434529 204642 434595 204645
rect 278681 204640 284954 204642
rect 278681 204584 278686 204640
rect 278742 204584 284954 204640
rect 278681 204582 284954 204584
rect 278681 204579 278747 204582
rect 284894 204506 284954 204582
rect 311758 204582 323594 204642
rect 289813 204506 289879 204509
rect 284894 204504 289879 204506
rect 284894 204448 289818 204504
rect 289874 204448 289879 204504
rect 284894 204446 289879 204448
rect 289813 204443 289879 204446
rect 300945 204370 301011 204373
rect 311758 204370 311818 204582
rect 323534 204506 323594 204582
rect 386462 204582 398850 204642
rect 362902 204506 362908 204508
rect 323534 204446 328562 204506
rect 300945 204368 311818 204370
rect 300945 204312 300950 204368
rect 301006 204312 311818 204368
rect 300945 204310 311818 204312
rect 328502 204370 328562 204446
rect 346580 204446 362908 204506
rect 336733 204370 336799 204373
rect 328502 204368 336799 204370
rect 328502 204312 336738 204368
rect 336794 204312 336799 204368
rect 328502 204310 336799 204312
rect 300945 204307 301011 204310
rect 336733 204307 336799 204310
rect 338113 204370 338179 204373
rect 346580 204370 346640 204446
rect 362902 204444 362908 204446
rect 362972 204444 362978 204508
rect 372470 204444 372476 204508
rect 372540 204506 372546 204508
rect 375189 204506 375255 204509
rect 372540 204504 375255 204506
rect 372540 204448 375194 204504
rect 375250 204448 375255 204504
rect 372540 204446 375255 204448
rect 372540 204444 372546 204446
rect 375189 204443 375255 204446
rect 384941 204506 385007 204509
rect 386462 204506 386522 204582
rect 384941 204504 386522 204506
rect 384941 204448 384946 204504
rect 385002 204448 386522 204504
rect 384941 204446 386522 204448
rect 384941 204443 385007 204446
rect 338113 204368 346640 204370
rect 338113 204312 338118 204368
rect 338174 204312 346640 204368
rect 338113 204310 346640 204312
rect 398790 204370 398850 204582
rect 434529 204640 437490 204642
rect 434529 204584 434534 204640
rect 434590 204584 437490 204640
rect 434529 204582 437490 204584
rect 434529 204579 434595 204582
rect 418061 204506 418127 204509
rect 408542 204504 418127 204506
rect 408542 204448 418066 204504
rect 418122 204448 418127 204504
rect 408542 204446 418127 204448
rect 408542 204370 408602 204446
rect 418061 204443 418127 204446
rect 425053 204370 425119 204373
rect 398790 204310 408602 204370
rect 424918 204368 425119 204370
rect 424918 204312 425058 204368
rect 425114 204312 425119 204368
rect 424918 204310 425119 204312
rect 437430 204370 437490 204582
rect 456566 204506 456626 204718
rect 463366 204716 463372 204718
rect 463436 204716 463442 204780
rect 502006 204778 502012 204780
rect 495206 204718 502012 204778
rect 495206 204506 495266 204718
rect 502006 204716 502012 204718
rect 502076 204716 502082 204780
rect 531262 204716 531268 204780
rect 531332 204778 531338 204780
rect 540881 204778 540947 204781
rect 531332 204776 540947 204778
rect 531332 204720 540886 204776
rect 540942 204720 540947 204776
rect 531332 204718 540947 204720
rect 531332 204716 531338 204718
rect 540881 204715 540947 204718
rect 560201 204642 560267 204645
rect 560201 204640 563162 204642
rect 560201 204584 560206 204640
rect 560262 204584 563162 204640
rect 560201 204582 563162 204584
rect 560201 204579 560267 204582
rect 514569 204506 514635 204509
rect 447182 204446 456626 204506
rect 466502 204446 482938 204506
rect 447182 204370 447242 204446
rect 437430 204310 447242 204370
rect 338113 204307 338179 204310
rect 418061 204098 418127 204101
rect 424918 204098 424978 204310
rect 425053 204307 425119 204310
rect 463550 204308 463556 204372
rect 463620 204370 463626 204372
rect 466502 204370 466562 204446
rect 463620 204310 466562 204370
rect 482878 204370 482938 204446
rect 485822 204446 495266 204506
rect 505142 204504 514635 204506
rect 505142 204448 514574 204504
rect 514630 204448 514635 204504
rect 505142 204446 514635 204448
rect 485822 204370 485882 204446
rect 482878 204310 485882 204370
rect 463620 204308 463626 204310
rect 502190 204308 502196 204372
rect 502260 204370 502266 204372
rect 505142 204370 505202 204446
rect 514569 204443 514635 204446
rect 526437 204506 526503 204509
rect 531262 204506 531268 204508
rect 526437 204504 531268 204506
rect 526437 204448 526442 204504
rect 526498 204448 531268 204504
rect 526437 204446 531268 204448
rect 526437 204443 526503 204446
rect 531262 204444 531268 204446
rect 531332 204444 531338 204508
rect 550582 204506 550588 204508
rect 543782 204446 550588 204506
rect 521653 204370 521719 204373
rect 502260 204310 505202 204370
rect 521518 204368 521719 204370
rect 521518 204312 521658 204368
rect 521714 204312 521719 204368
rect 521518 204310 521719 204312
rect 502260 204308 502266 204310
rect 418061 204096 424978 204098
rect 418061 204040 418066 204096
rect 418122 204040 424978 204096
rect 418061 204038 424978 204040
rect 514569 204098 514635 204101
rect 521518 204098 521578 204310
rect 521653 204307 521719 204310
rect 540881 204370 540947 204373
rect 543782 204370 543842 204446
rect 550582 204444 550588 204446
rect 550652 204444 550658 204508
rect 540881 204368 543842 204370
rect 540881 204312 540886 204368
rect 540942 204312 543842 204368
rect 540881 204310 543842 204312
rect 563102 204370 563162 204582
rect 572621 204506 572687 204509
rect 583342 204506 583402 205262
rect 583520 205172 584960 205262
rect 569910 204504 572687 204506
rect 569910 204448 572626 204504
rect 572682 204448 572687 204504
rect 569910 204446 572687 204448
rect 569910 204370 569970 204446
rect 572621 204443 572687 204446
rect 576902 204446 583402 204506
rect 563102 204310 569970 204370
rect 572713 204370 572779 204373
rect 576902 204370 576962 204446
rect 572713 204368 576962 204370
rect 572713 204312 572718 204368
rect 572774 204312 576962 204368
rect 572713 204310 576962 204312
rect 540881 204307 540947 204310
rect 572713 204307 572779 204310
rect 550582 204172 550588 204236
rect 550652 204234 550658 204236
rect 560201 204234 560267 204237
rect 550652 204232 560267 204234
rect 550652 204176 560206 204232
rect 560262 204176 560267 204232
rect 550652 204174 560267 204176
rect 550652 204172 550658 204174
rect 560201 204171 560267 204174
rect 514569 204096 521578 204098
rect 514569 204040 514574 204096
rect 514630 204040 521578 204096
rect 514569 204038 521578 204040
rect 418061 204035 418127 204038
rect 514569 204035 514635 204038
rect 252829 202874 252895 202877
rect 253013 202874 253079 202877
rect 252829 202872 253079 202874
rect 252829 202816 252834 202872
rect 252890 202816 253018 202872
rect 253074 202816 253079 202872
rect 252829 202814 253079 202816
rect 252829 202811 252895 202814
rect 253013 202811 253079 202814
rect 281717 202874 281783 202877
rect 281901 202874 281967 202877
rect 281717 202872 281967 202874
rect 281717 202816 281722 202872
rect 281778 202816 281906 202872
rect 281962 202816 281967 202872
rect 281717 202814 281967 202816
rect 281717 202811 281783 202814
rect 281901 202811 281967 202814
rect 288433 202874 288499 202877
rect 288617 202874 288683 202877
rect 288433 202872 288683 202874
rect 288433 202816 288438 202872
rect 288494 202816 288622 202872
rect 288678 202816 288683 202872
rect 288433 202814 288683 202816
rect 288433 202811 288499 202814
rect 288617 202811 288683 202814
rect 305177 202874 305243 202877
rect 305361 202874 305427 202877
rect 305177 202872 305427 202874
rect 305177 202816 305182 202872
rect 305238 202816 305366 202872
rect 305422 202816 305427 202872
rect 305177 202814 305427 202816
rect 305177 202811 305243 202814
rect 305361 202811 305427 202814
rect 308121 202874 308187 202877
rect 308305 202874 308371 202877
rect 308121 202872 308371 202874
rect 308121 202816 308126 202872
rect 308182 202816 308310 202872
rect 308366 202816 308371 202872
rect 308121 202814 308371 202816
rect 308121 202811 308187 202814
rect 308305 202811 308371 202814
rect 346577 202874 346643 202877
rect 346761 202874 346827 202877
rect 346577 202872 346827 202874
rect 346577 202816 346582 202872
rect 346638 202816 346766 202872
rect 346822 202816 346827 202872
rect 346577 202814 346827 202816
rect 346577 202811 346643 202814
rect 346761 202811 346827 202814
rect 382273 202874 382339 202877
rect 382457 202874 382523 202877
rect 382273 202872 382523 202874
rect 382273 202816 382278 202872
rect 382334 202816 382462 202872
rect 382518 202816 382523 202872
rect 382273 202814 382523 202816
rect 382273 202811 382339 202814
rect 382457 202811 382523 202814
rect 408677 202874 408743 202877
rect 408953 202874 409019 202877
rect 408677 202872 409019 202874
rect 408677 202816 408682 202872
rect 408738 202816 408958 202872
rect 409014 202816 409019 202872
rect 408677 202814 409019 202816
rect 408677 202811 408743 202814
rect 408953 202811 409019 202814
rect 416865 202874 416931 202877
rect 417141 202874 417207 202877
rect 416865 202872 417207 202874
rect 416865 202816 416870 202872
rect 416926 202816 417146 202872
rect 417202 202816 417207 202872
rect 416865 202814 417207 202816
rect 416865 202811 416931 202814
rect 417141 202811 417207 202814
rect 472065 202874 472131 202877
rect 472341 202874 472407 202877
rect 472065 202872 472407 202874
rect 472065 202816 472070 202872
rect 472126 202816 472346 202872
rect 472402 202816 472407 202872
rect 472065 202814 472407 202816
rect 472065 202811 472131 202814
rect 472341 202811 472407 202814
rect 255313 201514 255379 201517
rect 255589 201514 255655 201517
rect 255313 201512 255655 201514
rect 255313 201456 255318 201512
rect 255374 201456 255594 201512
rect 255650 201456 255655 201512
rect 255313 201454 255655 201456
rect 255313 201451 255379 201454
rect 255589 201451 255655 201454
rect 287145 201514 287211 201517
rect 287329 201514 287395 201517
rect 287145 201512 287395 201514
rect 287145 201456 287150 201512
rect 287206 201456 287334 201512
rect 287390 201456 287395 201512
rect 287145 201454 287395 201456
rect 287145 201451 287211 201454
rect 287329 201451 287395 201454
rect 351821 201514 351887 201517
rect 352097 201514 352163 201517
rect 351821 201512 352163 201514
rect 351821 201456 351826 201512
rect 351882 201456 352102 201512
rect 352158 201456 352163 201512
rect 351821 201454 352163 201456
rect 351821 201451 351887 201454
rect 352097 201451 352163 201454
rect 332685 200290 332751 200293
rect 332685 200288 332794 200290
rect 332685 200232 332690 200288
rect 332746 200232 332794 200288
rect 332685 200227 332794 200232
rect 359038 200228 359044 200292
rect 359108 200290 359114 200292
rect 359181 200290 359247 200293
rect 359108 200288 359247 200290
rect 359108 200232 359186 200288
rect 359242 200232 359247 200288
rect 359108 200230 359247 200232
rect 359108 200228 359114 200230
rect 359181 200227 359247 200230
rect 332734 200157 332794 200227
rect 331121 200154 331187 200157
rect 331397 200154 331463 200157
rect 331121 200152 331463 200154
rect 331121 200096 331126 200152
rect 331182 200096 331402 200152
rect 331458 200096 331463 200152
rect 331121 200094 331463 200096
rect 332734 200152 332843 200157
rect 332734 200096 332782 200152
rect 332838 200096 332843 200152
rect 332734 200094 332843 200096
rect 331121 200091 331187 200094
rect 331397 200091 331463 200094
rect 332777 200091 332843 200094
rect 359089 198796 359155 198797
rect 359038 198732 359044 198796
rect 359108 198794 359155 198796
rect 359108 198792 359200 198794
rect 359150 198736 359200 198792
rect 359108 198734 359200 198736
rect 359108 198732 359155 198734
rect 359089 198731 359155 198732
rect 234337 197570 234403 197573
rect 234294 197568 234403 197570
rect 234294 197512 234342 197568
rect 234398 197512 234403 197568
rect 234294 197507 234403 197512
rect 234294 197436 234354 197507
rect 234286 197372 234292 197436
rect 234356 197372 234362 197436
rect -960 193898 480 193988
rect 3969 193898 4035 193901
rect -960 193896 4035 193898
rect -960 193840 3974 193896
rect 4030 193840 4035 193896
rect -960 193838 4035 193840
rect -960 193748 480 193838
rect 3969 193835 4035 193838
rect 583520 193476 584960 193716
rect 252829 193218 252895 193221
rect 253013 193218 253079 193221
rect 252829 193216 253079 193218
rect 252829 193160 252834 193216
rect 252890 193160 253018 193216
rect 253074 193160 253079 193216
rect 252829 193158 253079 193160
rect 252829 193155 252895 193158
rect 253013 193155 253079 193158
rect 254117 193218 254183 193221
rect 254301 193218 254367 193221
rect 254117 193216 254367 193218
rect 254117 193160 254122 193216
rect 254178 193160 254306 193216
rect 254362 193160 254367 193216
rect 254117 193158 254367 193160
rect 254117 193155 254183 193158
rect 254301 193155 254367 193158
rect 259637 193218 259703 193221
rect 259821 193218 259887 193221
rect 259637 193216 259887 193218
rect 259637 193160 259642 193216
rect 259698 193160 259826 193216
rect 259882 193160 259887 193216
rect 259637 193158 259887 193160
rect 259637 193155 259703 193158
rect 259821 193155 259887 193158
rect 292757 193218 292823 193221
rect 292941 193218 293007 193221
rect 292757 193216 293007 193218
rect 292757 193160 292762 193216
rect 292818 193160 292946 193216
rect 293002 193160 293007 193216
rect 292757 193158 293007 193160
rect 292757 193155 292823 193158
rect 292941 193155 293007 193158
rect 321737 191858 321803 191861
rect 321921 191858 321987 191861
rect 321737 191856 321987 191858
rect 321737 191800 321742 191856
rect 321798 191800 321926 191856
rect 321982 191800 321987 191856
rect 321737 191798 321987 191800
rect 321737 191795 321803 191798
rect 321921 191795 321987 191798
rect 324497 191858 324563 191861
rect 324681 191858 324747 191861
rect 324497 191856 324747 191858
rect 324497 191800 324502 191856
rect 324558 191800 324686 191856
rect 324742 191800 324747 191856
rect 324497 191798 324747 191800
rect 324497 191795 324563 191798
rect 324681 191795 324747 191798
rect 342713 191858 342779 191861
rect 342897 191858 342963 191861
rect 342713 191856 342963 191858
rect 342713 191800 342718 191856
rect 342774 191800 342902 191856
rect 342958 191800 342963 191856
rect 342713 191798 342963 191800
rect 342713 191795 342779 191798
rect 342897 191795 342963 191798
rect 365713 191858 365779 191861
rect 365897 191858 365963 191861
rect 365713 191856 365963 191858
rect 365713 191800 365718 191856
rect 365774 191800 365902 191856
rect 365958 191800 365963 191856
rect 365713 191798 365963 191800
rect 365713 191795 365779 191798
rect 365897 191795 365963 191798
rect 364609 190498 364675 190501
rect 364793 190498 364859 190501
rect 364609 190496 364859 190498
rect 364609 190440 364614 190496
rect 364670 190440 364798 190496
rect 364854 190440 364859 190496
rect 364609 190438 364859 190440
rect 364609 190435 364675 190438
rect 364793 190435 364859 190438
rect 234286 187716 234292 187780
rect 234356 187778 234362 187780
rect 234470 187778 234476 187780
rect 234356 187718 234476 187778
rect 234356 187716 234362 187718
rect 234470 187716 234476 187718
rect 234540 187716 234546 187780
rect 234521 187508 234587 187509
rect 234470 187506 234476 187508
rect 234430 187446 234476 187506
rect 234540 187504 234587 187508
rect 234582 187448 234587 187504
rect 234470 187444 234476 187446
rect 234540 187444 234587 187448
rect 234521 187443 234587 187444
rect 243077 183698 243143 183701
rect 281993 183698 282059 183701
rect 243077 183696 243186 183698
rect 243077 183640 243082 183696
rect 243138 183640 243186 183696
rect 243077 183635 243186 183640
rect 241789 183562 241855 183565
rect 241973 183562 242039 183565
rect 241789 183560 242039 183562
rect 241789 183504 241794 183560
rect 241850 183504 241978 183560
rect 242034 183504 242039 183560
rect 241789 183502 242039 183504
rect 243126 183562 243186 183635
rect 281950 183696 282059 183698
rect 281950 183640 281998 183696
rect 282054 183640 282059 183696
rect 281950 183635 282059 183640
rect 243261 183562 243327 183565
rect 243126 183560 243327 183562
rect 243126 183504 243266 183560
rect 243322 183504 243327 183560
rect 243126 183502 243327 183504
rect 241789 183499 241855 183502
rect 241973 183499 242039 183502
rect 243261 183499 243327 183502
rect 266997 183562 267063 183565
rect 267181 183562 267247 183565
rect 266997 183560 267247 183562
rect 266997 183504 267002 183560
rect 267058 183504 267186 183560
rect 267242 183504 267247 183560
rect 266997 183502 267247 183504
rect 266997 183499 267063 183502
rect 267181 183499 267247 183502
rect 281950 183429 282010 183635
rect 288433 183562 288499 183565
rect 288617 183562 288683 183565
rect 288433 183560 288683 183562
rect 288433 183504 288438 183560
rect 288494 183504 288622 183560
rect 288678 183504 288683 183560
rect 288433 183502 288683 183504
rect 288433 183499 288499 183502
rect 288617 183499 288683 183502
rect 310697 183562 310763 183565
rect 310881 183562 310947 183565
rect 310697 183560 310947 183562
rect 310697 183504 310702 183560
rect 310758 183504 310886 183560
rect 310942 183504 310947 183560
rect 310697 183502 310947 183504
rect 310697 183499 310763 183502
rect 310881 183499 310947 183502
rect 408677 183562 408743 183565
rect 408953 183562 409019 183565
rect 408677 183560 409019 183562
rect 408677 183504 408682 183560
rect 408738 183504 408958 183560
rect 409014 183504 409019 183560
rect 408677 183502 409019 183504
rect 408677 183499 408743 183502
rect 408953 183499 409019 183502
rect 422385 183562 422451 183565
rect 422661 183562 422727 183565
rect 422385 183560 422727 183562
rect 422385 183504 422390 183560
rect 422446 183504 422666 183560
rect 422722 183504 422727 183560
rect 422385 183502 422727 183504
rect 422385 183499 422451 183502
rect 422661 183499 422727 183502
rect 472065 183562 472131 183565
rect 472341 183562 472407 183565
rect 472065 183560 472407 183562
rect 472065 183504 472070 183560
rect 472126 183504 472346 183560
rect 472402 183504 472407 183560
rect 472065 183502 472407 183504
rect 472065 183499 472131 183502
rect 472341 183499 472407 183502
rect 281950 183424 282059 183429
rect 281950 183368 281998 183424
rect 282054 183368 282059 183424
rect 281950 183366 282059 183368
rect 281993 183363 282059 183366
rect 382273 182202 382339 182205
rect 382457 182202 382523 182205
rect 382273 182200 382523 182202
rect 382273 182144 382278 182200
rect 382334 182144 382462 182200
rect 382518 182144 382523 182200
rect 382273 182142 382523 182144
rect 382273 182139 382339 182142
rect 382457 182139 382523 182142
rect 583520 181930 584960 182020
rect 583342 181870 584960 181930
rect 343541 181388 343607 181389
rect 343541 181386 343588 181388
rect 343500 181384 343588 181386
rect 343500 181328 343546 181384
rect 343500 181326 343588 181328
rect 343541 181324 343588 181326
rect 343652 181324 343658 181388
rect 343541 181323 343607 181324
rect 309041 181250 309107 181253
rect 343541 181250 343607 181253
rect 372613 181250 372679 181253
rect 294646 181248 309107 181250
rect 294646 181192 309046 181248
rect 309102 181192 309107 181248
rect 294646 181190 309107 181192
rect 257838 180916 257844 180980
rect 257908 180978 257914 180980
rect 294646 180978 294706 181190
rect 309041 181187 309107 181190
rect 334022 181248 343607 181250
rect 334022 181192 343546 181248
rect 343602 181192 343607 181248
rect 334022 181190 343607 181192
rect 318742 181114 318748 181116
rect 257908 180918 294706 180978
rect 313966 181054 318748 181114
rect 257908 180916 257914 180918
rect 309041 180842 309107 180845
rect 313966 180842 314026 181054
rect 318742 181052 318748 181054
rect 318812 181052 318818 181116
rect 334022 181114 334082 181190
rect 343541 181187 343607 181190
rect 372478 181248 372679 181250
rect 372478 181192 372618 181248
rect 372674 181192 372679 181248
rect 372478 181190 372679 181192
rect 331814 181054 334082 181114
rect 331814 180978 331874 181054
rect 343582 181052 343588 181116
rect 343652 181114 343658 181116
rect 343652 181054 360394 181114
rect 343652 181052 343658 181054
rect 323718 180918 331874 180978
rect 360334 180978 360394 181054
rect 361614 180978 361620 180980
rect 360334 180918 361620 180978
rect 309041 180840 314026 180842
rect 309041 180784 309046 180840
rect 309102 180784 314026 180840
rect 309041 180782 314026 180784
rect 309041 180779 309107 180782
rect 318742 180780 318748 180844
rect 318812 180842 318818 180844
rect 323718 180842 323778 180918
rect 361614 180916 361620 180918
rect 361684 180916 361690 180980
rect 371141 180978 371207 180981
rect 372478 180978 372538 181190
rect 372613 181187 372679 181190
rect 456566 181190 463618 181250
rect 434529 181114 434595 181117
rect 389222 181054 398850 181114
rect 371141 180976 372538 180978
rect 371141 180920 371146 180976
rect 371202 180920 372538 180976
rect 371141 180918 372538 180920
rect 382181 180978 382247 180981
rect 389222 180978 389282 181054
rect 382181 180976 389282 180978
rect 382181 180920 382186 180976
rect 382242 180920 389282 180976
rect 382181 180918 389282 180920
rect 371141 180915 371207 180918
rect 382181 180915 382247 180918
rect 318812 180782 323778 180842
rect 398790 180842 398850 181054
rect 434529 181112 437490 181114
rect 434529 181056 434534 181112
rect 434590 181056 437490 181112
rect 434529 181054 437490 181056
rect 434529 181051 434595 181054
rect 408542 180918 417986 180978
rect 408542 180842 408602 180918
rect 398790 180782 408602 180842
rect 417926 180842 417986 180918
rect 425053 180842 425119 180845
rect 417926 180840 425119 180842
rect 417926 180784 425058 180840
rect 425114 180784 425119 180840
rect 417926 180782 425119 180784
rect 437430 180842 437490 181054
rect 456566 180978 456626 181190
rect 463558 181116 463618 181190
rect 492630 181190 502258 181250
rect 463550 181052 463556 181116
rect 463620 181052 463626 181116
rect 475929 180978 475995 180981
rect 447182 180918 456626 180978
rect 466502 180976 475995 180978
rect 466502 180920 475934 180976
rect 475990 180920 475995 180976
rect 466502 180918 475995 180920
rect 447182 180842 447242 180918
rect 437430 180782 447242 180842
rect 318812 180780 318818 180782
rect 425053 180779 425119 180782
rect 463550 180780 463556 180844
rect 463620 180842 463626 180844
rect 466502 180842 466562 180918
rect 475929 180915 475995 180918
rect 476113 180978 476179 180981
rect 492630 180978 492690 181190
rect 502198 181116 502258 181190
rect 531262 181188 531268 181252
rect 531332 181250 531338 181252
rect 540881 181250 540947 181253
rect 531332 181248 540947 181250
rect 531332 181192 540886 181248
rect 540942 181192 540947 181248
rect 531332 181190 540947 181192
rect 531332 181188 531338 181190
rect 540881 181187 540947 181190
rect 502190 181052 502196 181116
rect 502260 181052 502266 181116
rect 583342 181114 583402 181870
rect 583520 181780 584960 181870
rect 572670 181054 583402 181114
rect 514569 180978 514635 180981
rect 476113 180976 482938 180978
rect 476113 180920 476118 180976
rect 476174 180920 482938 180976
rect 476113 180918 482938 180920
rect 476113 180915 476179 180918
rect 463620 180782 466562 180842
rect 482878 180842 482938 180918
rect 485822 180918 492690 180978
rect 505142 180976 514635 180978
rect 505142 180920 514574 180976
rect 514630 180920 514635 180976
rect 505142 180918 514635 180920
rect 485822 180842 485882 180918
rect 482878 180782 485882 180842
rect 463620 180780 463626 180782
rect 502190 180780 502196 180844
rect 502260 180842 502266 180844
rect 505142 180842 505202 180918
rect 514569 180915 514635 180918
rect 526437 180978 526503 180981
rect 531262 180978 531268 180980
rect 526437 180976 531268 180978
rect 526437 180920 526442 180976
rect 526498 180920 531268 180976
rect 526437 180918 531268 180920
rect 526437 180915 526503 180918
rect 531262 180916 531268 180918
rect 531332 180916 531338 180980
rect 553301 180978 553367 180981
rect 543782 180976 553367 180978
rect 543782 180920 553306 180976
rect 553362 180920 553367 180976
rect 543782 180918 553367 180920
rect 521653 180842 521719 180845
rect 502260 180782 505202 180842
rect 521518 180840 521719 180842
rect 521518 180784 521658 180840
rect 521714 180784 521719 180840
rect 521518 180782 521719 180784
rect 502260 180780 502266 180782
rect 3325 180706 3391 180709
rect 258758 180706 258764 180708
rect 3325 180704 258764 180706
rect 3325 180648 3330 180704
rect 3386 180648 258764 180704
rect 3325 180646 258764 180648
rect 3325 180643 3391 180646
rect 258758 180644 258764 180646
rect 258828 180644 258834 180708
rect 361614 180644 361620 180708
rect 361684 180706 361690 180708
rect 371141 180706 371207 180709
rect 361684 180704 371207 180706
rect 361684 180648 371146 180704
rect 371202 180648 371207 180704
rect 361684 180646 371207 180648
rect 361684 180644 361690 180646
rect 371141 180643 371207 180646
rect 514569 180570 514635 180573
rect 521518 180570 521578 180782
rect 521653 180779 521719 180782
rect 540881 180842 540947 180845
rect 543782 180842 543842 180918
rect 553301 180915 553367 180918
rect 554957 180978 555023 180981
rect 554957 180976 562978 180978
rect 554957 180920 554962 180976
rect 555018 180920 562978 180976
rect 554957 180918 562978 180920
rect 554957 180915 555023 180918
rect 540881 180840 543842 180842
rect 540881 180784 540886 180840
rect 540942 180784 543842 180840
rect 540881 180782 543842 180784
rect 562918 180842 562978 180918
rect 572670 180842 572730 181054
rect 562918 180782 572730 180842
rect 540881 180779 540947 180782
rect 514569 180568 521578 180570
rect 514569 180512 514574 180568
rect 514630 180512 521578 180568
rect 514569 180510 521578 180512
rect 514569 180507 514635 180510
rect -960 179482 480 179572
rect 3325 179482 3391 179485
rect -960 179480 3391 179482
rect -960 179424 3330 179480
rect 3386 179424 3391 179480
rect -960 179422 3391 179424
rect -960 179332 480 179422
rect 3325 179419 3391 179422
rect 234521 178122 234587 178125
rect 234654 178122 234660 178124
rect 234521 178120 234660 178122
rect 234521 178064 234526 178120
rect 234582 178064 234660 178120
rect 234521 178062 234660 178064
rect 234521 178059 234587 178062
rect 234654 178060 234660 178062
rect 234724 178060 234730 178124
rect 265249 177308 265315 177309
rect 265198 177244 265204 177308
rect 265268 177306 265315 177308
rect 265268 177304 265360 177306
rect 265310 177248 265360 177304
rect 265268 177246 265360 177248
rect 265268 177244 265315 177246
rect 265249 177243 265315 177244
rect 266445 173906 266511 173909
rect 266629 173906 266695 173909
rect 266445 173904 266695 173906
rect 266445 173848 266450 173904
rect 266506 173848 266634 173904
rect 266690 173848 266695 173904
rect 266445 173846 266695 173848
rect 266445 173843 266511 173846
rect 266629 173843 266695 173846
rect 287237 172546 287303 172549
rect 287421 172546 287487 172549
rect 287237 172544 287487 172546
rect 287237 172488 287242 172544
rect 287298 172488 287426 172544
rect 287482 172488 287487 172544
rect 287237 172486 287487 172488
rect 287237 172483 287303 172486
rect 287421 172483 287487 172486
rect 298185 172546 298251 172549
rect 298461 172546 298527 172549
rect 298185 172544 298527 172546
rect 298185 172488 298190 172544
rect 298246 172488 298466 172544
rect 298522 172488 298527 172544
rect 298185 172486 298527 172488
rect 298185 172483 298251 172486
rect 298461 172483 298527 172486
rect 342529 172546 342595 172549
rect 342897 172546 342963 172549
rect 342529 172544 342963 172546
rect 342529 172488 342534 172544
rect 342590 172488 342902 172544
rect 342958 172488 342963 172544
rect 342529 172486 342963 172488
rect 342529 172483 342595 172486
rect 342897 172483 342963 172486
rect 365713 172546 365779 172549
rect 365897 172546 365963 172549
rect 365713 172544 365963 172546
rect 365713 172488 365718 172544
rect 365774 172488 365902 172544
rect 365958 172488 365963 172544
rect 365713 172486 365963 172488
rect 365713 172483 365779 172486
rect 365897 172483 365963 172486
rect 261334 171260 261340 171324
rect 261404 171322 261410 171324
rect 268929 171322 268995 171325
rect 261404 171320 268995 171322
rect 261404 171264 268934 171320
rect 268990 171264 268995 171320
rect 261404 171262 268995 171264
rect 261404 171260 261410 171262
rect 268929 171259 268995 171262
rect 350398 170174 350642 170234
rect 268929 170098 268995 170101
rect 288341 170098 288407 170101
rect 268929 170096 288407 170098
rect 268929 170040 268934 170096
rect 268990 170040 288346 170096
rect 288402 170040 288407 170096
rect 268929 170038 288407 170040
rect 268929 170035 268995 170038
rect 288341 170035 288407 170038
rect 296621 170098 296687 170101
rect 298001 170098 298067 170101
rect 296621 170096 298067 170098
rect 296621 170040 296626 170096
rect 296682 170040 298006 170096
rect 298062 170040 298067 170096
rect 296621 170038 298067 170040
rect 296621 170035 296687 170038
rect 298001 170035 298067 170038
rect 317321 170098 317387 170101
rect 328361 170098 328427 170101
rect 317321 170096 328427 170098
rect 317321 170040 317326 170096
rect 317382 170040 328366 170096
rect 328422 170040 328427 170096
rect 317321 170038 328427 170040
rect 317321 170035 317387 170038
rect 328361 170035 328427 170038
rect 336641 170098 336707 170101
rect 336641 170096 342914 170098
rect 336641 170040 336646 170096
rect 336702 170040 342914 170096
rect 336641 170038 342914 170040
rect 336641 170035 336707 170038
rect 342854 169962 342914 170038
rect 350398 169962 350458 170174
rect 350582 170098 350642 170174
rect 495206 170174 502258 170234
rect 379329 170098 379395 170101
rect 350582 170038 357450 170098
rect 342854 169902 350458 169962
rect 357390 169962 357450 170038
rect 375238 170096 379395 170098
rect 375238 170040 379334 170096
rect 379390 170040 379395 170096
rect 375238 170038 379395 170040
rect 365713 169962 365779 169965
rect 357390 169960 365779 169962
rect 357390 169904 365718 169960
rect 365774 169904 365779 169960
rect 357390 169902 365779 169904
rect 365713 169899 365779 169902
rect 368289 169962 368355 169965
rect 375238 169962 375298 170038
rect 379329 170035 379395 170038
rect 379513 170098 379579 170101
rect 434529 170098 434595 170101
rect 379513 170096 381554 170098
rect 379513 170040 379518 170096
rect 379574 170040 381554 170096
rect 379513 170038 381554 170040
rect 379513 170035 379579 170038
rect 368289 169960 375298 169962
rect 368289 169904 368294 169960
rect 368350 169904 375298 169960
rect 368289 169902 375298 169904
rect 381494 169962 381554 170038
rect 386462 170038 398850 170098
rect 386462 169962 386522 170038
rect 381494 169902 386522 169962
rect 368289 169899 368355 169902
rect 298001 169826 298067 169829
rect 309041 169826 309107 169829
rect 298001 169824 298202 169826
rect 298001 169768 298006 169824
rect 298062 169768 298202 169824
rect 298001 169766 298202 169768
rect 298001 169763 298067 169766
rect 298142 169690 298202 169766
rect 307710 169824 309107 169826
rect 307710 169768 309046 169824
rect 309102 169768 309107 169824
rect 307710 169766 309107 169768
rect 398790 169826 398850 170038
rect 434529 170096 437490 170098
rect 434529 170040 434534 170096
rect 434590 170040 437490 170096
rect 434529 170038 437490 170040
rect 434529 170035 434595 170038
rect 418061 169962 418127 169965
rect 408542 169960 418127 169962
rect 408542 169904 418066 169960
rect 418122 169904 418127 169960
rect 408542 169902 418127 169904
rect 408542 169826 408602 169902
rect 418061 169899 418127 169902
rect 425053 169826 425119 169829
rect 398790 169766 408602 169826
rect 424918 169824 425119 169826
rect 424918 169768 425058 169824
rect 425114 169768 425119 169824
rect 424918 169766 425119 169768
rect 437430 169826 437490 170038
rect 454033 169962 454099 169965
rect 447182 169960 454099 169962
rect 447182 169904 454038 169960
rect 454094 169904 454099 169960
rect 447182 169902 454099 169904
rect 447182 169826 447242 169902
rect 454033 169899 454099 169902
rect 458173 169962 458239 169965
rect 475929 169962 475995 169965
rect 458173 169960 463618 169962
rect 458173 169904 458178 169960
rect 458234 169904 463618 169960
rect 458173 169902 463618 169904
rect 458173 169899 458239 169902
rect 437430 169766 447242 169826
rect 463558 169826 463618 169902
rect 466502 169960 475995 169962
rect 466502 169904 475934 169960
rect 475990 169904 475995 169960
rect 466502 169902 475995 169904
rect 466502 169826 466562 169902
rect 475929 169899 475995 169902
rect 476113 169962 476179 169965
rect 495206 169962 495266 170174
rect 476113 169960 482938 169962
rect 476113 169904 476118 169960
rect 476174 169904 482938 169960
rect 476113 169902 482938 169904
rect 476113 169899 476179 169902
rect 463558 169766 466562 169826
rect 482878 169826 482938 169902
rect 485822 169902 495266 169962
rect 485822 169826 485882 169902
rect 482878 169766 485882 169826
rect 502198 169826 502258 170174
rect 531262 170172 531268 170236
rect 531332 170234 531338 170236
rect 540881 170234 540947 170237
rect 531332 170232 540947 170234
rect 531332 170176 540886 170232
rect 540942 170176 540947 170232
rect 531332 170174 540947 170176
rect 531332 170172 531338 170174
rect 540881 170171 540947 170174
rect 560201 170098 560267 170101
rect 583520 170098 584960 170188
rect 560201 170096 563162 170098
rect 560201 170040 560206 170096
rect 560262 170040 563162 170096
rect 560201 170038 563162 170040
rect 560201 170035 560267 170038
rect 514569 169962 514635 169965
rect 505142 169960 514635 169962
rect 505142 169904 514574 169960
rect 514630 169904 514635 169960
rect 505142 169902 514635 169904
rect 505142 169826 505202 169902
rect 514569 169899 514635 169902
rect 516869 169962 516935 169965
rect 526437 169962 526503 169965
rect 531262 169962 531268 169964
rect 516869 169960 521578 169962
rect 516869 169904 516874 169960
rect 516930 169904 521578 169960
rect 516869 169902 521578 169904
rect 516869 169899 516935 169902
rect 502198 169766 505202 169826
rect 521518 169826 521578 169902
rect 526437 169960 531268 169962
rect 526437 169904 526442 169960
rect 526498 169904 531268 169960
rect 526437 169902 531268 169904
rect 526437 169899 526503 169902
rect 531262 169900 531268 169902
rect 531332 169900 531338 169964
rect 550582 169962 550588 169964
rect 543782 169902 550588 169962
rect 524229 169826 524295 169829
rect 521518 169824 524295 169826
rect 521518 169768 524234 169824
rect 524290 169768 524295 169824
rect 521518 169766 524295 169768
rect 299381 169690 299447 169693
rect 298142 169688 299447 169690
rect 298142 169632 299386 169688
rect 299442 169632 299447 169688
rect 298142 169630 299447 169632
rect 299381 169627 299447 169630
rect 302969 169690 303035 169693
rect 307710 169690 307770 169766
rect 309041 169763 309107 169766
rect 302969 169688 307770 169690
rect 302969 169632 302974 169688
rect 303030 169632 307770 169688
rect 302969 169630 307770 169632
rect 302969 169627 303035 169630
rect 418061 169554 418127 169557
rect 424918 169554 424978 169766
rect 425053 169763 425119 169766
rect 524229 169763 524295 169766
rect 540881 169826 540947 169829
rect 543782 169826 543842 169902
rect 550582 169900 550588 169902
rect 550652 169900 550658 169964
rect 540881 169824 543842 169826
rect 540881 169768 540886 169824
rect 540942 169768 543842 169824
rect 540881 169766 543842 169768
rect 563102 169826 563162 170038
rect 583342 170038 584960 170098
rect 572621 169962 572687 169965
rect 583342 169962 583402 170038
rect 569910 169960 572687 169962
rect 569910 169904 572626 169960
rect 572682 169904 572687 169960
rect 569910 169902 572687 169904
rect 569910 169826 569970 169902
rect 572621 169899 572687 169902
rect 576902 169902 583402 169962
rect 583520 169948 584960 170038
rect 563102 169766 569970 169826
rect 572713 169826 572779 169829
rect 576902 169826 576962 169902
rect 572713 169824 576962 169826
rect 572713 169768 572718 169824
rect 572774 169768 576962 169824
rect 572713 169766 576962 169768
rect 540881 169763 540947 169766
rect 572713 169763 572779 169766
rect 550582 169628 550588 169692
rect 550652 169690 550658 169692
rect 560201 169690 560267 169693
rect 550652 169688 560267 169690
rect 550652 169632 560206 169688
rect 560262 169632 560267 169688
rect 550652 169630 560267 169632
rect 550652 169628 550658 169630
rect 560201 169627 560267 169630
rect 418061 169552 424978 169554
rect 418061 169496 418066 169552
rect 418122 169496 424978 169552
rect 418061 169494 424978 169496
rect 418061 169491 418127 169494
rect -960 165066 480 165156
rect 2773 165066 2839 165069
rect -960 165064 2839 165066
rect -960 165008 2778 165064
rect 2834 165008 2839 165064
rect -960 165006 2839 165008
rect -960 164916 480 165006
rect 2773 165003 2839 165006
rect 321553 164386 321619 164389
rect 321510 164384 321619 164386
rect 321510 164328 321558 164384
rect 321614 164328 321619 164384
rect 321510 164323 321619 164328
rect 321510 164253 321570 164323
rect 265249 164252 265315 164253
rect 234286 164188 234292 164252
rect 234356 164250 234362 164252
rect 234654 164250 234660 164252
rect 234356 164190 234660 164250
rect 234356 164188 234362 164190
rect 234654 164188 234660 164190
rect 234724 164188 234730 164252
rect 265198 164250 265204 164252
rect 265158 164190 265204 164250
rect 265268 164248 265315 164252
rect 265310 164192 265315 164248
rect 265198 164188 265204 164190
rect 265268 164188 265315 164192
rect 265249 164187 265315 164188
rect 266997 164250 267063 164253
rect 267181 164250 267247 164253
rect 266997 164248 267247 164250
rect 266997 164192 267002 164248
rect 267058 164192 267186 164248
rect 267242 164192 267247 164248
rect 266997 164190 267247 164192
rect 321510 164248 321619 164253
rect 321510 164192 321558 164248
rect 321614 164192 321619 164248
rect 321510 164190 321619 164192
rect 266997 164187 267063 164190
rect 267181 164187 267247 164190
rect 321553 164187 321619 164190
rect 329925 164250 329991 164253
rect 330109 164250 330175 164253
rect 329925 164248 330175 164250
rect 329925 164192 329930 164248
rect 329986 164192 330114 164248
rect 330170 164192 330175 164248
rect 329925 164190 330175 164192
rect 329925 164187 329991 164190
rect 330109 164187 330175 164190
rect 376937 164250 377003 164253
rect 377121 164250 377187 164253
rect 376937 164248 377187 164250
rect 376937 164192 376942 164248
rect 376998 164192 377126 164248
rect 377182 164192 377187 164248
rect 376937 164190 377187 164192
rect 376937 164187 377003 164190
rect 377121 164187 377187 164190
rect 480345 164250 480411 164253
rect 480529 164250 480595 164253
rect 480345 164248 480595 164250
rect 480345 164192 480350 164248
rect 480406 164192 480534 164248
rect 480590 164192 480595 164248
rect 480345 164190 480595 164192
rect 480345 164187 480411 164190
rect 480529 164187 480595 164190
rect 236453 163026 236519 163029
rect 236272 163024 236519 163026
rect 236272 162968 236458 163024
rect 236514 162968 236519 163024
rect 236272 162966 236519 162968
rect 236272 162893 236332 162966
rect 236453 162963 236519 162966
rect 236269 162888 236335 162893
rect 236269 162832 236274 162888
rect 236330 162832 236335 162888
rect 236269 162827 236335 162832
rect 451825 162890 451891 162893
rect 452009 162890 452075 162893
rect 451825 162888 452075 162890
rect 451825 162832 451830 162888
rect 451886 162832 452014 162888
rect 452070 162832 452075 162888
rect 451825 162830 452075 162832
rect 451825 162827 451891 162830
rect 452009 162827 452075 162830
rect 583520 158402 584960 158492
rect 583342 158342 584960 158402
rect 307702 157796 307708 157860
rect 307772 157858 307778 157860
rect 317321 157858 317387 157861
rect 307772 157856 317387 157858
rect 307772 157800 317326 157856
rect 317382 157800 317387 157856
rect 307772 157798 317387 157800
rect 307772 157796 307778 157798
rect 317321 157795 317387 157798
rect 384982 157796 384988 157860
rect 385052 157858 385058 157860
rect 502006 157858 502012 157860
rect 385052 157798 386522 157858
rect 385052 157796 385058 157798
rect 386462 157722 386522 157798
rect 495206 157798 502012 157858
rect 405733 157722 405799 157725
rect 292438 157662 292682 157722
rect 255078 157524 255084 157588
rect 255148 157586 255154 157588
rect 278681 157586 278747 157589
rect 255148 157584 278747 157586
rect 255148 157528 278686 157584
rect 278742 157528 278747 157584
rect 255148 157526 278747 157528
rect 255148 157524 255154 157526
rect 278681 157523 278747 157526
rect 278681 157450 278747 157453
rect 292438 157450 292498 157662
rect 292622 157586 292682 157662
rect 333102 157662 333530 157722
rect 299422 157586 299428 157588
rect 292622 157526 299428 157586
rect 299422 157524 299428 157526
rect 299492 157524 299498 157588
rect 317321 157586 317387 157589
rect 317321 157584 323594 157586
rect 317321 157528 317326 157584
rect 317382 157528 323594 157584
rect 317321 157526 323594 157528
rect 317321 157523 317387 157526
rect 278681 157448 292498 157450
rect 278681 157392 278686 157448
rect 278742 157392 292498 157448
rect 278681 157390 292498 157392
rect 278681 157387 278747 157390
rect 299422 157388 299428 157452
rect 299492 157450 299498 157452
rect 307702 157450 307708 157452
rect 299492 157390 307708 157450
rect 299492 157388 299498 157390
rect 307702 157388 307708 157390
rect 307772 157388 307778 157452
rect 323534 157450 323594 157526
rect 333102 157450 333162 157662
rect 333470 157586 333530 157662
rect 340462 157662 340890 157722
rect 386462 157720 405799 157722
rect 386462 157664 405738 157720
rect 405794 157664 405799 157720
rect 386462 157662 405799 157664
rect 340462 157586 340522 157662
rect 333470 157526 340522 157586
rect 340830 157586 340890 157662
rect 405733 157659 405799 157662
rect 415301 157722 415367 157725
rect 417926 157722 418354 157756
rect 415301 157720 427738 157722
rect 415301 157664 415306 157720
rect 415362 157696 427738 157720
rect 415362 157664 417986 157696
rect 415301 157662 417986 157664
rect 418294 157662 427738 157696
rect 415301 157659 415367 157662
rect 375465 157586 375531 157589
rect 340830 157584 375531 157586
rect 340830 157528 375470 157584
rect 375526 157528 375531 157584
rect 340830 157526 375531 157528
rect 375465 157523 375531 157526
rect 323534 157390 333162 157450
rect 427678 157450 427738 157662
rect 427862 157662 437490 157722
rect 427862 157450 427922 157662
rect 427678 157390 427922 157450
rect 437430 157450 437490 157662
rect 456701 157586 456767 157589
rect 447182 157584 456767 157586
rect 447182 157528 456706 157584
rect 456762 157528 456767 157584
rect 447182 157526 456767 157528
rect 447182 157450 447242 157526
rect 456701 157523 456767 157526
rect 456885 157586 456951 157589
rect 495206 157586 495266 157798
rect 502006 157796 502012 157798
rect 502076 157796 502082 157860
rect 531262 157796 531268 157860
rect 531332 157858 531338 157860
rect 540881 157858 540947 157861
rect 531332 157856 540947 157858
rect 531332 157800 540886 157856
rect 540942 157800 540947 157856
rect 531332 157798 540947 157800
rect 531332 157796 531338 157798
rect 540881 157795 540947 157798
rect 560201 157722 560267 157725
rect 560201 157720 563162 157722
rect 560201 157664 560206 157720
rect 560262 157664 563162 157720
rect 560201 157662 563162 157664
rect 560201 157659 560267 157662
rect 514569 157586 514635 157589
rect 456885 157584 466378 157586
rect 456885 157528 456890 157584
rect 456946 157528 466378 157584
rect 456885 157526 466378 157528
rect 456885 157523 456951 157526
rect 437430 157390 447242 157450
rect 466318 157450 466378 157526
rect 466502 157526 475946 157586
rect 466502 157450 466562 157526
rect 466318 157390 466562 157450
rect 475886 157450 475946 157526
rect 485822 157526 495266 157586
rect 505142 157584 514635 157586
rect 505142 157528 514574 157584
rect 514630 157528 514635 157584
rect 505142 157526 514635 157528
rect 485822 157450 485882 157526
rect 475886 157390 485882 157450
rect 502190 157388 502196 157452
rect 502260 157450 502266 157452
rect 505142 157450 505202 157526
rect 514569 157523 514635 157526
rect 526437 157586 526503 157589
rect 531262 157586 531268 157588
rect 526437 157584 531268 157586
rect 526437 157528 526442 157584
rect 526498 157528 531268 157584
rect 526437 157526 531268 157528
rect 526437 157523 526503 157526
rect 531262 157524 531268 157526
rect 531332 157524 531338 157588
rect 550582 157586 550588 157588
rect 543782 157526 550588 157586
rect 521653 157450 521719 157453
rect 502260 157390 505202 157450
rect 521518 157448 521719 157450
rect 521518 157392 521658 157448
rect 521714 157392 521719 157448
rect 521518 157390 521719 157392
rect 502260 157388 502266 157390
rect 375465 157314 375531 157317
rect 384798 157314 384804 157316
rect 375465 157312 384804 157314
rect 375465 157256 375470 157312
rect 375526 157256 384804 157312
rect 375465 157254 384804 157256
rect 375465 157251 375531 157254
rect 384798 157252 384804 157254
rect 384868 157252 384874 157316
rect 514569 157178 514635 157181
rect 521518 157178 521578 157390
rect 521653 157387 521719 157390
rect 540881 157450 540947 157453
rect 543782 157450 543842 157526
rect 550582 157524 550588 157526
rect 550652 157524 550658 157588
rect 540881 157448 543842 157450
rect 540881 157392 540886 157448
rect 540942 157392 543842 157448
rect 540881 157390 543842 157392
rect 563102 157450 563162 157662
rect 572621 157586 572687 157589
rect 583342 157586 583402 158342
rect 583520 158252 584960 158342
rect 569910 157584 572687 157586
rect 569910 157528 572626 157584
rect 572682 157528 572687 157584
rect 569910 157526 572687 157528
rect 569910 157450 569970 157526
rect 572621 157523 572687 157526
rect 576902 157526 583402 157586
rect 563102 157390 569970 157450
rect 572713 157450 572779 157453
rect 576902 157450 576962 157526
rect 572713 157448 576962 157450
rect 572713 157392 572718 157448
rect 572774 157392 576962 157448
rect 572713 157390 576962 157392
rect 540881 157387 540947 157390
rect 572713 157387 572779 157390
rect 550582 157252 550588 157316
rect 550652 157314 550658 157316
rect 560201 157314 560267 157317
rect 550652 157312 560267 157314
rect 550652 157256 560206 157312
rect 560262 157256 560267 157312
rect 550652 157254 560267 157256
rect 550652 157252 550658 157254
rect 560201 157251 560267 157254
rect 514569 157176 521578 157178
rect 514569 157120 514574 157176
rect 514630 157120 521578 157176
rect 514569 157118 521578 157120
rect 514569 157115 514635 157118
rect 240225 154730 240291 154733
rect 283097 154730 283163 154733
rect 240182 154728 240291 154730
rect 240182 154672 240230 154728
rect 240286 154672 240291 154728
rect 240182 154667 240291 154672
rect 283054 154728 283163 154730
rect 283054 154672 283102 154728
rect 283158 154672 283163 154728
rect 283054 154667 283163 154672
rect 305177 154730 305243 154733
rect 309501 154730 309567 154733
rect 305177 154728 305378 154730
rect 305177 154672 305182 154728
rect 305238 154672 305378 154728
rect 305177 154670 305378 154672
rect 305177 154667 305243 154670
rect 240182 154597 240242 154667
rect 283054 154597 283114 154667
rect 234286 154532 234292 154596
rect 234356 154594 234362 154596
rect 234470 154594 234476 154596
rect 234356 154534 234476 154594
rect 234356 154532 234362 154534
rect 234470 154532 234476 154534
rect 234540 154532 234546 154596
rect 240182 154592 240291 154597
rect 240182 154536 240230 154592
rect 240286 154536 240291 154592
rect 240182 154534 240291 154536
rect 240225 154531 240291 154534
rect 266905 154594 266971 154597
rect 267089 154594 267155 154597
rect 266905 154592 267155 154594
rect 266905 154536 266910 154592
rect 266966 154536 267094 154592
rect 267150 154536 267155 154592
rect 266905 154534 267155 154536
rect 283054 154592 283163 154597
rect 283054 154536 283102 154592
rect 283158 154536 283163 154592
rect 283054 154534 283163 154536
rect 266905 154531 266971 154534
rect 267089 154531 267155 154534
rect 283097 154531 283163 154534
rect 305177 154594 305243 154597
rect 305318 154594 305378 154670
rect 305177 154592 305378 154594
rect 305177 154536 305182 154592
rect 305238 154536 305378 154592
rect 305177 154534 305378 154536
rect 309182 154728 309567 154730
rect 309182 154672 309506 154728
rect 309562 154672 309567 154728
rect 309182 154670 309567 154672
rect 309182 154594 309242 154670
rect 309501 154667 309567 154670
rect 392117 154730 392183 154733
rect 392117 154728 392226 154730
rect 392117 154672 392122 154728
rect 392178 154672 392226 154728
rect 392117 154667 392226 154672
rect 392166 154597 392226 154667
rect 309317 154594 309383 154597
rect 309182 154592 309383 154594
rect 309182 154536 309322 154592
rect 309378 154536 309383 154592
rect 309182 154534 309383 154536
rect 305177 154531 305243 154534
rect 309317 154531 309383 154534
rect 310697 154594 310763 154597
rect 310881 154594 310947 154597
rect 310697 154592 310947 154594
rect 310697 154536 310702 154592
rect 310758 154536 310886 154592
rect 310942 154536 310947 154592
rect 310697 154534 310947 154536
rect 310697 154531 310763 154534
rect 310881 154531 310947 154534
rect 331397 154594 331463 154597
rect 331581 154594 331647 154597
rect 331397 154592 331647 154594
rect 331397 154536 331402 154592
rect 331458 154536 331586 154592
rect 331642 154536 331647 154592
rect 331397 154534 331647 154536
rect 331397 154531 331463 154534
rect 331581 154531 331647 154534
rect 342345 154594 342411 154597
rect 342529 154594 342595 154597
rect 342345 154592 342595 154594
rect 342345 154536 342350 154592
rect 342406 154536 342534 154592
rect 342590 154536 342595 154592
rect 342345 154534 342595 154536
rect 342345 154531 342411 154534
rect 342529 154531 342595 154534
rect 386597 154594 386663 154597
rect 386781 154594 386847 154597
rect 386597 154592 386847 154594
rect 386597 154536 386602 154592
rect 386658 154536 386786 154592
rect 386842 154536 386847 154592
rect 386597 154534 386847 154536
rect 386597 154531 386663 154534
rect 386781 154531 386847 154534
rect 392117 154592 392226 154597
rect 392117 154536 392122 154592
rect 392178 154536 392226 154592
rect 392117 154534 392226 154536
rect 408401 154594 408467 154597
rect 408677 154594 408743 154597
rect 408401 154592 408743 154594
rect 408401 154536 408406 154592
rect 408462 154536 408682 154592
rect 408738 154536 408743 154592
rect 408401 154534 408743 154536
rect 392117 154531 392183 154534
rect 408401 154531 408467 154534
rect 408677 154531 408743 154534
rect 472157 154594 472223 154597
rect 472341 154594 472407 154597
rect 472157 154592 472407 154594
rect 472157 154536 472162 154592
rect 472218 154536 472346 154592
rect 472402 154536 472407 154592
rect 472157 154534 472407 154536
rect 472157 154531 472223 154534
rect 472341 154531 472407 154534
rect 252553 153234 252619 153237
rect 252829 153234 252895 153237
rect 252553 153232 252895 153234
rect 252553 153176 252558 153232
rect 252614 153176 252834 153232
rect 252890 153176 252895 153232
rect 252553 153174 252895 153176
rect 252553 153171 252619 153174
rect 252829 153171 252895 153174
rect 308213 153234 308279 153237
rect 308397 153234 308463 153237
rect 308213 153232 308463 153234
rect 308213 153176 308218 153232
rect 308274 153176 308402 153232
rect 308458 153176 308463 153232
rect 308213 153174 308463 153176
rect 308213 153171 308279 153174
rect 308397 153171 308463 153174
rect 327257 153234 327323 153237
rect 327441 153234 327507 153237
rect 327257 153232 327507 153234
rect 327257 153176 327262 153232
rect 327318 153176 327446 153232
rect 327502 153176 327507 153232
rect 327257 153174 327507 153176
rect 327257 153171 327323 153174
rect 327441 153171 327507 153174
rect 3325 151738 3391 151741
rect 258574 151738 258580 151740
rect 3325 151736 258580 151738
rect 3325 151680 3330 151736
rect 3386 151680 258580 151736
rect 3325 151678 258580 151680
rect 3325 151675 3391 151678
rect 258574 151676 258580 151678
rect 258644 151676 258650 151740
rect -960 150786 480 150876
rect 3325 150786 3391 150789
rect -960 150784 3391 150786
rect -960 150728 3330 150784
rect 3386 150728 3391 150784
rect -960 150726 3391 150728
rect -960 150636 480 150726
rect 3325 150723 3391 150726
rect 583520 146556 584960 146796
rect 266537 145074 266603 145077
rect 287237 145074 287303 145077
rect 305269 145074 305335 145077
rect 330109 145074 330175 145077
rect 266310 145072 266603 145074
rect 266310 145016 266542 145072
rect 266598 145016 266603 145072
rect 266310 145014 266603 145016
rect 234286 144876 234292 144940
rect 234356 144938 234362 144940
rect 234470 144938 234476 144940
rect 234356 144878 234476 144938
rect 234356 144876 234362 144878
rect 234470 144876 234476 144878
rect 234540 144876 234546 144940
rect 266310 144938 266370 145014
rect 266537 145011 266603 145014
rect 287102 145072 287303 145074
rect 287102 145016 287242 145072
rect 287298 145016 287303 145072
rect 287102 145014 287303 145016
rect 266445 144938 266511 144941
rect 266310 144936 266511 144938
rect 266310 144880 266450 144936
rect 266506 144880 266511 144936
rect 266310 144878 266511 144880
rect 287102 144938 287162 145014
rect 287237 145011 287303 145014
rect 304950 145072 305335 145074
rect 304950 145016 305274 145072
rect 305330 145016 305335 145072
rect 304950 145014 305335 145016
rect 287237 144938 287303 144941
rect 287102 144936 287303 144938
rect 287102 144880 287242 144936
rect 287298 144880 287303 144936
rect 287102 144878 287303 144880
rect 266445 144875 266511 144878
rect 287237 144875 287303 144878
rect 298277 144938 298343 144941
rect 298461 144938 298527 144941
rect 298277 144936 298527 144938
rect 298277 144880 298282 144936
rect 298338 144880 298466 144936
rect 298522 144880 298527 144936
rect 298277 144878 298527 144880
rect 304950 144938 305010 145014
rect 305269 145011 305335 145014
rect 329974 145072 330175 145074
rect 329974 145016 330114 145072
rect 330170 145016 330175 145072
rect 329974 145014 330175 145016
rect 329974 144941 330034 145014
rect 330109 145011 330175 145014
rect 305085 144938 305151 144941
rect 304950 144936 305151 144938
rect 304950 144880 305090 144936
rect 305146 144880 305151 144936
rect 304950 144878 305151 144880
rect 329974 144936 330083 144941
rect 356421 144938 356487 144941
rect 329974 144880 330022 144936
rect 330078 144880 330083 144936
rect 329974 144878 330083 144880
rect 298277 144875 298343 144878
rect 298461 144875 298527 144878
rect 305085 144875 305151 144878
rect 330017 144875 330083 144878
rect 356286 144936 356487 144938
rect 356286 144880 356426 144936
rect 356482 144880 356487 144936
rect 356286 144878 356487 144880
rect 356286 144802 356346 144878
rect 356421 144875 356487 144878
rect 357525 144938 357591 144941
rect 357709 144938 357775 144941
rect 357525 144936 357775 144938
rect 357525 144880 357530 144936
rect 357586 144880 357714 144936
rect 357770 144880 357775 144936
rect 357525 144878 357775 144880
rect 357525 144875 357591 144878
rect 357709 144875 357775 144878
rect 358997 144938 359063 144941
rect 359181 144938 359247 144941
rect 358997 144936 359247 144938
rect 358997 144880 359002 144936
rect 359058 144880 359186 144936
rect 359242 144880 359247 144936
rect 358997 144878 359247 144880
rect 358997 144875 359063 144878
rect 359181 144875 359247 144878
rect 356421 144802 356487 144805
rect 356286 144800 356487 144802
rect 356286 144744 356426 144800
rect 356482 144744 356487 144800
rect 356286 144742 356487 144744
rect 356421 144739 356487 144742
rect 240317 143578 240383 143581
rect 240501 143578 240567 143581
rect 240317 143576 240567 143578
rect 240317 143520 240322 143576
rect 240378 143520 240506 143576
rect 240562 143520 240567 143576
rect 240317 143518 240567 143520
rect 240317 143515 240383 143518
rect 240501 143515 240567 143518
rect 234337 138684 234403 138685
rect 234286 138682 234292 138684
rect 234246 138622 234292 138682
rect 234356 138680 234403 138684
rect 234398 138624 234403 138680
rect 234286 138620 234292 138622
rect 234356 138620 234403 138624
rect 234337 138619 234403 138620
rect 392209 138276 392275 138277
rect 392158 138274 392164 138276
rect 392118 138214 392164 138274
rect 392228 138272 392275 138276
rect 392270 138216 392275 138272
rect 392158 138212 392164 138214
rect 392228 138212 392275 138216
rect 392209 138211 392275 138212
rect -960 136370 480 136460
rect 3877 136370 3943 136373
rect -960 136368 3943 136370
rect -960 136312 3882 136368
rect 3938 136312 3943 136368
rect -960 136310 3943 136312
rect -960 136220 480 136310
rect 3877 136307 3943 136310
rect 244457 135418 244523 135421
rect 244414 135416 244523 135418
rect 244414 135360 244462 135416
rect 244518 135360 244523 135416
rect 244414 135355 244523 135360
rect 265157 135418 265223 135421
rect 324497 135418 324563 135421
rect 367369 135418 367435 135421
rect 386781 135418 386847 135421
rect 265157 135416 265266 135418
rect 265157 135360 265162 135416
rect 265218 135360 265266 135416
rect 265157 135355 265266 135360
rect 243077 135282 243143 135285
rect 243261 135282 243327 135285
rect 243077 135280 243327 135282
rect 243077 135224 243082 135280
rect 243138 135224 243266 135280
rect 243322 135224 243327 135280
rect 243077 135222 243327 135224
rect 243077 135219 243143 135222
rect 243261 135219 243327 135222
rect 244414 135149 244474 135355
rect 265206 135285 265266 135355
rect 324454 135416 324563 135418
rect 324454 135360 324502 135416
rect 324558 135360 324563 135416
rect 324454 135355 324563 135360
rect 367326 135416 367435 135418
rect 367326 135360 367374 135416
rect 367430 135360 367435 135416
rect 367326 135355 367435 135360
rect 386462 135416 386847 135418
rect 386462 135360 386786 135416
rect 386842 135360 386847 135416
rect 386462 135358 386847 135360
rect 324454 135285 324514 135355
rect 367326 135285 367386 135355
rect 265157 135280 265266 135285
rect 265157 135224 265162 135280
rect 265218 135224 265266 135280
rect 265157 135222 265266 135224
rect 270677 135282 270743 135285
rect 270861 135282 270927 135285
rect 270677 135280 270927 135282
rect 270677 135224 270682 135280
rect 270738 135224 270866 135280
rect 270922 135224 270927 135280
rect 270677 135222 270927 135224
rect 265157 135219 265223 135222
rect 270677 135219 270743 135222
rect 270861 135219 270927 135222
rect 295517 135282 295583 135285
rect 295701 135282 295767 135285
rect 295517 135280 295767 135282
rect 295517 135224 295522 135280
rect 295578 135224 295706 135280
rect 295762 135224 295767 135280
rect 295517 135222 295767 135224
rect 324454 135280 324563 135285
rect 324454 135224 324502 135280
rect 324558 135224 324563 135280
rect 324454 135222 324563 135224
rect 367326 135280 367435 135285
rect 367326 135224 367374 135280
rect 367430 135224 367435 135280
rect 367326 135222 367435 135224
rect 295517 135219 295583 135222
rect 295701 135219 295767 135222
rect 324497 135219 324563 135222
rect 367369 135219 367435 135222
rect 370037 135282 370103 135285
rect 370221 135282 370287 135285
rect 370037 135280 370287 135282
rect 370037 135224 370042 135280
rect 370098 135224 370226 135280
rect 370282 135224 370287 135280
rect 370037 135222 370287 135224
rect 386462 135282 386522 135358
rect 386781 135355 386847 135358
rect 386597 135282 386663 135285
rect 392117 135284 392183 135285
rect 392117 135282 392164 135284
rect 386462 135280 386663 135282
rect 386462 135224 386602 135280
rect 386658 135224 386663 135280
rect 386462 135222 386663 135224
rect 392072 135280 392164 135282
rect 392072 135224 392122 135280
rect 392072 135222 392164 135224
rect 370037 135219 370103 135222
rect 370221 135219 370287 135222
rect 386597 135219 386663 135222
rect 392117 135220 392164 135222
rect 392228 135220 392234 135284
rect 408861 135282 408927 135285
rect 409045 135282 409111 135285
rect 408861 135280 409111 135282
rect 408861 135224 408866 135280
rect 408922 135224 409050 135280
rect 409106 135224 409111 135280
rect 408861 135222 409111 135224
rect 392117 135219 392183 135220
rect 408861 135219 408927 135222
rect 409045 135219 409111 135222
rect 416773 135282 416839 135285
rect 416957 135282 417023 135285
rect 416773 135280 417023 135282
rect 416773 135224 416778 135280
rect 416834 135224 416962 135280
rect 417018 135224 417023 135280
rect 416773 135222 417023 135224
rect 416773 135219 416839 135222
rect 416957 135219 417023 135222
rect 427721 135282 427787 135285
rect 427905 135282 427971 135285
rect 427721 135280 427971 135282
rect 427721 135224 427726 135280
rect 427782 135224 427910 135280
rect 427966 135224 427971 135280
rect 427721 135222 427971 135224
rect 427721 135219 427787 135222
rect 427905 135219 427971 135222
rect 471973 135282 472039 135285
rect 472157 135282 472223 135285
rect 471973 135280 472223 135282
rect 471973 135224 471978 135280
rect 472034 135224 472162 135280
rect 472218 135224 472223 135280
rect 471973 135222 472223 135224
rect 471973 135219 472039 135222
rect 472157 135219 472223 135222
rect 244414 135144 244523 135149
rect 244414 135088 244462 135144
rect 244518 135088 244523 135144
rect 244414 135086 244523 135088
rect 244457 135083 244523 135086
rect 583520 134874 584960 134964
rect 583342 134814 584960 134874
rect 324262 134404 324268 134468
rect 324332 134466 324338 134468
rect 333881 134466 333947 134469
rect 324332 134464 333947 134466
rect 324332 134408 333886 134464
rect 333942 134408 333947 134464
rect 324332 134406 333947 134408
rect 324332 134404 324338 134406
rect 333881 134403 333947 134406
rect 402881 134330 402947 134333
rect 405641 134330 405707 134333
rect 417877 134330 417943 134333
rect 402881 134328 405707 134330
rect 402881 134272 402886 134328
rect 402942 134272 405646 134328
rect 405702 134272 405707 134328
rect 402881 134270 405707 134272
rect 402881 134267 402947 134270
rect 405641 134267 405707 134270
rect 415350 134328 417943 134330
rect 415350 134272 417882 134328
rect 417938 134272 417943 134328
rect 415350 134270 417943 134272
rect 267733 134194 267799 134197
rect 278681 134194 278747 134197
rect 267733 134192 278747 134194
rect 267733 134136 267738 134192
rect 267794 134136 278686 134192
rect 278742 134136 278747 134192
rect 267733 134134 278747 134136
rect 267733 134131 267799 134134
rect 278681 134131 278747 134134
rect 295241 134194 295307 134197
rect 298001 134194 298067 134197
rect 295241 134192 298067 134194
rect 295241 134136 295246 134192
rect 295302 134136 298006 134192
rect 298062 134136 298067 134192
rect 295241 134134 298067 134136
rect 295241 134131 295307 134134
rect 298001 134131 298067 134134
rect 301589 134194 301655 134197
rect 324262 134194 324268 134196
rect 301589 134192 306482 134194
rect 301589 134136 301594 134192
rect 301650 134136 306482 134192
rect 301589 134134 306482 134136
rect 301589 134131 301655 134134
rect 236361 134058 236427 134061
rect 267733 134058 267799 134061
rect 236318 134056 236427 134058
rect 236318 134000 236366 134056
rect 236422 134000 236427 134056
rect 236318 133995 236427 134000
rect 253798 134056 267799 134058
rect 253798 134000 267738 134056
rect 267794 134000 267799 134056
rect 253798 133998 267799 134000
rect 306422 134058 306482 134134
rect 323718 134134 324268 134194
rect 307569 134058 307635 134061
rect 306422 134056 307635 134058
rect 306422 134000 307574 134056
rect 307630 134000 307635 134056
rect 306422 133998 307635 134000
rect 236318 133925 236378 133995
rect 236269 133920 236378 133925
rect 236269 133864 236274 133920
rect 236330 133864 236378 133920
rect 236269 133862 236378 133864
rect 236269 133859 236335 133862
rect 249006 133860 249012 133924
rect 249076 133922 249082 133924
rect 253798 133922 253858 133998
rect 267733 133995 267799 133998
rect 307569 133995 307635 133998
rect 307753 134058 307819 134061
rect 318742 134058 318748 134060
rect 307753 134056 318748 134058
rect 307753 134000 307758 134056
rect 307814 134000 318748 134056
rect 307753 133998 318748 134000
rect 307753 133995 307819 133998
rect 318742 133996 318748 133998
rect 318812 133996 318818 134060
rect 249076 133862 253858 133922
rect 278681 133922 278747 133925
rect 285622 133922 285628 133924
rect 278681 133920 285628 133922
rect 278681 133864 278686 133920
rect 278742 133864 285628 133920
rect 278681 133862 285628 133864
rect 249076 133860 249082 133862
rect 278681 133859 278747 133862
rect 285622 133860 285628 133862
rect 285692 133860 285698 133924
rect 309501 133922 309567 133925
rect 309685 133922 309751 133925
rect 309501 133920 309751 133922
rect 309501 133864 309506 133920
rect 309562 133864 309690 133920
rect 309746 133864 309751 133920
rect 309501 133862 309751 133864
rect 309501 133859 309567 133862
rect 309685 133859 309751 133862
rect 318742 133724 318748 133788
rect 318812 133786 318818 133788
rect 323718 133786 323778 134134
rect 324262 134132 324268 134134
rect 324332 134132 324338 134196
rect 385217 134194 385283 134197
rect 393262 134194 393268 134196
rect 367142 134134 375482 134194
rect 333881 134058 333947 134061
rect 338021 134058 338087 134061
rect 333881 134056 338087 134058
rect 333881 134000 333886 134056
rect 333942 134000 338026 134056
rect 338082 134000 338087 134056
rect 333881 133998 338087 134000
rect 333881 133995 333947 133998
rect 338021 133995 338087 133998
rect 347957 134058 348023 134061
rect 353477 134058 353543 134061
rect 356421 134058 356487 134061
rect 347957 134056 348066 134058
rect 347957 134000 347962 134056
rect 348018 134000 348066 134056
rect 347957 133995 348066 134000
rect 353477 134056 353586 134058
rect 353477 134000 353482 134056
rect 353538 134000 353586 134056
rect 353477 133995 353586 134000
rect 356421 134056 356530 134058
rect 356421 134000 356426 134056
rect 356482 134000 356530 134056
rect 356421 133995 356530 134000
rect 348006 133925 348066 133995
rect 353526 133925 353586 133995
rect 356470 133925 356530 133995
rect 347957 133920 348066 133925
rect 347957 133864 347962 133920
rect 348018 133864 348066 133920
rect 347957 133862 348066 133864
rect 353477 133920 353586 133925
rect 353477 133864 353482 133920
rect 353538 133864 353586 133920
rect 353477 133862 353586 133864
rect 356421 133920 356530 133925
rect 356421 133864 356426 133920
rect 356482 133864 356530 133920
rect 356421 133862 356530 133864
rect 347957 133859 348023 133862
rect 353477 133859 353543 133862
rect 356421 133859 356487 133862
rect 357382 133860 357388 133924
rect 357452 133922 357458 133924
rect 367142 133922 367202 134134
rect 375422 134058 375482 134134
rect 385217 134192 393268 134194
rect 385217 134136 385222 134192
rect 385278 134136 393268 134192
rect 385217 134134 393268 134136
rect 385217 134131 385283 134134
rect 393262 134132 393268 134134
rect 393332 134132 393338 134196
rect 405733 134194 405799 134197
rect 415350 134194 415410 134270
rect 417877 134267 417943 134270
rect 492630 134270 502258 134330
rect 405733 134192 415410 134194
rect 405733 134136 405738 134192
rect 405794 134136 415410 134192
rect 405733 134134 415410 134136
rect 418245 134194 418311 134197
rect 418245 134192 427738 134194
rect 418245 134136 418250 134192
rect 418306 134136 427738 134192
rect 418245 134134 427738 134136
rect 405733 134131 405799 134134
rect 418245 134131 418311 134134
rect 383653 134058 383719 134061
rect 375422 134056 383719 134058
rect 375422 134000 383658 134056
rect 383714 134000 383719 134056
rect 375422 133998 383719 134000
rect 383653 133995 383719 133998
rect 357452 133862 367202 133922
rect 357452 133860 357458 133862
rect 393262 133860 393268 133924
rect 393332 133922 393338 133924
rect 402881 133922 402947 133925
rect 393332 133920 402947 133922
rect 393332 133864 402886 133920
rect 402942 133864 402947 133920
rect 393332 133862 402947 133864
rect 427678 133922 427738 134134
rect 427862 134134 437490 134194
rect 427862 133922 427922 134134
rect 427678 133862 427922 133922
rect 437430 133922 437490 134134
rect 456701 134058 456767 134061
rect 447182 134056 456767 134058
rect 447182 134000 456706 134056
rect 456762 134000 456767 134056
rect 447182 133998 456767 134000
rect 447182 133922 447242 133998
rect 456701 133995 456767 133998
rect 456885 134058 456951 134061
rect 473302 134058 473308 134060
rect 456885 134056 466378 134058
rect 456885 134000 456890 134056
rect 456946 134000 466378 134056
rect 456885 133998 466378 134000
rect 456885 133995 456951 133998
rect 437430 133862 447242 133922
rect 466318 133922 466378 133998
rect 466502 133998 473308 134058
rect 466502 133922 466562 133998
rect 473302 133996 473308 133998
rect 473372 133996 473378 134060
rect 492630 134058 492690 134270
rect 502198 134196 502258 134270
rect 531262 134268 531268 134332
rect 531332 134330 531338 134332
rect 540881 134330 540947 134333
rect 531332 134328 540947 134330
rect 531332 134272 540886 134328
rect 540942 134272 540947 134328
rect 531332 134270 540947 134272
rect 531332 134268 531338 134270
rect 540881 134267 540947 134270
rect 502190 134132 502196 134196
rect 502260 134132 502266 134196
rect 560201 134194 560267 134197
rect 560201 134192 563162 134194
rect 560201 134136 560206 134192
rect 560262 134136 563162 134192
rect 560201 134134 563162 134136
rect 560201 134131 560267 134134
rect 514569 134058 514635 134061
rect 485822 133998 492690 134058
rect 505142 134056 514635 134058
rect 505142 134000 514574 134056
rect 514630 134000 514635 134056
rect 505142 133998 514635 134000
rect 485822 133922 485882 133998
rect 466318 133862 466562 133922
rect 482878 133862 485882 133922
rect 393332 133860 393338 133862
rect 402881 133859 402947 133862
rect 318812 133726 323778 133786
rect 318812 133724 318818 133726
rect 285622 133588 285628 133652
rect 285692 133650 285698 133652
rect 295241 133650 295307 133653
rect 357382 133650 357388 133652
rect 285692 133648 295307 133650
rect 285692 133592 295246 133648
rect 295302 133592 295307 133648
rect 285692 133590 295307 133592
rect 285692 133588 285698 133590
rect 295241 133587 295307 133590
rect 348006 133590 357388 133650
rect 338113 133514 338179 133517
rect 348006 133514 348066 133590
rect 357382 133588 357388 133590
rect 357452 133588 357458 133652
rect 473302 133588 473308 133652
rect 473372 133650 473378 133652
rect 482878 133650 482938 133862
rect 502190 133860 502196 133924
rect 502260 133922 502266 133924
rect 505142 133922 505202 133998
rect 514569 133995 514635 133998
rect 526437 134058 526503 134061
rect 531262 134058 531268 134060
rect 526437 134056 531268 134058
rect 526437 134000 526442 134056
rect 526498 134000 531268 134056
rect 526437 133998 531268 134000
rect 526437 133995 526503 133998
rect 531262 133996 531268 133998
rect 531332 133996 531338 134060
rect 550582 134058 550588 134060
rect 543782 133998 550588 134058
rect 521653 133922 521719 133925
rect 502260 133862 505202 133922
rect 521518 133920 521719 133922
rect 521518 133864 521658 133920
rect 521714 133864 521719 133920
rect 521518 133862 521719 133864
rect 502260 133860 502266 133862
rect 473372 133590 482938 133650
rect 514569 133650 514635 133653
rect 521518 133650 521578 133862
rect 521653 133859 521719 133862
rect 540881 133922 540947 133925
rect 543782 133922 543842 133998
rect 550582 133996 550588 133998
rect 550652 133996 550658 134060
rect 540881 133920 543842 133922
rect 540881 133864 540886 133920
rect 540942 133864 543842 133920
rect 540881 133862 543842 133864
rect 563102 133922 563162 134134
rect 572621 134058 572687 134061
rect 583342 134058 583402 134814
rect 583520 134724 584960 134814
rect 569910 134056 572687 134058
rect 569910 134000 572626 134056
rect 572682 134000 572687 134056
rect 569910 133998 572687 134000
rect 569910 133922 569970 133998
rect 572621 133995 572687 133998
rect 576902 133998 583402 134058
rect 563102 133862 569970 133922
rect 572713 133922 572779 133925
rect 576902 133922 576962 133998
rect 572713 133920 576962 133922
rect 572713 133864 572718 133920
rect 572774 133864 576962 133920
rect 572713 133862 576962 133864
rect 540881 133859 540947 133862
rect 572713 133859 572779 133862
rect 550582 133724 550588 133788
rect 550652 133786 550658 133788
rect 560201 133786 560267 133789
rect 550652 133784 560267 133786
rect 550652 133728 560206 133784
rect 560262 133728 560267 133784
rect 550652 133726 560267 133728
rect 550652 133724 550658 133726
rect 560201 133723 560267 133726
rect 514569 133648 521578 133650
rect 514569 133592 514574 133648
rect 514630 133592 521578 133648
rect 514569 133590 521578 133592
rect 473372 133588 473378 133590
rect 514569 133587 514635 133590
rect 338113 133512 348066 133514
rect 338113 133456 338118 133512
rect 338174 133456 348066 133512
rect 338113 133454 348066 133456
rect 338113 133451 338179 133454
rect 249977 125900 250043 125901
rect 249926 125898 249932 125900
rect 249886 125838 249932 125898
rect 249996 125896 250043 125900
rect 250038 125840 250043 125896
rect 249926 125836 249932 125838
rect 249996 125836 250043 125840
rect 249977 125835 250043 125836
rect 283097 125762 283163 125765
rect 283054 125760 283163 125762
rect 283054 125704 283102 125760
rect 283158 125704 283163 125760
rect 283054 125699 283163 125704
rect 287237 125762 287303 125765
rect 288617 125762 288683 125765
rect 294137 125762 294203 125765
rect 287237 125760 287346 125762
rect 287237 125704 287242 125760
rect 287298 125704 287346 125760
rect 287237 125699 287346 125704
rect 283054 125629 283114 125699
rect 287286 125629 287346 125699
rect 249977 125628 250043 125629
rect 249926 125564 249932 125628
rect 249996 125626 250043 125628
rect 252921 125626 252987 125629
rect 249996 125624 250088 125626
rect 250038 125568 250088 125624
rect 249996 125566 250088 125568
rect 252694 125624 252987 125626
rect 252694 125568 252926 125624
rect 252982 125568 252987 125624
rect 252694 125566 252987 125568
rect 249996 125564 250043 125566
rect 249977 125563 250043 125564
rect 252553 125354 252619 125357
rect 252694 125354 252754 125566
rect 252921 125563 252987 125566
rect 271873 125626 271939 125629
rect 272057 125626 272123 125629
rect 271873 125624 272123 125626
rect 271873 125568 271878 125624
rect 271934 125568 272062 125624
rect 272118 125568 272123 125624
rect 271873 125566 272123 125568
rect 283054 125624 283163 125629
rect 283054 125568 283102 125624
rect 283158 125568 283163 125624
rect 283054 125566 283163 125568
rect 271873 125563 271939 125566
rect 272057 125563 272123 125566
rect 283097 125563 283163 125566
rect 287237 125624 287346 125629
rect 287237 125568 287242 125624
rect 287298 125568 287346 125624
rect 287237 125566 287346 125568
rect 288574 125760 288683 125762
rect 288574 125704 288622 125760
rect 288678 125704 288683 125760
rect 288574 125699 288683 125704
rect 294094 125760 294203 125762
rect 294094 125704 294142 125760
rect 294198 125704 294203 125760
rect 294094 125699 294203 125704
rect 324497 125760 324563 125765
rect 352097 125762 352163 125765
rect 357617 125762 357683 125765
rect 324497 125704 324502 125760
rect 324558 125704 324563 125760
rect 324497 125699 324563 125704
rect 352054 125760 352163 125762
rect 352054 125704 352102 125760
rect 352158 125704 352163 125760
rect 352054 125699 352163 125704
rect 357574 125760 357683 125762
rect 357574 125704 357622 125760
rect 357678 125704 357683 125760
rect 357574 125699 357683 125704
rect 393221 125762 393287 125765
rect 408861 125762 408927 125765
rect 393221 125760 393330 125762
rect 393221 125704 393226 125760
rect 393282 125704 393330 125760
rect 393221 125699 393330 125704
rect 288574 125629 288634 125699
rect 294094 125629 294154 125699
rect 324500 125629 324560 125699
rect 352054 125629 352114 125699
rect 288574 125624 288683 125629
rect 288574 125568 288622 125624
rect 288678 125568 288683 125624
rect 288574 125566 288683 125568
rect 287237 125563 287303 125566
rect 288617 125563 288683 125566
rect 294045 125624 294154 125629
rect 294045 125568 294050 125624
rect 294106 125568 294154 125624
rect 294045 125566 294154 125568
rect 324497 125624 324563 125629
rect 324497 125568 324502 125624
rect 324558 125568 324563 125624
rect 294045 125563 294111 125566
rect 324497 125563 324563 125568
rect 352005 125624 352114 125629
rect 352005 125568 352010 125624
rect 352066 125568 352114 125624
rect 352005 125566 352114 125568
rect 357574 125629 357634 125699
rect 393270 125629 393330 125699
rect 357574 125624 357683 125629
rect 357574 125568 357622 125624
rect 357678 125568 357683 125624
rect 357574 125566 357683 125568
rect 352005 125563 352071 125566
rect 357617 125563 357683 125566
rect 367369 125626 367435 125629
rect 367553 125626 367619 125629
rect 367369 125624 367619 125626
rect 367369 125568 367374 125624
rect 367430 125568 367558 125624
rect 367614 125568 367619 125624
rect 367369 125566 367619 125568
rect 367369 125563 367435 125566
rect 367553 125563 367619 125566
rect 393221 125624 393330 125629
rect 393221 125568 393226 125624
rect 393282 125568 393330 125624
rect 393221 125566 393330 125568
rect 408542 125760 408927 125762
rect 408542 125704 408866 125760
rect 408922 125704 408927 125760
rect 408542 125702 408927 125704
rect 408542 125626 408602 125702
rect 408861 125699 408927 125702
rect 408677 125626 408743 125629
rect 408542 125624 408743 125626
rect 408542 125568 408682 125624
rect 408738 125568 408743 125624
rect 408542 125566 408743 125568
rect 393221 125563 393287 125566
rect 408677 125563 408743 125566
rect 252553 125352 252754 125354
rect 252553 125296 252558 125352
rect 252614 125296 252754 125352
rect 252553 125294 252754 125296
rect 252553 125291 252619 125294
rect 359089 124266 359155 124269
rect 359046 124264 359155 124266
rect 359046 124208 359094 124264
rect 359150 124208 359155 124264
rect 359046 124203 359155 124208
rect 359046 124132 359106 124203
rect 359038 124068 359044 124132
rect 359108 124068 359114 124132
rect 365662 123388 365668 123452
rect 365732 123450 365738 123452
rect 365732 123390 375298 123450
rect 365732 123388 365738 123390
rect 307702 123252 307708 123316
rect 307772 123314 307778 123316
rect 344921 123314 344987 123317
rect 345933 123314 345999 123317
rect 307772 123254 322306 123314
rect 307772 123252 307778 123254
rect 252318 123116 252324 123180
rect 252388 123178 252394 123180
rect 322246 123178 322306 123254
rect 344921 123312 345999 123314
rect 344921 123256 344926 123312
rect 344982 123256 345938 123312
rect 345994 123256 345999 123312
rect 344921 123254 345999 123256
rect 375238 123314 375298 123390
rect 375238 123254 379714 123314
rect 344921 123251 344987 123254
rect 345933 123251 345999 123254
rect 335302 123178 335308 123180
rect 252388 123118 278698 123178
rect 252388 123116 252394 123118
rect 278638 123042 278698 123118
rect 292438 123118 302066 123178
rect 322246 123118 335308 123178
rect 292438 123042 292498 123118
rect 278638 122982 292498 123042
rect 302006 123042 302066 123118
rect 335302 123116 335308 123118
rect 335372 123116 335378 123180
rect 354581 123178 354647 123181
rect 354581 123176 360946 123178
rect 354581 123120 354586 123176
rect 354642 123120 360946 123176
rect 354581 123118 360946 123120
rect 354581 123115 354647 123118
rect 307702 123042 307708 123044
rect 302006 122982 307708 123042
rect 307702 122980 307708 122982
rect 307772 122980 307778 123044
rect 360886 123042 360946 123118
rect 365662 123042 365668 123044
rect 360886 122982 365668 123042
rect 365662 122980 365668 122982
rect 365732 122980 365738 123044
rect 379654 123042 379714 123254
rect 495206 123254 502258 123314
rect 434529 123178 434595 123181
rect 394006 123118 398850 123178
rect 394006 123042 394066 123118
rect 379654 122982 394066 123042
rect 335302 122844 335308 122908
rect 335372 122906 335378 122908
rect 344921 122906 344987 122909
rect 335372 122904 344987 122906
rect 335372 122848 344926 122904
rect 344982 122848 344987 122904
rect 335372 122846 344987 122848
rect 398790 122906 398850 123118
rect 434529 123176 437490 123178
rect 434529 123120 434534 123176
rect 434590 123120 437490 123176
rect 434529 123118 437490 123120
rect 434529 123115 434595 123118
rect 408542 122982 418170 123042
rect 408542 122906 408602 122982
rect 398790 122846 408602 122906
rect 418110 122906 418170 122982
rect 425053 122906 425119 122909
rect 418110 122904 425119 122906
rect 418110 122848 425058 122904
rect 425114 122848 425119 122904
rect 418110 122846 425119 122848
rect 437430 122906 437490 123118
rect 454033 123042 454099 123045
rect 447182 123040 454099 123042
rect 447182 122984 454038 123040
rect 454094 122984 454099 123040
rect 447182 122982 454099 122984
rect 447182 122906 447242 122982
rect 454033 122979 454099 122982
rect 458173 123042 458239 123045
rect 475929 123042 475995 123045
rect 458173 123040 463618 123042
rect 458173 122984 458178 123040
rect 458234 122984 463618 123040
rect 458173 122982 463618 122984
rect 458173 122979 458239 122982
rect 437430 122846 447242 122906
rect 463558 122906 463618 122982
rect 466502 123040 475995 123042
rect 466502 122984 475934 123040
rect 475990 122984 475995 123040
rect 466502 122982 475995 122984
rect 466502 122906 466562 122982
rect 475929 122979 475995 122982
rect 478137 123042 478203 123045
rect 495206 123042 495266 123254
rect 478137 123040 482938 123042
rect 478137 122984 478142 123040
rect 478198 122984 482938 123040
rect 478137 122982 482938 122984
rect 478137 122979 478203 122982
rect 463558 122846 466562 122906
rect 482878 122906 482938 122982
rect 485822 122982 495266 123042
rect 485822 122906 485882 122982
rect 482878 122846 485882 122906
rect 502198 122906 502258 123254
rect 531262 123252 531268 123316
rect 531332 123314 531338 123316
rect 540881 123314 540947 123317
rect 531332 123312 540947 123314
rect 531332 123256 540886 123312
rect 540942 123256 540947 123312
rect 531332 123254 540947 123256
rect 531332 123252 531338 123254
rect 540881 123251 540947 123254
rect 560201 123178 560267 123181
rect 583520 123178 584960 123268
rect 560201 123176 563162 123178
rect 560201 123120 560206 123176
rect 560262 123120 563162 123176
rect 560201 123118 563162 123120
rect 560201 123115 560267 123118
rect 514569 123042 514635 123045
rect 505142 123040 514635 123042
rect 505142 122984 514574 123040
rect 514630 122984 514635 123040
rect 505142 122982 514635 122984
rect 505142 122906 505202 122982
rect 514569 122979 514635 122982
rect 516869 123042 516935 123045
rect 526437 123042 526503 123045
rect 531262 123042 531268 123044
rect 516869 123040 521578 123042
rect 516869 122984 516874 123040
rect 516930 122984 521578 123040
rect 516869 122982 521578 122984
rect 516869 122979 516935 122982
rect 502198 122846 505202 122906
rect 521518 122906 521578 122982
rect 526437 123040 531268 123042
rect 526437 122984 526442 123040
rect 526498 122984 531268 123040
rect 526437 122982 531268 122984
rect 526437 122979 526503 122982
rect 531262 122980 531268 122982
rect 531332 122980 531338 123044
rect 550582 123042 550588 123044
rect 543782 122982 550588 123042
rect 524229 122906 524295 122909
rect 521518 122904 524295 122906
rect 521518 122848 524234 122904
rect 524290 122848 524295 122904
rect 521518 122846 524295 122848
rect 335372 122844 335378 122846
rect 344921 122843 344987 122846
rect 425053 122843 425119 122846
rect 524229 122843 524295 122846
rect 540881 122906 540947 122909
rect 543782 122906 543842 122982
rect 550582 122980 550588 122982
rect 550652 122980 550658 123044
rect 540881 122904 543842 122906
rect 540881 122848 540886 122904
rect 540942 122848 543842 122904
rect 540881 122846 543842 122848
rect 563102 122906 563162 123118
rect 583342 123118 584960 123178
rect 572621 123042 572687 123045
rect 583342 123042 583402 123118
rect 569910 123040 572687 123042
rect 569910 122984 572626 123040
rect 572682 122984 572687 123040
rect 569910 122982 572687 122984
rect 569910 122906 569970 122982
rect 572621 122979 572687 122982
rect 576902 122982 583402 123042
rect 583520 123028 584960 123118
rect 563102 122846 569970 122906
rect 572713 122906 572779 122909
rect 576902 122906 576962 122982
rect 572713 122904 576962 122906
rect 572713 122848 572718 122904
rect 572774 122848 576962 122904
rect 572713 122846 576962 122848
rect 540881 122843 540947 122846
rect 572713 122843 572779 122846
rect 550582 122708 550588 122772
rect 550652 122770 550658 122772
rect 560201 122770 560267 122773
rect 550652 122768 560267 122770
rect 550652 122712 560206 122768
rect 560262 122712 560267 122768
rect 550652 122710 560267 122712
rect 550652 122708 550658 122710
rect 560201 122707 560267 122710
rect -960 122090 480 122180
rect 2957 122090 3023 122093
rect -960 122088 3023 122090
rect -960 122032 2962 122088
rect 3018 122032 3023 122088
rect -960 122030 3023 122032
rect -960 121940 480 122030
rect 2957 122027 3023 122030
rect 234337 121818 234403 121821
rect 234337 121816 234538 121818
rect 234337 121760 234342 121816
rect 234398 121760 234538 121816
rect 234337 121758 234538 121760
rect 234337 121755 234403 121758
rect 234478 121684 234538 121758
rect 234470 121620 234476 121684
rect 234540 121620 234546 121684
rect 234705 121412 234771 121413
rect 234654 121410 234660 121412
rect 234614 121350 234660 121410
rect 234724 121408 234771 121412
rect 234766 121352 234771 121408
rect 234654 121348 234660 121350
rect 234724 121348 234771 121352
rect 234705 121347 234771 121348
rect 277577 116106 277643 116109
rect 277534 116104 277643 116106
rect 277534 116048 277582 116104
rect 277638 116048 277643 116104
rect 277534 116043 277643 116048
rect 277534 115973 277594 116043
rect 265065 115970 265131 115973
rect 265249 115970 265315 115973
rect 265065 115968 265315 115970
rect 265065 115912 265070 115968
rect 265126 115912 265254 115968
rect 265310 115912 265315 115968
rect 265065 115910 265315 115912
rect 265065 115907 265131 115910
rect 265249 115907 265315 115910
rect 277485 115968 277594 115973
rect 277485 115912 277490 115968
rect 277546 115912 277594 115968
rect 277485 115910 277594 115912
rect 304901 115970 304967 115973
rect 305085 115970 305151 115973
rect 304901 115968 305151 115970
rect 304901 115912 304906 115968
rect 304962 115912 305090 115968
rect 305146 115912 305151 115968
rect 304901 115910 305151 115912
rect 277485 115907 277551 115910
rect 304901 115907 304967 115910
rect 305085 115907 305151 115910
rect 397729 115970 397795 115973
rect 397913 115970 397979 115973
rect 397729 115968 397979 115970
rect 397729 115912 397734 115968
rect 397790 115912 397918 115968
rect 397974 115912 397979 115968
rect 397729 115910 397979 115912
rect 397729 115907 397795 115910
rect 397913 115907 397979 115910
rect 416773 115970 416839 115973
rect 416957 115970 417023 115973
rect 416773 115968 417023 115970
rect 416773 115912 416778 115968
rect 416834 115912 416962 115968
rect 417018 115912 417023 115968
rect 416773 115910 417023 115912
rect 416773 115907 416839 115910
rect 416957 115907 417023 115910
rect 471973 115970 472039 115973
rect 472157 115970 472223 115973
rect 471973 115968 472223 115970
rect 471973 115912 471978 115968
rect 472034 115912 472162 115968
rect 472218 115912 472223 115968
rect 471973 115910 472223 115912
rect 471973 115907 472039 115910
rect 472157 115907 472223 115910
rect 480253 115970 480319 115973
rect 480437 115970 480503 115973
rect 480253 115968 480503 115970
rect 480253 115912 480258 115968
rect 480314 115912 480442 115968
rect 480498 115912 480503 115968
rect 480253 115910 480503 115912
rect 480253 115907 480319 115910
rect 480437 115907 480503 115910
rect 319069 114610 319135 114613
rect 318934 114608 319135 114610
rect 318934 114552 319074 114608
rect 319130 114552 319135 114608
rect 318934 114550 319135 114552
rect 318934 114474 318994 114550
rect 319069 114547 319135 114550
rect 359038 114548 359044 114612
rect 359108 114548 359114 114612
rect 319069 114474 319135 114477
rect 353477 114474 353543 114477
rect 318934 114472 319135 114474
rect 318934 114416 319074 114472
rect 319130 114416 319135 114472
rect 318934 114414 319135 114416
rect 319069 114411 319135 114414
rect 353342 114472 353543 114474
rect 353342 114416 353482 114472
rect 353538 114416 353543 114472
rect 353342 114414 353543 114416
rect 359046 114474 359106 114548
rect 359181 114474 359247 114477
rect 359046 114472 359247 114474
rect 359046 114416 359186 114472
rect 359242 114416 359247 114472
rect 359046 114414 359247 114416
rect 353342 114338 353402 114414
rect 353477 114411 353543 114414
rect 359181 114411 359247 114414
rect 353569 114338 353635 114341
rect 353342 114336 353635 114338
rect 353342 114280 353574 114336
rect 353630 114280 353635 114336
rect 353342 114278 353635 114280
rect 353569 114275 353635 114278
rect 234705 112980 234771 112981
rect 234654 112916 234660 112980
rect 234724 112978 234771 112980
rect 234724 112976 234816 112978
rect 234766 112920 234816 112976
rect 234724 112918 234816 112920
rect 234724 112916 234771 112918
rect 234705 112915 234771 112916
rect 583520 111482 584960 111572
rect 583342 111422 584960 111482
rect 327022 111012 327028 111076
rect 327092 111074 327098 111076
rect 327092 111014 336658 111074
rect 327092 111012 327098 111014
rect 278773 110938 278839 110941
rect 269070 110936 278839 110938
rect 269070 110880 278778 110936
rect 278834 110880 278839 110936
rect 269070 110878 278839 110880
rect 247534 110604 247540 110668
rect 247604 110666 247610 110668
rect 269070 110666 269130 110878
rect 278773 110875 278839 110878
rect 298001 110802 298067 110805
rect 327022 110802 327028 110804
rect 298001 110800 298202 110802
rect 298001 110744 298006 110800
rect 298062 110744 298202 110800
rect 298001 110742 298202 110744
rect 298001 110739 298067 110742
rect 298142 110668 298202 110742
rect 311758 110742 327028 110802
rect 247604 110606 269130 110666
rect 247604 110604 247610 110606
rect 298134 110604 298140 110668
rect 298204 110604 298210 110668
rect 278773 110530 278839 110533
rect 298001 110530 298067 110533
rect 278773 110528 298067 110530
rect 278773 110472 278778 110528
rect 278834 110472 298006 110528
rect 298062 110472 298067 110528
rect 278773 110470 298067 110472
rect 278773 110467 278839 110470
rect 298001 110467 298067 110470
rect 298134 110468 298140 110532
rect 298204 110530 298210 110532
rect 311758 110530 311818 110742
rect 327022 110740 327028 110742
rect 327092 110740 327098 110804
rect 336598 110802 336658 111014
rect 463366 110938 463372 110940
rect 456566 110878 463372 110938
rect 336733 110802 336799 110805
rect 357382 110802 357388 110804
rect 336598 110800 336799 110802
rect 336598 110744 336738 110800
rect 336794 110744 336799 110800
rect 336598 110742 336799 110744
rect 336733 110739 336799 110742
rect 351134 110742 357388 110802
rect 298204 110470 311818 110530
rect 346209 110530 346275 110533
rect 351134 110530 351194 110742
rect 357382 110740 357388 110742
rect 357452 110740 357458 110804
rect 434529 110802 434595 110805
rect 394006 110742 398850 110802
rect 394006 110666 394066 110742
rect 367326 110606 394066 110666
rect 346209 110528 351194 110530
rect 346209 110472 346214 110528
rect 346270 110472 351194 110528
rect 346209 110470 351194 110472
rect 298204 110468 298210 110470
rect 346209 110467 346275 110470
rect 357566 110468 357572 110532
rect 357636 110530 357642 110532
rect 367326 110530 367386 110606
rect 357636 110470 367386 110530
rect 398790 110530 398850 110742
rect 434529 110800 437490 110802
rect 434529 110744 434534 110800
rect 434590 110744 437490 110800
rect 434529 110742 437490 110744
rect 434529 110739 434595 110742
rect 418061 110666 418127 110669
rect 408542 110664 418127 110666
rect 408542 110608 418066 110664
rect 418122 110608 418127 110664
rect 408542 110606 418127 110608
rect 408542 110530 408602 110606
rect 418061 110603 418127 110606
rect 425053 110530 425119 110533
rect 398790 110470 408602 110530
rect 424918 110528 425119 110530
rect 424918 110472 425058 110528
rect 425114 110472 425119 110528
rect 424918 110470 425119 110472
rect 437430 110530 437490 110742
rect 456566 110666 456626 110878
rect 463366 110876 463372 110878
rect 463436 110876 463442 110940
rect 502006 110938 502012 110940
rect 495206 110878 502012 110938
rect 495206 110666 495266 110878
rect 502006 110876 502012 110878
rect 502076 110876 502082 110940
rect 531262 110876 531268 110940
rect 531332 110938 531338 110940
rect 540881 110938 540947 110941
rect 531332 110936 540947 110938
rect 531332 110880 540886 110936
rect 540942 110880 540947 110936
rect 531332 110878 540947 110880
rect 531332 110876 531338 110878
rect 540881 110875 540947 110878
rect 560201 110802 560267 110805
rect 560201 110800 563162 110802
rect 560201 110744 560206 110800
rect 560262 110744 563162 110800
rect 560201 110742 563162 110744
rect 560201 110739 560267 110742
rect 514569 110666 514635 110669
rect 447182 110606 456626 110666
rect 466502 110606 475946 110666
rect 447182 110530 447242 110606
rect 437430 110470 447242 110530
rect 357636 110468 357642 110470
rect 418061 110258 418127 110261
rect 424918 110258 424978 110470
rect 425053 110467 425119 110470
rect 463550 110468 463556 110532
rect 463620 110530 463626 110532
rect 466502 110530 466562 110606
rect 463620 110470 466562 110530
rect 475886 110530 475946 110606
rect 485822 110606 495266 110666
rect 505142 110664 514635 110666
rect 505142 110608 514574 110664
rect 514630 110608 514635 110664
rect 505142 110606 514635 110608
rect 485822 110530 485882 110606
rect 475886 110470 485882 110530
rect 463620 110468 463626 110470
rect 502190 110468 502196 110532
rect 502260 110530 502266 110532
rect 505142 110530 505202 110606
rect 514569 110603 514635 110606
rect 526437 110666 526503 110669
rect 531262 110666 531268 110668
rect 526437 110664 531268 110666
rect 526437 110608 526442 110664
rect 526498 110608 531268 110664
rect 526437 110606 531268 110608
rect 526437 110603 526503 110606
rect 531262 110604 531268 110606
rect 531332 110604 531338 110668
rect 550582 110666 550588 110668
rect 543782 110606 550588 110666
rect 521653 110530 521719 110533
rect 502260 110470 505202 110530
rect 521518 110528 521719 110530
rect 521518 110472 521658 110528
rect 521714 110472 521719 110528
rect 521518 110470 521719 110472
rect 502260 110468 502266 110470
rect 418061 110256 424978 110258
rect 418061 110200 418066 110256
rect 418122 110200 424978 110256
rect 418061 110198 424978 110200
rect 514569 110258 514635 110261
rect 521518 110258 521578 110470
rect 521653 110467 521719 110470
rect 540881 110530 540947 110533
rect 543782 110530 543842 110606
rect 550582 110604 550588 110606
rect 550652 110604 550658 110668
rect 540881 110528 543842 110530
rect 540881 110472 540886 110528
rect 540942 110472 543842 110528
rect 540881 110470 543842 110472
rect 563102 110530 563162 110742
rect 572621 110666 572687 110669
rect 583342 110666 583402 111422
rect 583520 111332 584960 111422
rect 569910 110664 572687 110666
rect 569910 110608 572626 110664
rect 572682 110608 572687 110664
rect 569910 110606 572687 110608
rect 569910 110530 569970 110606
rect 572621 110603 572687 110606
rect 576902 110606 583402 110666
rect 563102 110470 569970 110530
rect 572713 110530 572779 110533
rect 576902 110530 576962 110606
rect 572713 110528 576962 110530
rect 572713 110472 572718 110528
rect 572774 110472 576962 110528
rect 572713 110470 576962 110472
rect 540881 110467 540947 110470
rect 572713 110467 572779 110470
rect 550582 110332 550588 110396
rect 550652 110394 550658 110396
rect 560201 110394 560267 110397
rect 550652 110392 560267 110394
rect 550652 110336 560206 110392
rect 560262 110336 560267 110392
rect 550652 110334 560267 110336
rect 550652 110332 550658 110334
rect 560201 110331 560267 110334
rect 514569 110256 521578 110258
rect 514569 110200 514574 110256
rect 514630 110200 521578 110256
rect 514569 110198 521578 110200
rect 418061 110195 418127 110198
rect 514569 110195 514635 110198
rect -960 107674 480 107764
rect 3785 107674 3851 107677
rect -960 107672 3851 107674
rect -960 107616 3790 107672
rect 3846 107616 3851 107672
rect -960 107614 3851 107616
rect -960 107524 480 107614
rect 3785 107611 3851 107614
rect 281625 106314 281691 106317
rect 281809 106314 281875 106317
rect 281625 106312 281875 106314
rect 281625 106256 281630 106312
rect 281686 106256 281814 106312
rect 281870 106256 281875 106312
rect 281625 106254 281875 106256
rect 281625 106251 281691 106254
rect 281809 106251 281875 106254
rect 305177 106280 305243 106283
rect 305177 106278 305378 106280
rect 305177 106222 305182 106278
rect 305238 106222 305378 106278
rect 305177 106220 305378 106222
rect 305177 106217 305243 106220
rect 305318 106045 305378 106220
rect 305269 106040 305378 106045
rect 305269 105984 305274 106040
rect 305330 105984 305378 106040
rect 305269 105982 305378 105984
rect 305269 105979 305335 105982
rect 351821 104818 351887 104821
rect 352005 104818 352071 104821
rect 351821 104816 352071 104818
rect 351821 104760 351826 104816
rect 351882 104760 352010 104816
rect 352066 104760 352071 104816
rect 351821 104758 352071 104760
rect 351821 104755 351887 104758
rect 352005 104755 352071 104758
rect 583520 99636 584960 99876
rect 451641 99516 451707 99517
rect 451590 99514 451596 99516
rect 451550 99454 451596 99514
rect 451660 99512 451707 99516
rect 451702 99456 451707 99512
rect 451590 99452 451596 99454
rect 451660 99452 451707 99456
rect 451641 99451 451707 99452
rect 234286 96596 234292 96660
rect 234356 96658 234362 96660
rect 234470 96658 234476 96660
rect 234356 96598 234476 96658
rect 234356 96596 234362 96598
rect 234470 96596 234476 96598
rect 234540 96596 234546 96660
rect 241789 96658 241855 96661
rect 241973 96658 242039 96661
rect 241789 96656 242039 96658
rect 241789 96600 241794 96656
rect 241850 96600 241978 96656
rect 242034 96600 242039 96656
rect 241789 96598 242039 96600
rect 241789 96595 241855 96598
rect 241973 96595 242039 96598
rect 388069 96658 388135 96661
rect 392025 96658 392091 96661
rect 392209 96658 392275 96661
rect 388069 96656 388178 96658
rect 388069 96600 388074 96656
rect 388130 96600 388178 96656
rect 388069 96595 388178 96600
rect 392025 96656 392275 96658
rect 392025 96600 392030 96656
rect 392086 96600 392214 96656
rect 392270 96600 392275 96656
rect 392025 96598 392275 96600
rect 392025 96595 392091 96598
rect 392209 96595 392275 96598
rect 416773 96658 416839 96661
rect 416957 96658 417023 96661
rect 451641 96660 451707 96661
rect 416773 96656 417023 96658
rect 416773 96600 416778 96656
rect 416834 96600 416962 96656
rect 417018 96600 417023 96656
rect 416773 96598 417023 96600
rect 416773 96595 416839 96598
rect 416957 96595 417023 96598
rect 451590 96596 451596 96660
rect 451660 96658 451707 96660
rect 471973 96658 472039 96661
rect 472157 96658 472223 96661
rect 451660 96656 451752 96658
rect 451702 96600 451752 96656
rect 451660 96598 451752 96600
rect 471973 96656 472223 96658
rect 471973 96600 471978 96656
rect 472034 96600 472162 96656
rect 472218 96600 472223 96656
rect 471973 96598 472223 96600
rect 451660 96596 451707 96598
rect 451641 96595 451707 96596
rect 471973 96595 472039 96598
rect 472157 96595 472223 96598
rect 387977 96522 388043 96525
rect 388118 96522 388178 96595
rect 387977 96520 388178 96522
rect 387977 96464 387982 96520
rect 388038 96464 388178 96520
rect 387977 96462 388178 96464
rect 387977 96459 388043 96462
rect 270769 95434 270835 95437
rect 270542 95432 270835 95434
rect 270542 95376 270774 95432
rect 270830 95376 270835 95432
rect 270542 95374 270835 95376
rect 270542 95298 270602 95374
rect 270769 95371 270835 95374
rect 270677 95298 270743 95301
rect 270542 95296 270743 95298
rect 270542 95240 270682 95296
rect 270738 95240 270743 95296
rect 270542 95238 270743 95240
rect 270677 95235 270743 95238
rect 356421 94072 356487 94077
rect 356421 94016 356426 94072
rect 356482 94016 356487 94072
rect 356421 94011 356487 94016
rect 356424 93941 356484 94011
rect 356421 93936 356487 93941
rect 356421 93880 356426 93936
rect 356482 93880 356487 93936
rect 356421 93875 356487 93880
rect -960 93258 480 93348
rect 3693 93258 3759 93261
rect -960 93256 3759 93258
rect -960 93200 3698 93256
rect 3754 93200 3759 93256
rect -960 93198 3759 93200
rect -960 93108 480 93198
rect 3693 93195 3759 93198
rect 234470 89858 234476 89860
rect 234294 89798 234476 89858
rect 234294 89588 234354 89798
rect 234470 89796 234476 89798
rect 234540 89796 234546 89860
rect 234286 89524 234292 89588
rect 234356 89524 234362 89588
rect 583520 87954 584960 88044
rect 583342 87894 584960 87954
rect 550582 87484 550588 87548
rect 550652 87546 550658 87548
rect 560201 87546 560267 87549
rect 550652 87544 560267 87546
rect 550652 87488 560206 87544
rect 560262 87488 560267 87544
rect 550652 87486 560267 87488
rect 550652 87484 550658 87486
rect 560201 87483 560267 87486
rect 299422 87410 299428 87412
rect 292254 87350 299428 87410
rect 242750 87076 242756 87140
rect 242820 87138 242826 87140
rect 259361 87138 259427 87141
rect 267733 87138 267799 87141
rect 242820 87078 248522 87138
rect 242820 87076 242826 87078
rect 248462 87002 248522 87078
rect 259361 87136 267799 87138
rect 259361 87080 259366 87136
rect 259422 87080 267738 87136
rect 267794 87080 267799 87136
rect 259361 87078 267799 87080
rect 259361 87075 259427 87078
rect 267733 87075 267799 87078
rect 273713 87138 273779 87141
rect 292254 87138 292314 87350
rect 299422 87348 299428 87350
rect 299492 87348 299498 87412
rect 317454 87348 317460 87412
rect 317524 87410 317530 87412
rect 321461 87410 321527 87413
rect 536097 87410 536163 87413
rect 317524 87408 321527 87410
rect 317524 87352 321466 87408
rect 321522 87352 321527 87408
rect 317524 87350 321527 87352
rect 317524 87348 317530 87350
rect 321461 87347 321527 87350
rect 456566 87350 463618 87410
rect 338021 87274 338087 87277
rect 340781 87274 340847 87277
rect 338021 87272 340847 87274
rect 338021 87216 338026 87272
rect 338082 87216 340786 87272
rect 340842 87216 340847 87272
rect 338021 87214 340847 87216
rect 338021 87211 338087 87214
rect 340781 87211 340847 87214
rect 354581 87274 354647 87277
rect 365621 87274 365687 87277
rect 384941 87276 385007 87277
rect 384941 87274 384988 87276
rect 354581 87272 365687 87274
rect 354581 87216 354586 87272
rect 354642 87216 365626 87272
rect 365682 87216 365687 87272
rect 354581 87214 365687 87216
rect 384900 87272 384988 87274
rect 384900 87216 384946 87272
rect 384900 87214 384988 87216
rect 354581 87211 354647 87214
rect 365621 87211 365687 87214
rect 384941 87212 384988 87214
rect 385052 87212 385058 87276
rect 385166 87212 385172 87276
rect 385236 87274 385242 87276
rect 434529 87274 434595 87277
rect 385236 87214 398850 87274
rect 385236 87212 385242 87214
rect 384941 87211 385007 87212
rect 273713 87136 292314 87138
rect 273713 87080 273718 87136
rect 273774 87080 292314 87136
rect 273713 87078 292314 87080
rect 273713 87075 273779 87078
rect 299422 87076 299428 87140
rect 299492 87138 299498 87140
rect 317454 87138 317460 87140
rect 299492 87078 317460 87138
rect 299492 87076 299498 87078
rect 317454 87076 317460 87078
rect 317524 87076 317530 87140
rect 321461 87138 321527 87141
rect 328545 87138 328611 87141
rect 321461 87136 328611 87138
rect 321461 87080 321466 87136
rect 321522 87080 328550 87136
rect 328606 87080 328611 87136
rect 321461 87078 328611 87080
rect 321461 87075 321527 87078
rect 328545 87075 328611 87078
rect 373901 87138 373967 87141
rect 375414 87138 375420 87140
rect 373901 87136 375420 87138
rect 373901 87080 373906 87136
rect 373962 87080 375420 87136
rect 373901 87078 375420 87080
rect 373901 87075 373967 87078
rect 375414 87076 375420 87078
rect 375484 87076 375490 87140
rect 257981 87002 258047 87005
rect 248462 87000 258047 87002
rect 248462 86944 257986 87000
rect 258042 86944 258047 87000
rect 248462 86942 258047 86944
rect 257981 86939 258047 86942
rect 357525 87002 357591 87005
rect 357709 87002 357775 87005
rect 357525 87000 357775 87002
rect 357525 86944 357530 87000
rect 357586 86944 357714 87000
rect 357770 86944 357775 87000
rect 357525 86942 357775 86944
rect 398790 87002 398850 87214
rect 434529 87272 437490 87274
rect 434529 87216 434534 87272
rect 434590 87216 437490 87272
rect 434529 87214 437490 87216
rect 434529 87211 434595 87214
rect 415393 87138 415459 87141
rect 408542 87136 415459 87138
rect 408542 87080 415398 87136
rect 415454 87080 415459 87136
rect 408542 87078 415459 87080
rect 408542 87002 408602 87078
rect 415393 87075 415459 87078
rect 398790 86942 408602 87002
rect 424869 87002 424935 87005
rect 425053 87002 425119 87005
rect 424869 87000 425119 87002
rect 424869 86944 424874 87000
rect 424930 86944 425058 87000
rect 425114 86944 425119 87000
rect 424869 86942 425119 86944
rect 437430 87002 437490 87214
rect 456566 87138 456626 87350
rect 463558 87276 463618 87350
rect 492630 87350 502258 87410
rect 463550 87212 463556 87276
rect 463620 87212 463626 87276
rect 475929 87138 475995 87141
rect 447182 87078 456626 87138
rect 466502 87136 475995 87138
rect 466502 87080 475934 87136
rect 475990 87080 475995 87136
rect 466502 87078 475995 87080
rect 447182 87002 447242 87078
rect 437430 86942 447242 87002
rect 357525 86939 357591 86942
rect 357709 86939 357775 86942
rect 424869 86939 424935 86942
rect 425053 86939 425119 86942
rect 463550 86940 463556 87004
rect 463620 87002 463626 87004
rect 466502 87002 466562 87078
rect 475929 87075 475995 87078
rect 476113 87138 476179 87141
rect 492630 87138 492690 87350
rect 502198 87276 502258 87350
rect 531270 87408 536163 87410
rect 531270 87352 536102 87408
rect 536158 87352 536163 87408
rect 531270 87350 536163 87352
rect 502190 87212 502196 87276
rect 502260 87212 502266 87276
rect 531270 87138 531330 87350
rect 536097 87347 536163 87350
rect 560201 87274 560267 87277
rect 560201 87272 563162 87274
rect 560201 87216 560206 87272
rect 560262 87216 563162 87272
rect 560201 87214 563162 87216
rect 560201 87211 560267 87214
rect 550582 87138 550588 87140
rect 476113 87136 482938 87138
rect 476113 87080 476118 87136
rect 476174 87080 482938 87136
rect 476113 87078 482938 87080
rect 476113 87075 476179 87078
rect 463620 86942 466562 87002
rect 482878 87002 482938 87078
rect 485822 87078 492690 87138
rect 505142 87078 516794 87138
rect 485822 87002 485882 87078
rect 482878 86942 485882 87002
rect 463620 86940 463626 86942
rect 502190 86940 502196 87004
rect 502260 87002 502266 87004
rect 505142 87002 505202 87078
rect 502260 86942 505202 87002
rect 516734 87002 516794 87078
rect 529798 87078 531330 87138
rect 543782 87078 550588 87138
rect 520222 87002 520228 87004
rect 516734 86942 520228 87002
rect 502260 86940 502266 86942
rect 520222 86940 520228 86942
rect 520292 86940 520298 87004
rect 525057 87002 525123 87005
rect 529798 87002 529858 87078
rect 525057 87000 529858 87002
rect 525057 86944 525062 87000
rect 525118 86944 529858 87000
rect 525057 86942 529858 86944
rect 536097 87002 536163 87005
rect 543782 87002 543842 87078
rect 550582 87076 550588 87078
rect 550652 87076 550658 87140
rect 536097 87000 543842 87002
rect 536097 86944 536102 87000
rect 536158 86944 543842 87000
rect 536097 86942 543842 86944
rect 563102 87002 563162 87214
rect 572621 87138 572687 87141
rect 569910 87136 572687 87138
rect 569910 87080 572626 87136
rect 572682 87080 572687 87136
rect 569910 87078 572687 87080
rect 569910 87002 569970 87078
rect 572621 87075 572687 87078
rect 576761 87138 576827 87141
rect 583342 87138 583402 87894
rect 583520 87804 584960 87894
rect 576761 87136 583402 87138
rect 576761 87080 576766 87136
rect 576822 87080 583402 87136
rect 576761 87078 583402 87080
rect 576761 87075 576827 87078
rect 563102 86942 569970 87002
rect 525057 86939 525123 86942
rect 536097 86939 536163 86942
rect 257981 86866 258047 86869
rect 259361 86866 259427 86869
rect 257981 86864 259427 86866
rect 257981 86808 257986 86864
rect 258042 86808 259366 86864
rect 259422 86808 259427 86864
rect 257981 86806 259427 86808
rect 257981 86803 258047 86806
rect 259361 86803 259427 86806
rect 375414 86804 375420 86868
rect 375484 86866 375490 86868
rect 384941 86866 385007 86869
rect 375484 86864 385007 86866
rect 375484 86808 384946 86864
rect 385002 86808 385007 86864
rect 375484 86806 385007 86808
rect 375484 86804 375490 86806
rect 384941 86803 385007 86806
rect 520222 86668 520228 86732
rect 520292 86730 520298 86732
rect 525057 86730 525123 86733
rect 520292 86728 525123 86730
rect 520292 86672 525062 86728
rect 525118 86672 525123 86728
rect 520292 86670 525123 86672
rect 520292 86668 520298 86670
rect 525057 86667 525123 86670
rect 266445 82786 266511 82789
rect 266310 82784 266511 82786
rect 266310 82728 266450 82784
rect 266506 82728 266511 82784
rect 266310 82726 266511 82728
rect 266310 82650 266370 82726
rect 266445 82723 266511 82726
rect 266629 82650 266695 82653
rect 266310 82648 266695 82650
rect 266310 82592 266634 82648
rect 266690 82592 266695 82648
rect 266310 82590 266695 82592
rect 266629 82587 266695 82590
rect 234286 80684 234292 80748
rect 234356 80746 234362 80748
rect 234654 80746 234660 80748
rect 234356 80686 234660 80746
rect 234356 80684 234362 80686
rect 234654 80684 234660 80686
rect 234724 80684 234730 80748
rect -960 78978 480 79068
rect 3325 78978 3391 78981
rect -960 78976 3391 78978
rect -960 78920 3330 78976
rect 3386 78920 3391 78976
rect -960 78918 3391 78920
rect -960 78828 480 78918
rect 3325 78915 3391 78918
rect 253105 76530 253171 76533
rect 253105 76528 258090 76530
rect 253105 76472 253110 76528
rect 253166 76472 258090 76528
rect 253105 76470 258090 76472
rect 253105 76467 253171 76470
rect 258030 76394 258090 76470
rect 258030 76334 263794 76394
rect 263734 76122 263794 76334
rect 318934 76334 341442 76394
rect 309041 76258 309107 76261
rect 304214 76256 309107 76258
rect 304214 76200 309046 76256
rect 309102 76200 309107 76256
rect 304214 76198 309107 76200
rect 263734 76062 273362 76122
rect 244038 75924 244044 75988
rect 244108 75986 244114 75988
rect 253105 75986 253171 75989
rect 244108 75984 253171 75986
rect 244108 75928 253110 75984
rect 253166 75928 253171 75984
rect 244108 75926 253171 75928
rect 273302 75986 273362 76062
rect 283465 75986 283531 75989
rect 273302 75984 283531 75986
rect 273302 75928 283470 75984
rect 283526 75928 283531 75984
rect 273302 75926 283531 75928
rect 244108 75924 244114 75926
rect 253105 75923 253171 75926
rect 283465 75923 283531 75926
rect 298277 75986 298343 75989
rect 298553 75986 298619 75989
rect 298277 75984 298619 75986
rect 298277 75928 298282 75984
rect 298338 75928 298558 75984
rect 298614 75928 298619 75984
rect 298277 75926 298619 75928
rect 298277 75923 298343 75926
rect 298553 75923 298619 75926
rect 234470 75788 234476 75852
rect 234540 75850 234546 75852
rect 234654 75850 234660 75852
rect 234540 75790 234660 75850
rect 234540 75788 234546 75790
rect 234654 75788 234660 75790
rect 234724 75788 234730 75852
rect 290549 75850 290615 75853
rect 304214 75850 304274 76198
rect 309041 76195 309107 76198
rect 317321 76258 317387 76261
rect 318701 76258 318767 76261
rect 318934 76258 318994 76334
rect 317321 76256 318994 76258
rect 317321 76200 317326 76256
rect 317382 76200 318706 76256
rect 318762 76200 318994 76256
rect 317321 76198 318994 76200
rect 317321 76195 317387 76198
rect 318701 76195 318810 76198
rect 318750 76125 318810 76195
rect 318701 76120 318810 76125
rect 318701 76064 318706 76120
rect 318762 76064 318810 76120
rect 318701 76062 318810 76064
rect 341382 76122 341442 76334
rect 357382 76332 357388 76396
rect 357452 76394 357458 76396
rect 357452 76334 370514 76394
rect 357452 76332 357458 76334
rect 357382 76122 357388 76124
rect 341382 76062 343098 76122
rect 318701 76059 318767 76062
rect 343038 75986 343098 76062
rect 350582 76062 357388 76122
rect 343038 75952 350458 75986
rect 350582 75952 350642 76062
rect 357382 76060 357388 76062
rect 357452 76060 357458 76124
rect 370454 76122 370514 76334
rect 425102 76334 427738 76394
rect 398741 76258 398807 76261
rect 389222 76256 398807 76258
rect 389222 76200 398746 76256
rect 398802 76200 398807 76256
rect 389222 76198 398807 76200
rect 376702 76122 376708 76124
rect 370454 76062 376708 76122
rect 376702 76060 376708 76062
rect 376772 76060 376778 76124
rect 376886 76060 376892 76124
rect 376956 76122 376962 76124
rect 389222 76122 389282 76198
rect 398741 76195 398807 76198
rect 405641 76258 405707 76261
rect 418061 76258 418127 76261
rect 425102 76258 425162 76334
rect 405641 76256 408418 76258
rect 405641 76200 405646 76256
rect 405702 76200 408418 76256
rect 405641 76198 408418 76200
rect 405641 76195 405707 76198
rect 376956 76062 389282 76122
rect 376956 76060 376962 76062
rect 343038 75926 350642 75952
rect 408358 75986 408418 76198
rect 415350 76256 418127 76258
rect 415350 76200 418066 76256
rect 418122 76200 418127 76256
rect 415350 76198 418127 76200
rect 415350 76122 415410 76198
rect 418061 76195 418127 76198
rect 424918 76198 425162 76258
rect 427678 76258 427738 76334
rect 495206 76334 502258 76394
rect 427678 76198 437490 76258
rect 408542 76062 415410 76122
rect 418153 76122 418219 76125
rect 424918 76122 424978 76198
rect 418153 76120 424978 76122
rect 418153 76064 418158 76120
rect 418214 76064 424978 76120
rect 418153 76062 424978 76064
rect 408542 75986 408602 76062
rect 418153 76059 418219 76062
rect 408358 75926 408602 75986
rect 437430 75986 437490 76198
rect 456701 76122 456767 76125
rect 447182 76120 456767 76122
rect 447182 76064 456706 76120
rect 456762 76064 456767 76120
rect 447182 76062 456767 76064
rect 447182 75986 447242 76062
rect 456701 76059 456767 76062
rect 456885 76122 456951 76125
rect 475929 76122 475995 76125
rect 456885 76120 466378 76122
rect 456885 76064 456890 76120
rect 456946 76064 466378 76120
rect 456885 76062 466378 76064
rect 456885 76059 456951 76062
rect 437430 75926 447242 75986
rect 466318 75986 466378 76062
rect 466502 76120 475995 76122
rect 466502 76064 475934 76120
rect 475990 76064 475995 76120
rect 466502 76062 475995 76064
rect 466502 75986 466562 76062
rect 475929 76059 475995 76062
rect 478137 76122 478203 76125
rect 495206 76122 495266 76334
rect 478137 76120 482938 76122
rect 478137 76064 478142 76120
rect 478198 76064 482938 76120
rect 478137 76062 482938 76064
rect 478137 76059 478203 76062
rect 466318 75926 466562 75986
rect 482878 75986 482938 76062
rect 485822 76062 495266 76122
rect 485822 75986 485882 76062
rect 482878 75926 485882 75986
rect 502198 75986 502258 76334
rect 531262 76332 531268 76396
rect 531332 76394 531338 76396
rect 540881 76394 540947 76397
rect 531332 76392 540947 76394
rect 531332 76336 540886 76392
rect 540942 76336 540947 76392
rect 531332 76334 540947 76336
rect 531332 76332 531338 76334
rect 540881 76331 540947 76334
rect 560201 76258 560267 76261
rect 583520 76258 584960 76348
rect 560201 76256 563162 76258
rect 560201 76200 560206 76256
rect 560262 76200 563162 76256
rect 560201 76198 563162 76200
rect 560201 76195 560267 76198
rect 514569 76122 514635 76125
rect 505142 76120 514635 76122
rect 505142 76064 514574 76120
rect 514630 76064 514635 76120
rect 505142 76062 514635 76064
rect 505142 75986 505202 76062
rect 514569 76059 514635 76062
rect 516869 76122 516935 76125
rect 526437 76122 526503 76125
rect 531262 76122 531268 76124
rect 516869 76120 521578 76122
rect 516869 76064 516874 76120
rect 516930 76064 521578 76120
rect 516869 76062 521578 76064
rect 516869 76059 516935 76062
rect 502198 75926 505202 75986
rect 521518 75986 521578 76062
rect 526437 76120 531268 76122
rect 526437 76064 526442 76120
rect 526498 76064 531268 76120
rect 526437 76062 531268 76064
rect 526437 76059 526503 76062
rect 531262 76060 531268 76062
rect 531332 76060 531338 76124
rect 550582 76122 550588 76124
rect 543782 76062 550588 76122
rect 524229 75986 524295 75989
rect 521518 75984 524295 75986
rect 521518 75928 524234 75984
rect 524290 75928 524295 75984
rect 521518 75926 524295 75928
rect 350398 75892 350642 75926
rect 524229 75923 524295 75926
rect 540881 75986 540947 75989
rect 543782 75986 543842 76062
rect 550582 76060 550588 76062
rect 550652 76060 550658 76124
rect 540881 75984 543842 75986
rect 540881 75928 540886 75984
rect 540942 75928 543842 75984
rect 540881 75926 543842 75928
rect 563102 75986 563162 76198
rect 583342 76198 584960 76258
rect 572621 76122 572687 76125
rect 583342 76122 583402 76198
rect 569910 76120 572687 76122
rect 569910 76064 572626 76120
rect 572682 76064 572687 76120
rect 569910 76062 572687 76064
rect 569910 75986 569970 76062
rect 572621 76059 572687 76062
rect 576902 76062 583402 76122
rect 583520 76108 584960 76198
rect 563102 75926 569970 75986
rect 572713 75986 572779 75989
rect 576902 75986 576962 76062
rect 572713 75984 576962 75986
rect 572713 75928 572718 75984
rect 572774 75928 576962 75984
rect 572713 75926 576962 75928
rect 540881 75923 540947 75926
rect 572713 75923 572779 75926
rect 290549 75848 304274 75850
rect 290549 75792 290554 75848
rect 290610 75792 304274 75848
rect 290549 75790 304274 75792
rect 290549 75787 290615 75790
rect 550582 75788 550588 75852
rect 550652 75850 550658 75852
rect 560201 75850 560267 75853
rect 550652 75848 560267 75850
rect 550652 75792 560206 75848
rect 560262 75792 560267 75848
rect 550652 75790 560267 75792
rect 550652 75788 550658 75790
rect 560201 75787 560267 75790
rect 353385 66330 353451 66333
rect 353385 66328 353586 66330
rect 353385 66272 353390 66328
rect 353446 66272 353586 66328
rect 353385 66270 353586 66272
rect 353385 66267 353451 66270
rect 353526 66058 353586 66270
rect 353661 66058 353727 66061
rect 353526 66056 353727 66058
rect 353526 66000 353666 66056
rect 353722 66000 353727 66056
rect 353526 65998 353727 66000
rect 353661 65995 353727 65998
rect 240041 64972 240107 64973
rect 239990 64970 239996 64972
rect 239950 64910 239996 64970
rect 240060 64968 240107 64972
rect 240102 64912 240107 64968
rect 239990 64908 239996 64910
rect 240060 64908 240107 64912
rect 240041 64907 240107 64908
rect -960 64562 480 64652
rect 3601 64562 3667 64565
rect 583520 64562 584960 64652
rect -960 64560 3667 64562
rect -960 64504 3606 64560
rect 3662 64504 3667 64560
rect -960 64502 3667 64504
rect -960 64412 480 64502
rect 3601 64499 3667 64502
rect 583342 64502 584960 64562
rect 253105 64290 253171 64293
rect 253105 64288 258090 64290
rect 253105 64232 253110 64288
rect 253166 64232 258090 64288
rect 253105 64230 258090 64232
rect 253105 64227 253171 64230
rect 258030 64154 258090 64230
rect 304257 64154 304323 64157
rect 258030 64094 263610 64154
rect 263550 63882 263610 64094
rect 299430 64152 304323 64154
rect 299430 64096 304262 64152
rect 304318 64096 304323 64152
rect 299430 64094 304323 64096
rect 267641 63882 267707 63885
rect 263550 63880 267707 63882
rect 263550 63824 267646 63880
rect 267702 63824 267707 63880
rect 263550 63822 267707 63824
rect 267641 63819 267707 63822
rect 275921 63882 275987 63885
rect 277301 63882 277367 63885
rect 299430 63882 299490 64094
rect 304257 64091 304323 64094
rect 502006 64018 502012 64020
rect 495206 63958 502012 64018
rect 275921 63880 277367 63882
rect 275921 63824 275926 63880
rect 275982 63824 277306 63880
rect 277362 63824 277367 63880
rect 275921 63822 277367 63824
rect 275921 63819 275987 63822
rect 277301 63819 277367 63822
rect 286918 63822 299490 63882
rect 346485 63882 346551 63885
rect 355501 63882 355567 63885
rect 346485 63880 355567 63882
rect 346485 63824 346490 63880
rect 346546 63824 355506 63880
rect 355562 63824 355567 63880
rect 346485 63822 355567 63824
rect 286918 63746 286978 63822
rect 346485 63819 346551 63822
rect 355501 63819 355567 63822
rect 405641 63882 405707 63885
rect 418061 63882 418127 63885
rect 405641 63880 408418 63882
rect 405641 63824 405646 63880
rect 405702 63824 408418 63880
rect 405641 63822 408418 63824
rect 405641 63819 405707 63822
rect 373942 63746 373948 63748
rect 277350 63686 286978 63746
rect 364382 63686 373948 63746
rect 277350 63613 277410 63686
rect 248321 63610 248387 63613
rect 248321 63608 248522 63610
rect 248321 63552 248326 63608
rect 248382 63552 248522 63608
rect 248321 63550 248522 63552
rect 248321 63547 248387 63550
rect 248462 63338 248522 63550
rect 277301 63608 277410 63613
rect 277301 63552 277306 63608
rect 277362 63552 277410 63608
rect 277301 63550 277410 63552
rect 304257 63610 304323 63613
rect 309174 63610 309180 63612
rect 304257 63608 309180 63610
rect 304257 63552 304262 63608
rect 304318 63552 309180 63608
rect 304257 63550 309180 63552
rect 277301 63547 277367 63550
rect 304257 63547 304323 63550
rect 309174 63548 309180 63550
rect 309244 63548 309250 63612
rect 337469 63610 337535 63613
rect 330342 63608 337535 63610
rect 330342 63552 337474 63608
rect 337530 63552 337535 63608
rect 330342 63550 337535 63552
rect 253105 63338 253171 63341
rect 248462 63336 253171 63338
rect 248462 63280 253110 63336
rect 253166 63280 253171 63336
rect 248462 63278 253171 63280
rect 253105 63275 253171 63278
rect 309174 63276 309180 63340
rect 309244 63338 309250 63340
rect 330342 63338 330402 63550
rect 337469 63547 337535 63550
rect 344921 63610 344987 63613
rect 346209 63610 346275 63613
rect 344921 63608 346275 63610
rect 344921 63552 344926 63608
rect 344982 63552 346214 63608
rect 346270 63552 346275 63608
rect 344921 63550 346275 63552
rect 344921 63547 344987 63550
rect 346209 63547 346275 63550
rect 360377 63610 360443 63613
rect 364382 63610 364442 63686
rect 373942 63684 373948 63686
rect 374012 63684 374018 63748
rect 383561 63746 383627 63749
rect 393313 63746 393379 63749
rect 383561 63744 393379 63746
rect 383561 63688 383566 63744
rect 383622 63688 393318 63744
rect 393374 63688 393379 63744
rect 383561 63686 393379 63688
rect 383561 63683 383627 63686
rect 393313 63683 393379 63686
rect 360377 63608 364442 63610
rect 360377 63552 360382 63608
rect 360438 63552 364442 63608
rect 360377 63550 364442 63552
rect 408358 63610 408418 63822
rect 415350 63880 418127 63882
rect 415350 63824 418066 63880
rect 418122 63824 418127 63880
rect 415350 63822 418127 63824
rect 415350 63746 415410 63822
rect 418061 63819 418127 63822
rect 424918 63822 427738 63882
rect 408542 63686 415410 63746
rect 418153 63746 418219 63749
rect 424918 63746 424978 63822
rect 418153 63744 424978 63746
rect 418153 63688 418158 63744
rect 418214 63688 424978 63744
rect 418153 63686 424978 63688
rect 408542 63610 408602 63686
rect 418153 63683 418219 63686
rect 408358 63550 408602 63610
rect 427678 63610 427738 63822
rect 427862 63822 437490 63882
rect 427862 63610 427922 63822
rect 427678 63550 427922 63610
rect 437430 63610 437490 63822
rect 456701 63746 456767 63749
rect 447182 63744 456767 63746
rect 447182 63688 456706 63744
rect 456762 63688 456767 63744
rect 447182 63686 456767 63688
rect 447182 63610 447242 63686
rect 456701 63683 456767 63686
rect 456885 63746 456951 63749
rect 495206 63746 495266 63958
rect 502006 63956 502012 63958
rect 502076 63956 502082 64020
rect 531262 63956 531268 64020
rect 531332 64018 531338 64020
rect 540881 64018 540947 64021
rect 531332 64016 540947 64018
rect 531332 63960 540886 64016
rect 540942 63960 540947 64016
rect 531332 63958 540947 63960
rect 531332 63956 531338 63958
rect 540881 63955 540947 63958
rect 560201 63882 560267 63885
rect 560201 63880 563162 63882
rect 560201 63824 560206 63880
rect 560262 63824 563162 63880
rect 560201 63822 563162 63824
rect 560201 63819 560267 63822
rect 514569 63746 514635 63749
rect 456885 63744 466378 63746
rect 456885 63688 456890 63744
rect 456946 63688 466378 63744
rect 456885 63686 466378 63688
rect 456885 63683 456951 63686
rect 437430 63550 447242 63610
rect 466318 63610 466378 63686
rect 466502 63686 482938 63746
rect 466502 63610 466562 63686
rect 466318 63550 466562 63610
rect 482878 63610 482938 63686
rect 485822 63686 495266 63746
rect 505142 63744 514635 63746
rect 505142 63688 514574 63744
rect 514630 63688 514635 63744
rect 505142 63686 514635 63688
rect 485822 63610 485882 63686
rect 482878 63550 485882 63610
rect 360377 63547 360443 63550
rect 502190 63548 502196 63612
rect 502260 63610 502266 63612
rect 505142 63610 505202 63686
rect 514569 63683 514635 63686
rect 526437 63746 526503 63749
rect 531262 63746 531268 63748
rect 526437 63744 531268 63746
rect 526437 63688 526442 63744
rect 526498 63688 531268 63744
rect 526437 63686 531268 63688
rect 526437 63683 526503 63686
rect 531262 63684 531268 63686
rect 531332 63684 531338 63748
rect 550582 63746 550588 63748
rect 543782 63686 550588 63746
rect 521653 63610 521719 63613
rect 502260 63550 505202 63610
rect 521518 63608 521719 63610
rect 521518 63552 521658 63608
rect 521714 63552 521719 63608
rect 521518 63550 521719 63552
rect 502260 63548 502266 63550
rect 373942 63412 373948 63476
rect 374012 63474 374018 63476
rect 383561 63474 383627 63477
rect 374012 63472 383627 63474
rect 374012 63416 383566 63472
rect 383622 63416 383627 63472
rect 374012 63414 383627 63416
rect 374012 63412 374018 63414
rect 383561 63411 383627 63414
rect 309244 63278 330402 63338
rect 514569 63338 514635 63341
rect 521518 63338 521578 63550
rect 521653 63547 521719 63550
rect 540881 63610 540947 63613
rect 543782 63610 543842 63686
rect 550582 63684 550588 63686
rect 550652 63684 550658 63748
rect 540881 63608 543842 63610
rect 540881 63552 540886 63608
rect 540942 63552 543842 63608
rect 540881 63550 543842 63552
rect 563102 63610 563162 63822
rect 572621 63746 572687 63749
rect 583342 63746 583402 64502
rect 583520 64412 584960 64502
rect 569910 63744 572687 63746
rect 569910 63688 572626 63744
rect 572682 63688 572687 63744
rect 569910 63686 572687 63688
rect 569910 63610 569970 63686
rect 572621 63683 572687 63686
rect 576902 63686 583402 63746
rect 563102 63550 569970 63610
rect 572713 63610 572779 63613
rect 576902 63610 576962 63686
rect 572713 63608 576962 63610
rect 572713 63552 572718 63608
rect 572774 63552 576962 63608
rect 572713 63550 576962 63552
rect 540881 63547 540947 63550
rect 572713 63547 572779 63550
rect 550582 63412 550588 63476
rect 550652 63474 550658 63476
rect 560201 63474 560267 63477
rect 550652 63472 560267 63474
rect 550652 63416 560206 63472
rect 560262 63416 560267 63472
rect 550652 63414 560267 63416
rect 550652 63412 550658 63414
rect 560201 63411 560267 63414
rect 514569 63336 521578 63338
rect 514569 63280 514574 63336
rect 514630 63280 521578 63336
rect 514569 63278 521578 63280
rect 309244 63276 309250 63278
rect 514569 63275 514635 63278
rect 367369 55450 367435 55453
rect 367142 55448 367435 55450
rect 367142 55392 367374 55448
rect 367430 55392 367435 55448
rect 367142 55390 367435 55392
rect 367142 55314 367202 55390
rect 367369 55387 367435 55390
rect 367277 55314 367343 55317
rect 367142 55312 367343 55314
rect 367142 55256 367282 55312
rect 367338 55256 367343 55312
rect 367142 55254 367343 55256
rect 367277 55251 367343 55254
rect 255497 55178 255563 55181
rect 255773 55178 255839 55181
rect 255497 55176 255839 55178
rect 255497 55120 255502 55176
rect 255558 55120 255778 55176
rect 255834 55120 255839 55176
rect 255497 55118 255839 55120
rect 255497 55115 255563 55118
rect 255773 55115 255839 55118
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3509 50146 3575 50149
rect -960 50144 3575 50146
rect -960 50088 3514 50144
rect 3570 50088 3575 50144
rect -960 50086 3575 50088
rect -960 49996 480 50086
rect 3509 50083 3575 50086
rect 310881 47018 310947 47021
rect 310654 47016 310947 47018
rect 310654 46960 310886 47016
rect 310942 46960 310947 47016
rect 310654 46958 310947 46960
rect 310654 46746 310714 46958
rect 310881 46955 310947 46958
rect 310789 46746 310855 46749
rect 310654 46744 310855 46746
rect 310654 46688 310794 46744
rect 310850 46688 310855 46744
rect 310654 46686 310855 46688
rect 310789 46683 310855 46686
rect 367369 45658 367435 45661
rect 367326 45656 367435 45658
rect 367326 45600 367374 45656
rect 367430 45600 367435 45656
rect 367326 45595 367435 45600
rect 367326 45522 367386 45595
rect 367461 45522 367527 45525
rect 367326 45520 367527 45522
rect 367326 45464 367466 45520
rect 367522 45464 367527 45520
rect 367326 45462 367527 45464
rect 367461 45459 367527 45462
rect 234102 43828 234108 43892
rect 234172 43890 234178 43892
rect 240041 43890 240107 43893
rect 234172 43888 240107 43890
rect 234172 43832 240046 43888
rect 240102 43832 240107 43888
rect 234172 43830 240107 43832
rect 234172 43828 234178 43830
rect 240041 43827 240107 43830
rect 583520 41034 584960 41124
rect 583342 40974 584960 41034
rect 258022 40490 258028 40492
rect 254534 40430 258028 40490
rect 240041 40218 240107 40221
rect 254534 40218 254594 40430
rect 258022 40428 258028 40430
rect 258092 40428 258098 40492
rect 349797 40490 349863 40493
rect 412449 40490 412515 40493
rect 413921 40490 413987 40493
rect 349797 40488 359658 40490
rect 349797 40432 349802 40488
rect 349858 40432 359658 40488
rect 349797 40430 359658 40432
rect 349797 40427 349863 40430
rect 267733 40354 267799 40357
rect 240041 40216 254594 40218
rect 240041 40160 240046 40216
rect 240102 40160 254594 40216
rect 240041 40158 254594 40160
rect 267598 40352 267799 40354
rect 267598 40296 267738 40352
rect 267794 40296 267799 40352
rect 267598 40294 267799 40296
rect 240041 40155 240107 40158
rect 258022 40020 258028 40084
rect 258092 40082 258098 40084
rect 267598 40082 267658 40294
rect 267733 40291 267799 40294
rect 277301 40354 277367 40357
rect 278681 40354 278747 40357
rect 277301 40352 278747 40354
rect 277301 40296 277306 40352
rect 277362 40296 278686 40352
rect 278742 40296 278747 40352
rect 277301 40294 278747 40296
rect 277301 40291 277367 40294
rect 278681 40291 278747 40294
rect 293174 40294 302986 40354
rect 258092 40022 267658 40082
rect 278681 40082 278747 40085
rect 293174 40082 293234 40294
rect 278681 40080 293234 40082
rect 278681 40024 278686 40080
rect 278742 40024 293234 40080
rect 278681 40022 293234 40024
rect 302926 40082 302986 40294
rect 317321 40218 317387 40221
rect 326797 40218 326863 40221
rect 317321 40216 326863 40218
rect 317321 40160 317326 40216
rect 317382 40160 326802 40216
rect 326858 40160 326863 40216
rect 317321 40158 326863 40160
rect 317321 40155 317387 40158
rect 326797 40155 326863 40158
rect 341057 40218 341123 40221
rect 349797 40218 349863 40221
rect 341057 40216 349863 40218
rect 341057 40160 341062 40216
rect 341118 40160 349802 40216
rect 349858 40160 349863 40216
rect 341057 40158 349863 40160
rect 341057 40155 341123 40158
rect 349797 40155 349863 40158
rect 311801 40082 311867 40085
rect 302926 40080 311867 40082
rect 302926 40024 311806 40080
rect 311862 40024 311867 40080
rect 302926 40022 311867 40024
rect 258092 40020 258098 40022
rect 278681 40019 278747 40022
rect 311801 40019 311867 40022
rect 326981 40082 327047 40085
rect 335302 40082 335308 40084
rect 326981 40080 335308 40082
rect 326981 40024 326986 40080
rect 327042 40024 335308 40080
rect 326981 40022 335308 40024
rect 326981 40019 327047 40022
rect 335302 40020 335308 40022
rect 335372 40020 335378 40084
rect 359598 40082 359658 40430
rect 412449 40488 413987 40490
rect 412449 40432 412454 40488
rect 412510 40432 413926 40488
rect 413982 40432 413987 40488
rect 412449 40430 413987 40432
rect 412449 40427 412515 40430
rect 413921 40427 413987 40430
rect 492630 40430 502258 40490
rect 383694 40292 383700 40356
rect 383764 40354 383770 40356
rect 402973 40354 403039 40357
rect 383764 40352 403039 40354
rect 383764 40296 402978 40352
rect 403034 40296 403039 40352
rect 383764 40294 403039 40296
rect 383764 40292 383770 40294
rect 402973 40291 403039 40294
rect 424918 40294 427738 40354
rect 383561 40218 383627 40221
rect 413921 40218 413987 40221
rect 424918 40218 424978 40294
rect 383561 40216 383762 40218
rect 383561 40160 383566 40216
rect 383622 40160 383762 40216
rect 383561 40158 383762 40160
rect 383561 40155 383627 40158
rect 383561 40082 383627 40085
rect 383702 40084 383762 40158
rect 413921 40216 424978 40218
rect 413921 40160 413926 40216
rect 413982 40160 424978 40216
rect 413921 40158 424978 40160
rect 413921 40155 413987 40158
rect 359598 40022 364442 40082
rect 364382 39946 364442 40022
rect 373950 40080 383627 40082
rect 373950 40024 383566 40080
rect 383622 40024 383627 40080
rect 373950 40022 383627 40024
rect 373950 39946 374010 40022
rect 383561 40019 383627 40022
rect 383694 40020 383700 40084
rect 383764 40020 383770 40084
rect 427678 40082 427738 40294
rect 427862 40294 437490 40354
rect 427862 40082 427922 40294
rect 427678 40022 427922 40082
rect 437430 40082 437490 40294
rect 456701 40218 456767 40221
rect 447182 40216 456767 40218
rect 447182 40160 456706 40216
rect 456762 40160 456767 40216
rect 447182 40158 456767 40160
rect 447182 40082 447242 40158
rect 456701 40155 456767 40158
rect 456885 40218 456951 40221
rect 492630 40218 492690 40430
rect 502198 40356 502258 40430
rect 531262 40428 531268 40492
rect 531332 40490 531338 40492
rect 540881 40490 540947 40493
rect 531332 40488 540947 40490
rect 531332 40432 540886 40488
rect 540942 40432 540947 40488
rect 531332 40430 540947 40432
rect 531332 40428 531338 40430
rect 540881 40427 540947 40430
rect 502190 40292 502196 40356
rect 502260 40292 502266 40356
rect 560201 40354 560267 40357
rect 560201 40352 563162 40354
rect 560201 40296 560206 40352
rect 560262 40296 563162 40352
rect 560201 40294 563162 40296
rect 560201 40291 560267 40294
rect 514569 40218 514635 40221
rect 456885 40216 466378 40218
rect 456885 40160 456890 40216
rect 456946 40160 466378 40216
rect 456885 40158 466378 40160
rect 456885 40155 456951 40158
rect 437430 40022 447242 40082
rect 466318 40082 466378 40158
rect 466502 40158 482938 40218
rect 466502 40082 466562 40158
rect 466318 40022 466562 40082
rect 482878 40082 482938 40158
rect 485822 40158 492690 40218
rect 505142 40216 514635 40218
rect 505142 40160 514574 40216
rect 514630 40160 514635 40216
rect 505142 40158 514635 40160
rect 485822 40082 485882 40158
rect 482878 40022 485882 40082
rect 502190 40020 502196 40084
rect 502260 40082 502266 40084
rect 505142 40082 505202 40158
rect 514569 40155 514635 40158
rect 526437 40218 526503 40221
rect 531262 40218 531268 40220
rect 526437 40216 531268 40218
rect 526437 40160 526442 40216
rect 526498 40160 531268 40216
rect 526437 40158 531268 40160
rect 526437 40155 526503 40158
rect 531262 40156 531268 40158
rect 531332 40156 531338 40220
rect 550582 40218 550588 40220
rect 543782 40158 550588 40218
rect 521653 40082 521719 40085
rect 502260 40022 505202 40082
rect 521518 40080 521719 40082
rect 521518 40024 521658 40080
rect 521714 40024 521719 40080
rect 521518 40022 521719 40024
rect 502260 40020 502266 40022
rect 364382 39886 374010 39946
rect 335302 39748 335308 39812
rect 335372 39810 335378 39812
rect 341057 39810 341123 39813
rect 335372 39808 341123 39810
rect 335372 39752 341062 39808
rect 341118 39752 341123 39808
rect 335372 39750 341123 39752
rect 335372 39748 335378 39750
rect 341057 39747 341123 39750
rect 514569 39810 514635 39813
rect 521518 39810 521578 40022
rect 521653 40019 521719 40022
rect 540881 40082 540947 40085
rect 543782 40082 543842 40158
rect 550582 40156 550588 40158
rect 550652 40156 550658 40220
rect 540881 40080 543842 40082
rect 540881 40024 540886 40080
rect 540942 40024 543842 40080
rect 540881 40022 543842 40024
rect 563102 40082 563162 40294
rect 572621 40218 572687 40221
rect 583342 40218 583402 40974
rect 583520 40884 584960 40974
rect 569910 40216 572687 40218
rect 569910 40160 572626 40216
rect 572682 40160 572687 40216
rect 569910 40158 572687 40160
rect 569910 40082 569970 40158
rect 572621 40155 572687 40158
rect 576902 40158 583402 40218
rect 563102 40022 569970 40082
rect 572713 40082 572779 40085
rect 576902 40082 576962 40158
rect 572713 40080 576962 40082
rect 572713 40024 572718 40080
rect 572774 40024 576962 40080
rect 572713 40022 576962 40024
rect 540881 40019 540947 40022
rect 572713 40019 572779 40022
rect 550582 39884 550588 39948
rect 550652 39946 550658 39948
rect 560201 39946 560267 39949
rect 550652 39944 560267 39946
rect 550652 39888 560206 39944
rect 560262 39888 560267 39944
rect 550652 39886 560267 39888
rect 550652 39884 550658 39886
rect 560201 39883 560267 39886
rect 514569 39808 521578 39810
rect 514569 39752 514574 39808
rect 514630 39752 521578 39808
rect 514569 39750 521578 39752
rect 514569 39747 514635 39750
rect -960 35866 480 35956
rect 3509 35866 3575 35869
rect -960 35864 3575 35866
rect -960 35808 3514 35864
rect 3570 35808 3575 35864
rect -960 35806 3575 35808
rect -960 35716 480 35806
rect 3509 35803 3575 35806
rect 338062 29548 338068 29612
rect 338132 29610 338138 29612
rect 338132 29550 345122 29610
rect 338132 29548 338138 29550
rect 317321 29474 317387 29477
rect 318701 29474 318767 29477
rect 246254 29414 256066 29474
rect 237230 29276 237236 29340
rect 237300 29338 237306 29340
rect 246254 29338 246314 29414
rect 237300 29278 246314 29338
rect 237300 29276 237306 29278
rect 256006 29202 256066 29414
rect 317321 29472 318767 29474
rect 317321 29416 317326 29472
rect 317382 29416 318706 29472
rect 318762 29416 318767 29472
rect 317321 29414 318767 29416
rect 345062 29474 345122 29550
rect 373942 29548 373948 29612
rect 374012 29610 374018 29612
rect 383561 29610 383627 29613
rect 374012 29608 383627 29610
rect 374012 29552 383566 29608
rect 383622 29552 383627 29608
rect 374012 29550 383627 29552
rect 374012 29548 374018 29550
rect 383561 29547 383627 29550
rect 453982 29548 453988 29612
rect 454052 29610 454058 29612
rect 454052 29550 463618 29610
rect 454052 29548 454058 29550
rect 350993 29474 351059 29477
rect 463558 29476 463618 29550
rect 550582 29548 550588 29612
rect 550652 29610 550658 29612
rect 560201 29610 560267 29613
rect 550652 29608 560267 29610
rect 550652 29552 560206 29608
rect 560262 29552 560267 29608
rect 550652 29550 560267 29552
rect 550652 29548 550658 29550
rect 560201 29547 560267 29550
rect 345062 29472 351059 29474
rect 345062 29416 350998 29472
rect 351054 29416 351059 29472
rect 345062 29414 351059 29416
rect 317321 29411 317387 29414
rect 318701 29411 318767 29414
rect 350993 29411 351059 29414
rect 413326 29414 417986 29474
rect 293217 29338 293283 29341
rect 318701 29340 318767 29341
rect 373901 29340 373967 29341
rect 293217 29336 299490 29338
rect 293217 29280 293222 29336
rect 293278 29280 299490 29336
rect 293217 29278 299490 29280
rect 293217 29275 293283 29278
rect 274081 29202 274147 29205
rect 256006 29200 274147 29202
rect 256006 29144 274086 29200
rect 274142 29144 274147 29200
rect 256006 29142 274147 29144
rect 274081 29139 274147 29142
rect 274265 29202 274331 29205
rect 278773 29202 278839 29205
rect 274265 29200 278839 29202
rect 274265 29144 274270 29200
rect 274326 29144 278778 29200
rect 278834 29144 278839 29200
rect 274265 29142 278839 29144
rect 274265 29139 274331 29142
rect 278773 29139 278839 29142
rect 283097 29202 283163 29205
rect 288382 29202 288388 29204
rect 283097 29200 288388 29202
rect 283097 29144 283102 29200
rect 283158 29144 288388 29200
rect 283097 29142 288388 29144
rect 283097 29139 283163 29142
rect 288382 29140 288388 29142
rect 288452 29140 288458 29204
rect 299430 29202 299490 29278
rect 318701 29336 318748 29340
rect 318812 29338 318818 29340
rect 338062 29338 338068 29340
rect 318701 29280 318706 29336
rect 318701 29276 318748 29280
rect 318812 29278 318894 29338
rect 331814 29278 338068 29338
rect 318812 29276 318818 29278
rect 318701 29275 318767 29276
rect 307702 29202 307708 29204
rect 299430 29142 307708 29202
rect 307702 29140 307708 29142
rect 307772 29140 307778 29204
rect 331814 29202 331874 29278
rect 338062 29276 338068 29278
rect 338132 29276 338138 29340
rect 373901 29336 373948 29340
rect 374012 29338 374018 29340
rect 373901 29280 373906 29336
rect 373901 29276 373948 29280
rect 374012 29278 374094 29338
rect 374012 29276 374018 29278
rect 373901 29275 373967 29276
rect 323718 29142 331874 29202
rect 350993 29202 351059 29205
rect 383561 29202 383627 29205
rect 395889 29202 395955 29205
rect 350993 29200 355978 29202
rect 350993 29144 350998 29200
rect 351054 29144 355978 29200
rect 350993 29142 355978 29144
rect 318742 29004 318748 29068
rect 318812 29066 318818 29068
rect 323718 29066 323778 29142
rect 350993 29139 351059 29142
rect 318812 29006 323778 29066
rect 318812 29004 318818 29006
rect 288382 28868 288388 28932
rect 288452 28930 288458 28932
rect 293217 28930 293283 28933
rect 288452 28928 293283 28930
rect 288452 28872 293222 28928
rect 293278 28872 293283 28928
rect 288452 28870 293283 28872
rect 288452 28868 288458 28870
rect 293217 28867 293283 28870
rect 307702 28868 307708 28932
rect 307772 28930 307778 28932
rect 317321 28930 317387 28933
rect 307772 28928 317387 28930
rect 307772 28872 317326 28928
rect 317382 28872 317387 28928
rect 307772 28870 317387 28872
rect 355918 28930 355978 29142
rect 383561 29200 395955 29202
rect 383561 29144 383566 29200
rect 383622 29144 395894 29200
rect 395950 29144 395955 29200
rect 383561 29142 395955 29144
rect 383561 29139 383627 29142
rect 395889 29139 395955 29142
rect 396073 29202 396139 29205
rect 413326 29202 413386 29414
rect 396073 29200 413386 29202
rect 396073 29144 396078 29200
rect 396134 29144 413386 29200
rect 396073 29142 413386 29144
rect 417926 29202 417986 29414
rect 463550 29412 463556 29476
rect 463620 29412 463626 29476
rect 502190 29474 502196 29476
rect 495206 29414 502196 29474
rect 473261 29338 473327 29341
rect 427678 29278 437490 29338
rect 417926 29142 418538 29202
rect 396073 29139 396139 29142
rect 418478 29066 418538 29142
rect 427678 29066 427738 29278
rect 418478 29006 427738 29066
rect 437430 29066 437490 29278
rect 473261 29336 476130 29338
rect 473261 29280 473266 29336
rect 473322 29280 476130 29336
rect 473261 29278 476130 29280
rect 473261 29275 473327 29278
rect 453982 29202 453988 29204
rect 447182 29142 453988 29202
rect 447182 29066 447242 29142
rect 453982 29140 453988 29142
rect 454052 29140 454058 29204
rect 437430 29006 447242 29066
rect 463550 29004 463556 29068
rect 463620 29066 463626 29068
rect 466269 29066 466335 29069
rect 463620 29064 466335 29066
rect 463620 29008 466274 29064
rect 466330 29008 466335 29064
rect 463620 29006 466335 29008
rect 476070 29066 476130 29278
rect 495206 29202 495266 29414
rect 502190 29412 502196 29414
rect 502260 29412 502266 29476
rect 521510 29474 521516 29476
rect 514526 29414 521516 29474
rect 514526 29202 514586 29414
rect 521510 29412 521516 29414
rect 521580 29412 521586 29476
rect 531262 29412 531268 29476
rect 531332 29474 531338 29476
rect 540789 29474 540855 29477
rect 531332 29472 540855 29474
rect 531332 29416 540794 29472
rect 540850 29416 540855 29472
rect 531332 29414 540855 29416
rect 531332 29412 531338 29414
rect 540789 29411 540855 29414
rect 560201 29338 560267 29341
rect 583520 29338 584960 29428
rect 560201 29336 563162 29338
rect 560201 29280 560206 29336
rect 560262 29280 563162 29336
rect 560201 29278 563162 29280
rect 560201 29275 560267 29278
rect 485822 29142 495266 29202
rect 505142 29142 514586 29202
rect 525885 29202 525951 29205
rect 531262 29202 531268 29204
rect 525885 29200 531268 29202
rect 525885 29144 525890 29200
rect 525946 29144 531268 29200
rect 525885 29142 531268 29144
rect 485822 29066 485882 29142
rect 476070 29006 485882 29066
rect 463620 29004 463626 29006
rect 466269 29003 466335 29006
rect 502190 29004 502196 29068
rect 502260 29066 502266 29068
rect 505142 29066 505202 29142
rect 525885 29139 525951 29142
rect 531262 29140 531268 29142
rect 531332 29140 531338 29204
rect 550582 29202 550588 29204
rect 543782 29142 550588 29202
rect 502260 29006 505202 29066
rect 502260 29004 502266 29006
rect 521510 29004 521516 29068
rect 521580 29066 521586 29068
rect 521653 29066 521719 29069
rect 521580 29064 521719 29066
rect 521580 29008 521658 29064
rect 521714 29008 521719 29064
rect 521580 29006 521719 29008
rect 521580 29004 521586 29006
rect 521653 29003 521719 29006
rect 540881 29066 540947 29069
rect 543782 29066 543842 29142
rect 550582 29140 550588 29142
rect 550652 29140 550658 29204
rect 540881 29064 543842 29066
rect 540881 29008 540886 29064
rect 540942 29008 543842 29064
rect 540881 29006 543842 29008
rect 563102 29066 563162 29278
rect 583342 29278 584960 29338
rect 572621 29202 572687 29205
rect 569910 29200 572687 29202
rect 569910 29144 572626 29200
rect 572682 29144 572687 29200
rect 569910 29142 572687 29144
rect 569910 29066 569970 29142
rect 572621 29139 572687 29142
rect 576761 29202 576827 29205
rect 583342 29202 583402 29278
rect 576761 29200 583402 29202
rect 576761 29144 576766 29200
rect 576822 29144 583402 29200
rect 583520 29188 584960 29278
rect 576761 29142 583402 29144
rect 576761 29139 576827 29142
rect 563102 29006 569970 29066
rect 540881 29003 540947 29006
rect 364198 28930 364442 28964
rect 373901 28930 373967 28933
rect 355918 28928 373967 28930
rect 355918 28904 373906 28928
rect 355918 28870 364258 28904
rect 364382 28872 373906 28904
rect 373962 28872 373967 28928
rect 364382 28870 373967 28872
rect 307772 28868 307778 28870
rect 317321 28867 317387 28870
rect 373901 28867 373967 28870
rect 408677 27570 408743 27573
rect 408542 27568 408743 27570
rect 408542 27512 408682 27568
rect 408738 27512 408743 27568
rect 408542 27510 408743 27512
rect 408542 27434 408602 27510
rect 408677 27507 408743 27510
rect 408769 27434 408835 27437
rect 408542 27432 408835 27434
rect 408542 27376 408774 27432
rect 408830 27376 408835 27432
rect 408542 27374 408835 27376
rect 408769 27371 408835 27374
rect 336549 24850 336615 24853
rect 336733 24850 336799 24853
rect 336549 24848 336799 24850
rect 336549 24792 336554 24848
rect 336610 24792 336738 24848
rect 336794 24792 336799 24848
rect 336549 24790 336799 24792
rect 336549 24787 336615 24790
rect 336733 24787 336799 24790
rect 356329 24850 356395 24853
rect 356513 24850 356579 24853
rect 356329 24848 356579 24850
rect 356329 24792 356334 24848
rect 356390 24792 356518 24848
rect 356574 24792 356579 24848
rect 356329 24790 356579 24792
rect 356329 24787 356395 24790
rect 356513 24787 356579 24790
rect 527214 21994 527220 21996
rect 614 21934 527220 21994
rect -960 21450 480 21540
rect 614 21450 674 21934
rect 527214 21932 527220 21934
rect 527284 21932 527290 21996
rect -960 21390 674 21450
rect -960 21300 480 21390
rect 309409 18186 309475 18189
rect 309182 18184 309475 18186
rect 309182 18128 309414 18184
rect 309470 18128 309475 18184
rect 309182 18126 309475 18128
rect 309182 18050 309242 18126
rect 309409 18123 309475 18126
rect 309317 18050 309383 18053
rect 309182 18048 309383 18050
rect 309182 17992 309322 18048
rect 309378 17992 309383 18048
rect 309182 17990 309383 17992
rect 309317 17987 309383 17990
rect 583520 17642 584960 17732
rect 583342 17582 584960 17642
rect 259494 17308 259500 17372
rect 259564 17370 259570 17372
rect 268878 17370 268884 17372
rect 259564 17310 268884 17370
rect 259564 17308 259570 17310
rect 268878 17308 268884 17310
rect 268948 17308 268954 17372
rect 355961 17234 356027 17237
rect 357382 17234 357388 17236
rect 355961 17232 357388 17234
rect 355961 17176 355966 17232
rect 356022 17176 357388 17232
rect 355961 17174 357388 17176
rect 355961 17171 356027 17174
rect 357382 17172 357388 17174
rect 357452 17172 357458 17236
rect 251081 17098 251147 17101
rect 259494 17098 259500 17100
rect 251081 17096 259500 17098
rect 251081 17040 251086 17096
rect 251142 17040 259500 17096
rect 251081 17038 259500 17040
rect 251081 17035 251147 17038
rect 259494 17036 259500 17038
rect 259564 17036 259570 17100
rect 367134 17036 367140 17100
rect 367204 17098 367210 17100
rect 367204 17038 367386 17098
rect 367204 17036 367210 17038
rect 306414 16962 306420 16964
rect 280110 16902 282930 16962
rect 231710 16764 231716 16828
rect 231780 16826 231786 16828
rect 240133 16826 240199 16829
rect 231780 16824 240199 16826
rect 231780 16768 240138 16824
rect 240194 16768 240199 16824
rect 231780 16766 240199 16768
rect 231780 16764 231786 16766
rect 240133 16763 240199 16766
rect 240225 16690 240291 16693
rect 251081 16690 251147 16693
rect 280110 16690 280170 16902
rect 240225 16688 251147 16690
rect 240225 16632 240230 16688
rect 240286 16632 251086 16688
rect 251142 16632 251147 16688
rect 240225 16630 251147 16632
rect 240225 16627 240291 16630
rect 251081 16627 251147 16630
rect 273302 16630 280170 16690
rect 282870 16690 282930 16902
rect 303846 16902 306420 16962
rect 282870 16630 289922 16690
rect 269062 16492 269068 16556
rect 269132 16554 269138 16556
rect 273302 16554 273362 16630
rect 269132 16494 273362 16554
rect 289862 16554 289922 16630
rect 303846 16554 303906 16902
rect 306414 16900 306420 16902
rect 306484 16900 306490 16964
rect 357382 16900 357388 16964
rect 357452 16962 357458 16964
rect 367326 16962 367386 17038
rect 425094 17036 425100 17100
rect 425164 17036 425170 17100
rect 502006 17098 502012 17100
rect 495206 17038 502012 17098
rect 405733 16962 405799 16965
rect 418061 16962 418127 16965
rect 357452 16902 357634 16962
rect 367326 16902 381554 16962
rect 357452 16900 357458 16902
rect 319621 16826 319687 16829
rect 347681 16826 347747 16829
rect 319621 16824 329114 16826
rect 319621 16768 319626 16824
rect 319682 16768 329114 16824
rect 319621 16766 329114 16768
rect 319621 16763 319687 16766
rect 306598 16628 306604 16692
rect 306668 16690 306674 16692
rect 318701 16690 318767 16693
rect 306668 16688 318767 16690
rect 306668 16632 318706 16688
rect 318762 16632 318767 16688
rect 306668 16630 318767 16632
rect 329054 16690 329114 16766
rect 346350 16824 347747 16826
rect 346350 16768 347686 16824
rect 347742 16768 347747 16824
rect 346350 16766 347747 16768
rect 357574 16826 357634 16902
rect 367134 16826 367140 16828
rect 357574 16766 367140 16826
rect 334065 16690 334131 16693
rect 329054 16688 334131 16690
rect 329054 16632 334070 16688
rect 334126 16632 334131 16688
rect 329054 16630 334131 16632
rect 306668 16628 306674 16630
rect 318701 16627 318767 16630
rect 334065 16627 334131 16630
rect 338113 16690 338179 16693
rect 346350 16690 346410 16766
rect 347681 16763 347747 16766
rect 367134 16764 367140 16766
rect 367204 16764 367210 16828
rect 381494 16826 381554 16902
rect 391062 16902 400874 16962
rect 391062 16826 391122 16902
rect 381494 16766 391122 16826
rect 400814 16826 400874 16902
rect 405733 16960 418127 16962
rect 405733 16904 405738 16960
rect 405794 16904 418066 16960
rect 418122 16904 418127 16960
rect 405733 16902 418127 16904
rect 405733 16899 405799 16902
rect 418061 16899 418127 16902
rect 418245 16962 418311 16965
rect 425102 16962 425162 17036
rect 418245 16960 425162 16962
rect 418245 16904 418250 16960
rect 418306 16904 425162 16960
rect 418245 16902 425162 16904
rect 427678 16902 437490 16962
rect 418245 16899 418311 16902
rect 405733 16826 405799 16829
rect 400814 16824 405799 16826
rect 400814 16768 405738 16824
rect 405794 16768 405799 16824
rect 400814 16766 405799 16768
rect 405733 16763 405799 16766
rect 425094 16764 425100 16828
rect 425164 16826 425170 16828
rect 427678 16826 427738 16902
rect 425164 16766 427738 16826
rect 425164 16764 425170 16766
rect 338113 16688 346410 16690
rect 338113 16632 338118 16688
rect 338174 16632 346410 16688
rect 338113 16630 346410 16632
rect 437430 16690 437490 16902
rect 456701 16826 456767 16829
rect 447182 16824 456767 16826
rect 447182 16768 456706 16824
rect 456762 16768 456767 16824
rect 447182 16766 456767 16768
rect 447182 16690 447242 16766
rect 456701 16763 456767 16766
rect 456885 16826 456951 16829
rect 495206 16826 495266 17038
rect 502006 17036 502012 17038
rect 502076 17036 502082 17100
rect 531262 17036 531268 17100
rect 531332 17098 531338 17100
rect 540881 17098 540947 17101
rect 531332 17096 540947 17098
rect 531332 17040 540886 17096
rect 540942 17040 540947 17096
rect 531332 17038 540947 17040
rect 531332 17036 531338 17038
rect 540881 17035 540947 17038
rect 560201 16962 560267 16965
rect 560201 16960 563162 16962
rect 560201 16904 560206 16960
rect 560262 16904 563162 16960
rect 560201 16902 563162 16904
rect 560201 16899 560267 16902
rect 514569 16826 514635 16829
rect 456885 16824 466378 16826
rect 456885 16768 456890 16824
rect 456946 16768 466378 16824
rect 456885 16766 466378 16768
rect 456885 16763 456951 16766
rect 437430 16630 447242 16690
rect 466318 16690 466378 16766
rect 466502 16766 482938 16826
rect 466502 16690 466562 16766
rect 466318 16630 466562 16690
rect 482878 16690 482938 16766
rect 485822 16766 495266 16826
rect 505142 16824 514635 16826
rect 505142 16768 514574 16824
rect 514630 16768 514635 16824
rect 505142 16766 514635 16768
rect 485822 16690 485882 16766
rect 482878 16630 485882 16690
rect 338113 16627 338179 16630
rect 502190 16628 502196 16692
rect 502260 16690 502266 16692
rect 505142 16690 505202 16766
rect 514569 16763 514635 16766
rect 516041 16826 516107 16829
rect 526437 16826 526503 16829
rect 531262 16826 531268 16828
rect 516041 16824 521578 16826
rect 516041 16768 516046 16824
rect 516102 16768 521578 16824
rect 516041 16766 521578 16768
rect 516041 16763 516107 16766
rect 502260 16630 505202 16690
rect 521518 16690 521578 16766
rect 526437 16824 531268 16826
rect 526437 16768 526442 16824
rect 526498 16768 531268 16824
rect 526437 16766 531268 16768
rect 526437 16763 526503 16766
rect 531262 16764 531268 16766
rect 531332 16764 531338 16828
rect 550582 16826 550588 16828
rect 543782 16766 550588 16826
rect 524229 16690 524295 16693
rect 521518 16688 524295 16690
rect 521518 16632 524234 16688
rect 524290 16632 524295 16688
rect 521518 16630 524295 16632
rect 502260 16628 502266 16630
rect 524229 16627 524295 16630
rect 540881 16690 540947 16693
rect 543782 16690 543842 16766
rect 550582 16764 550588 16766
rect 550652 16764 550658 16828
rect 540881 16688 543842 16690
rect 540881 16632 540886 16688
rect 540942 16632 543842 16688
rect 540881 16630 543842 16632
rect 563102 16690 563162 16902
rect 572621 16826 572687 16829
rect 583342 16826 583402 17582
rect 583520 17492 584960 17582
rect 569910 16824 572687 16826
rect 569910 16768 572626 16824
rect 572682 16768 572687 16824
rect 569910 16766 572687 16768
rect 569910 16690 569970 16766
rect 572621 16763 572687 16766
rect 576902 16766 583402 16826
rect 563102 16630 569970 16690
rect 572713 16690 572779 16693
rect 576902 16690 576962 16766
rect 572713 16688 576962 16690
rect 572713 16632 572718 16688
rect 572774 16632 576962 16688
rect 572713 16630 576962 16632
rect 540881 16627 540947 16630
rect 572713 16627 572779 16630
rect 289862 16494 303906 16554
rect 269132 16492 269138 16494
rect 550582 16492 550588 16556
rect 550652 16554 550658 16556
rect 560201 16554 560267 16557
rect 550652 16552 560267 16554
rect 550652 16496 560206 16552
rect 560262 16496 560267 16552
rect 550652 16494 560267 16496
rect 550652 16492 550658 16494
rect 560201 16491 560267 16494
rect 60641 10298 60707 10301
rect 259729 10298 259795 10301
rect 60641 10296 259795 10298
rect 60641 10240 60646 10296
rect 60702 10240 259734 10296
rect 259790 10240 259795 10296
rect 60641 10238 259795 10240
rect 60641 10235 60707 10238
rect 259729 10235 259795 10238
rect 136081 8938 136147 8941
rect 299565 8938 299631 8941
rect 136081 8936 299631 8938
rect 136081 8880 136086 8936
rect 136142 8880 299570 8936
rect 299626 8880 299631 8936
rect 136081 8878 299631 8880
rect 136081 8875 136147 8878
rect 299565 8875 299631 8878
rect 134885 7578 134951 7581
rect 298277 7578 298343 7581
rect 134885 7576 298343 7578
rect 134885 7520 134890 7576
rect 134946 7520 298282 7576
rect 298338 7520 298343 7576
rect 134885 7518 298343 7520
rect 134885 7515 134951 7518
rect 298277 7515 298343 7518
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 48129 6218 48195 6221
rect 253933 6218 253999 6221
rect 48129 6216 253999 6218
rect 48129 6160 48134 6216
rect 48190 6160 253938 6216
rect 253994 6160 253999 6216
rect 48129 6158 253999 6160
rect 48129 6155 48195 6158
rect 253933 6155 253999 6158
rect 583520 5796 584960 6036
rect 219341 4858 219407 4861
rect 342253 4858 342319 4861
rect 219341 4856 342319 4858
rect 219341 4800 219346 4856
rect 219402 4800 342258 4856
rect 342314 4800 342319 4856
rect 219341 4798 342319 4800
rect 219341 4795 219407 4798
rect 342253 4795 342319 4798
rect 408309 3634 408375 3637
rect 408585 3634 408651 3637
rect 408309 3632 408651 3634
rect 408309 3576 408314 3632
rect 408370 3576 408590 3632
rect 408646 3576 408651 3632
rect 408309 3574 408651 3576
rect 408309 3571 408375 3574
rect 408585 3571 408651 3574
rect 6453 3362 6519 3365
rect 231853 3362 231919 3365
rect 6453 3360 231919 3362
rect 6453 3304 6458 3360
rect 6514 3304 231858 3360
rect 231914 3304 231919 3360
rect 6453 3302 231919 3304
rect 6453 3299 6519 3302
rect 231853 3299 231919 3302
rect 356145 3362 356211 3365
rect 410517 3362 410583 3365
rect 356145 3360 410583 3362
rect 356145 3304 356150 3360
rect 356206 3304 410522 3360
rect 410578 3304 410583 3360
rect 356145 3302 410583 3304
rect 356145 3299 356211 3302
rect 410517 3299 410583 3302
rect 525701 3362 525767 3365
rect 575013 3362 575079 3365
rect 525701 3360 575079 3362
rect 525701 3304 525706 3360
rect 525762 3304 575018 3360
rect 575074 3304 575079 3360
rect 525701 3302 575079 3304
rect 525701 3299 525767 3302
rect 575013 3299 575079 3302
<< via3 >>
rect 527404 642772 527468 642836
rect 258948 642636 259012 642700
rect 261892 642500 261956 642564
rect 261708 642364 261772 642428
rect 261524 642228 261588 642292
rect 258764 642092 258828 642156
rect 527956 641956 528020 642020
rect 258580 641820 258644 641884
rect 402836 639644 402900 639708
rect 384988 639372 385052 639436
rect 231716 639236 231780 639300
rect 234476 639236 234540 639300
rect 237236 639236 237300 639300
rect 239996 639236 240060 639300
rect 242756 639236 242820 639300
rect 244044 639296 244108 639300
rect 244044 639240 244058 639296
rect 244058 639240 244108 639296
rect 244044 639236 244108 639240
rect 247540 639236 247604 639300
rect 249012 639236 249076 639300
rect 252324 639296 252388 639300
rect 252324 639240 252338 639296
rect 252338 639240 252388 639296
rect 252324 639236 252388 639240
rect 255084 639236 255148 639300
rect 257844 639236 257908 639300
rect 261340 639236 261404 639300
rect 263364 639236 263428 639300
rect 273116 639296 273180 639300
rect 273116 639240 273166 639296
rect 273166 639240 273180 639296
rect 273116 639236 273180 639240
rect 281212 639296 281276 639300
rect 281212 639240 281226 639296
rect 281226 639240 281276 639296
rect 281212 639236 281276 639240
rect 307524 639236 307588 639300
rect 342668 639236 342732 639300
rect 362172 639236 362236 639300
rect 365116 639236 365180 639300
rect 315988 639100 316052 639164
rect 325556 639100 325620 639164
rect 333284 639100 333348 639164
rect 336412 639100 336476 639164
rect 342484 639100 342548 639164
rect 355548 639100 355612 639164
rect 364196 639100 364260 639164
rect 257660 638964 257724 639028
rect 229876 638828 229940 638892
rect 277164 638964 277228 639028
rect 277532 638964 277596 639028
rect 286916 638964 286980 639028
rect 267780 638828 267844 638892
rect 277348 638828 277412 638892
rect 286732 638828 286796 638892
rect 335308 638964 335372 639028
rect 355180 638964 355244 639028
rect 362356 638964 362420 639028
rect 374868 639100 374932 639164
rect 384068 639100 384132 639164
rect 398604 639100 398668 639164
rect 398972 639100 399036 639164
rect 408540 639236 408604 639300
rect 408724 639236 408788 639300
rect 417740 639508 417804 639572
rect 422708 639508 422772 639572
rect 462268 639296 462332 639300
rect 462268 639240 462318 639296
rect 462318 639240 462332 639296
rect 462268 639236 462332 639240
rect 488580 639296 488644 639300
rect 488580 639240 488630 639296
rect 488630 639240 488644 639296
rect 488580 639236 488644 639240
rect 509740 639296 509804 639300
rect 509740 639240 509790 639296
rect 509790 639240 509804 639296
rect 509740 639236 509804 639240
rect 525380 639296 525444 639300
rect 525380 639240 525430 639296
rect 525430 639240 525444 639296
rect 525380 639236 525444 639240
rect 527220 639236 527284 639300
rect 342484 638828 342548 638892
rect 342668 638828 342732 638892
rect 374500 638964 374564 639028
rect 384436 638828 384500 638892
rect 333284 638556 333348 638620
rect 234292 638420 234356 638484
rect 239444 638420 239508 638484
rect 244228 638420 244292 638484
rect 258028 638420 258092 638484
rect 267596 638420 267660 638484
rect 277532 638420 277596 638484
rect 286732 638420 286796 638484
rect 296668 638420 296732 638484
rect 306604 638420 306668 638484
rect 315988 638420 316052 638484
rect 325556 638420 325620 638484
rect 335308 638420 335372 638484
rect 355180 638692 355244 638756
rect 355364 638692 355428 638756
rect 362172 638692 362236 638756
rect 362356 638692 362420 638756
rect 374500 638692 374564 638756
rect 374684 638692 374748 638756
rect 384252 638692 384316 638756
rect 402836 638964 402900 639028
rect 384804 638828 384868 638892
rect 384988 638828 385052 638892
rect 408540 638964 408604 639028
rect 408356 638828 408420 638892
rect 408540 638828 408604 638892
rect 437244 638964 437308 639028
rect 408724 638692 408788 638756
rect 417924 638828 417988 638892
rect 437428 638828 437492 638892
rect 422708 638692 422772 638756
rect 437244 638692 437308 638756
rect 456564 638964 456628 639028
rect 437796 638828 437860 638892
rect 456564 638692 456628 638756
rect 336412 638556 336476 638620
rect 355364 638420 355428 638484
rect 355548 638420 355612 638484
rect 364196 638420 364260 638484
rect 462268 638556 462332 638620
rect 365116 638420 365180 638484
rect 374684 638420 374748 638484
rect 374868 638420 374932 638484
rect 384068 638420 384132 638484
rect 384252 638420 384316 638484
rect 417740 638420 417804 638484
rect 417924 638420 417988 638484
rect 488580 638420 488644 638484
rect 525196 638420 525260 638484
rect 529060 638420 529124 638484
rect 509740 638284 509804 638348
rect 525564 638284 525628 638348
rect 525380 638148 525444 638212
rect 229876 638012 229940 638076
rect 257660 638012 257724 638076
rect 258028 638012 258092 638076
rect 267596 638012 267660 638076
rect 273116 638012 273180 638076
rect 525196 638012 525260 638076
rect 234292 637876 234356 637940
rect 239444 637876 239508 637940
rect 244228 637876 244292 637940
rect 267780 637876 267844 637940
rect 277164 637876 277228 637940
rect 281212 637876 281276 637940
rect 277348 637740 277412 637804
rect 286916 637740 286980 637804
rect 296668 637740 296732 637804
rect 306604 637740 306668 637804
rect 307524 637740 307588 637804
rect 525564 637740 525628 637804
rect 527588 637468 527652 637532
rect 528140 637332 528204 637396
rect 528140 628084 528204 628148
rect 527404 627948 527468 628012
rect 527404 621012 527468 621076
rect 528324 621012 528388 621076
rect 528324 618156 528388 618220
rect 528876 618020 528940 618084
rect 528508 608636 528572 608700
rect 528876 608636 528940 608700
rect 527588 601700 527652 601764
rect 528508 601700 528572 601764
rect 527588 592180 527652 592244
rect 527588 591908 527652 591972
rect 527404 589460 527468 589524
rect 527588 589460 527652 589524
rect 527220 570420 527284 570484
rect 527588 570148 527652 570212
rect 527220 570012 527284 570076
rect 527404 570012 527468 570076
rect 527404 568516 527468 568580
rect 528140 568516 528204 568580
rect 528140 559132 528204 559196
rect 527588 558996 527652 559060
rect 527588 553964 527652 554028
rect 527956 553692 528020 553756
rect 527956 553284 528020 553348
rect 527588 553012 527652 553076
rect 527588 533700 527652 533764
rect 527588 514796 527652 514860
rect 527588 514660 527652 514724
rect 527588 512212 527652 512276
rect 527772 512076 527836 512140
rect 527772 505140 527836 505204
rect 527404 504868 527468 504932
rect 527772 492492 527836 492556
rect 528140 492356 528204 492420
rect 527588 482972 527652 483036
rect 528140 482972 528204 483036
rect 527588 471820 527652 471884
rect 527956 471684 528020 471748
rect 527956 462300 528020 462364
rect 528140 462300 528204 462364
rect 527772 454004 527836 454068
rect 528140 454004 528204 454068
rect 527772 447204 527836 447268
rect 527588 446932 527652 446996
rect 527220 428300 527284 428364
rect 527772 428300 527836 428364
rect 527588 425036 527652 425100
rect 527588 424900 527652 424964
rect 527220 421636 527284 421700
rect 527772 421636 527836 421700
rect 527588 368732 527652 368796
rect 234292 336636 234356 336700
rect 234660 327116 234724 327180
rect 258948 324260 259012 324324
rect 234660 318956 234724 319020
rect 234292 318820 234356 318884
rect 234292 303104 234356 303108
rect 234292 303048 234306 303104
rect 234306 303048 234356 303104
rect 234292 303044 234356 303048
rect 234292 299508 234356 299572
rect 234292 290396 234356 290460
rect 234660 290396 234724 290460
rect 529060 274620 529124 274684
rect 234476 273396 234540 273460
rect 234108 273260 234172 273324
rect 261892 266188 261956 266252
rect 234108 263740 234172 263804
rect 233924 263468 233988 263532
rect 233924 262108 233988 262172
rect 234108 252588 234172 252652
rect 261708 252452 261772 252516
rect 234108 247692 234172 247756
rect 234476 247692 234540 247756
rect 234476 225116 234540 225180
rect 234292 224844 234356 224908
rect 263364 208524 263428 208588
rect 261524 208252 261588 208316
rect 234476 206892 234540 206956
rect 362908 204716 362972 204780
rect 372476 204716 372540 204780
rect 362908 204444 362972 204508
rect 372476 204444 372540 204508
rect 463372 204716 463436 204780
rect 502012 204716 502076 204780
rect 531268 204716 531332 204780
rect 463556 204308 463620 204372
rect 502196 204308 502260 204372
rect 531268 204444 531332 204508
rect 550588 204444 550652 204508
rect 550588 204172 550652 204236
rect 359044 200228 359108 200292
rect 359044 198792 359108 198796
rect 359044 198736 359094 198792
rect 359094 198736 359108 198792
rect 359044 198732 359108 198736
rect 234292 197372 234356 197436
rect 234292 187716 234356 187780
rect 234476 187716 234540 187780
rect 234476 187504 234540 187508
rect 234476 187448 234526 187504
rect 234526 187448 234540 187504
rect 234476 187444 234540 187448
rect 343588 181384 343652 181388
rect 343588 181328 343602 181384
rect 343602 181328 343652 181384
rect 343588 181324 343652 181328
rect 257844 180916 257908 180980
rect 318748 181052 318812 181116
rect 343588 181052 343652 181116
rect 318748 180780 318812 180844
rect 361620 180916 361684 180980
rect 463556 181052 463620 181116
rect 463556 180780 463620 180844
rect 531268 181188 531332 181252
rect 502196 181052 502260 181116
rect 502196 180780 502260 180844
rect 531268 180916 531332 180980
rect 258764 180644 258828 180708
rect 361620 180644 361684 180708
rect 234660 178060 234724 178124
rect 265204 177304 265268 177308
rect 265204 177248 265254 177304
rect 265254 177248 265268 177304
rect 265204 177244 265268 177248
rect 261340 171260 261404 171324
rect 531268 170172 531332 170236
rect 531268 169900 531332 169964
rect 550588 169900 550652 169964
rect 550588 169628 550652 169692
rect 234292 164188 234356 164252
rect 234660 164188 234724 164252
rect 265204 164248 265268 164252
rect 265204 164192 265254 164248
rect 265254 164192 265268 164248
rect 265204 164188 265268 164192
rect 307708 157796 307772 157860
rect 384988 157796 385052 157860
rect 255084 157524 255148 157588
rect 299428 157524 299492 157588
rect 299428 157388 299492 157452
rect 307708 157388 307772 157452
rect 502012 157796 502076 157860
rect 531268 157796 531332 157860
rect 502196 157388 502260 157452
rect 531268 157524 531332 157588
rect 384804 157252 384868 157316
rect 550588 157524 550652 157588
rect 550588 157252 550652 157316
rect 234292 154532 234356 154596
rect 234476 154532 234540 154596
rect 258580 151676 258644 151740
rect 234292 144876 234356 144940
rect 234476 144876 234540 144940
rect 234292 138680 234356 138684
rect 234292 138624 234342 138680
rect 234342 138624 234356 138680
rect 234292 138620 234356 138624
rect 392164 138272 392228 138276
rect 392164 138216 392214 138272
rect 392214 138216 392228 138272
rect 392164 138212 392228 138216
rect 392164 135280 392228 135284
rect 392164 135224 392178 135280
rect 392178 135224 392228 135280
rect 392164 135220 392228 135224
rect 324268 134404 324332 134468
rect 249012 133860 249076 133924
rect 318748 133996 318812 134060
rect 285628 133860 285692 133924
rect 318748 133724 318812 133788
rect 324268 134132 324332 134196
rect 357388 133860 357452 133924
rect 393268 134132 393332 134196
rect 393268 133860 393332 133924
rect 473308 133996 473372 134060
rect 531268 134268 531332 134332
rect 502196 134132 502260 134196
rect 285628 133588 285692 133652
rect 357388 133588 357452 133652
rect 473308 133588 473372 133652
rect 502196 133860 502260 133924
rect 531268 133996 531332 134060
rect 550588 133996 550652 134060
rect 550588 133724 550652 133788
rect 249932 125896 249996 125900
rect 249932 125840 249982 125896
rect 249982 125840 249996 125896
rect 249932 125836 249996 125840
rect 249932 125624 249996 125628
rect 249932 125568 249982 125624
rect 249982 125568 249996 125624
rect 249932 125564 249996 125568
rect 359044 124068 359108 124132
rect 365668 123388 365732 123452
rect 307708 123252 307772 123316
rect 252324 123116 252388 123180
rect 335308 123116 335372 123180
rect 307708 122980 307772 123044
rect 365668 122980 365732 123044
rect 335308 122844 335372 122908
rect 531268 123252 531332 123316
rect 531268 122980 531332 123044
rect 550588 122980 550652 123044
rect 550588 122708 550652 122772
rect 234476 121620 234540 121684
rect 234660 121408 234724 121412
rect 234660 121352 234710 121408
rect 234710 121352 234724 121408
rect 234660 121348 234724 121352
rect 359044 114548 359108 114612
rect 234660 112976 234724 112980
rect 234660 112920 234710 112976
rect 234710 112920 234724 112976
rect 234660 112916 234724 112920
rect 327028 111012 327092 111076
rect 247540 110604 247604 110668
rect 298140 110604 298204 110668
rect 298140 110468 298204 110532
rect 327028 110740 327092 110804
rect 357388 110740 357452 110804
rect 357572 110468 357636 110532
rect 463372 110876 463436 110940
rect 502012 110876 502076 110940
rect 531268 110876 531332 110940
rect 463556 110468 463620 110532
rect 502196 110468 502260 110532
rect 531268 110604 531332 110668
rect 550588 110604 550652 110668
rect 550588 110332 550652 110396
rect 451596 99512 451660 99516
rect 451596 99456 451646 99512
rect 451646 99456 451660 99512
rect 451596 99452 451660 99456
rect 234292 96596 234356 96660
rect 234476 96596 234540 96660
rect 451596 96656 451660 96660
rect 451596 96600 451646 96656
rect 451646 96600 451660 96656
rect 451596 96596 451660 96600
rect 234476 89796 234540 89860
rect 234292 89524 234356 89588
rect 550588 87484 550652 87548
rect 242756 87076 242820 87140
rect 299428 87348 299492 87412
rect 317460 87348 317524 87412
rect 384988 87272 385052 87276
rect 384988 87216 385002 87272
rect 385002 87216 385052 87272
rect 384988 87212 385052 87216
rect 385172 87212 385236 87276
rect 299428 87076 299492 87140
rect 317460 87076 317524 87140
rect 375420 87076 375484 87140
rect 463556 87212 463620 87276
rect 463556 86940 463620 87004
rect 502196 87212 502260 87276
rect 502196 86940 502260 87004
rect 520228 86940 520292 87004
rect 550588 87076 550652 87140
rect 375420 86804 375484 86868
rect 520228 86668 520292 86732
rect 234292 80684 234356 80748
rect 234660 80684 234724 80748
rect 244044 75924 244108 75988
rect 234476 75788 234540 75852
rect 234660 75788 234724 75852
rect 357388 76332 357452 76396
rect 357388 76060 357452 76124
rect 376708 76060 376772 76124
rect 376892 76060 376956 76124
rect 531268 76332 531332 76396
rect 531268 76060 531332 76124
rect 550588 76060 550652 76124
rect 550588 75788 550652 75852
rect 239996 64968 240060 64972
rect 239996 64912 240046 64968
rect 240046 64912 240060 64968
rect 239996 64908 240060 64912
rect 309180 63548 309244 63612
rect 309180 63276 309244 63340
rect 373948 63684 374012 63748
rect 502012 63956 502076 64020
rect 531268 63956 531332 64020
rect 502196 63548 502260 63612
rect 531268 63684 531332 63748
rect 373948 63412 374012 63476
rect 550588 63684 550652 63748
rect 550588 63412 550652 63476
rect 234108 43828 234172 43892
rect 258028 40428 258092 40492
rect 258028 40020 258092 40084
rect 335308 40020 335372 40084
rect 383700 40292 383764 40356
rect 383700 40020 383764 40084
rect 531268 40428 531332 40492
rect 502196 40292 502260 40356
rect 502196 40020 502260 40084
rect 531268 40156 531332 40220
rect 335308 39748 335372 39812
rect 550588 40156 550652 40220
rect 550588 39884 550652 39948
rect 338068 29548 338132 29612
rect 237236 29276 237300 29340
rect 373948 29548 374012 29612
rect 453988 29548 454052 29612
rect 550588 29548 550652 29612
rect 288388 29140 288452 29204
rect 318748 29336 318812 29340
rect 318748 29280 318762 29336
rect 318762 29280 318812 29336
rect 318748 29276 318812 29280
rect 307708 29140 307772 29204
rect 338068 29276 338132 29340
rect 373948 29336 374012 29340
rect 373948 29280 373962 29336
rect 373962 29280 374012 29336
rect 373948 29276 374012 29280
rect 318748 29004 318812 29068
rect 288388 28868 288452 28932
rect 307708 28868 307772 28932
rect 463556 29412 463620 29476
rect 453988 29140 454052 29204
rect 463556 29004 463620 29068
rect 502196 29412 502260 29476
rect 521516 29412 521580 29476
rect 531268 29412 531332 29476
rect 502196 29004 502260 29068
rect 531268 29140 531332 29204
rect 521516 29004 521580 29068
rect 550588 29140 550652 29204
rect 527220 21932 527284 21996
rect 259500 17308 259564 17372
rect 268884 17308 268948 17372
rect 357388 17172 357452 17236
rect 259500 17036 259564 17100
rect 367140 17036 367204 17100
rect 231716 16764 231780 16828
rect 269068 16492 269132 16556
rect 306420 16900 306484 16964
rect 357388 16900 357452 16964
rect 425100 17036 425164 17100
rect 306604 16628 306668 16692
rect 367140 16764 367204 16828
rect 425100 16764 425164 16828
rect 502012 17036 502076 17100
rect 531268 17036 531332 17100
rect 502196 16628 502260 16692
rect 531268 16764 531332 16828
rect 550588 16764 550652 16828
rect 550588 16492 550652 16556
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 231715 639300 231781 639301
rect 231715 639236 231716 639300
rect 231780 639236 231781 639300
rect 231715 639235 231781 639236
rect 234475 639300 234541 639301
rect 234475 639236 234476 639300
rect 234540 639236 234541 639300
rect 234475 639235 234541 639236
rect 229875 638892 229941 638893
rect 229875 638828 229876 638892
rect 229940 638828 229941 638892
rect 229875 638827 229941 638828
rect 229878 638077 229938 638827
rect 229875 638076 229941 638077
rect 229875 638012 229876 638076
rect 229940 638012 229941 638076
rect 229875 638011 229941 638012
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 231718 16829 231778 639235
rect 234291 638484 234357 638485
rect 234291 638420 234292 638484
rect 234356 638420 234357 638484
rect 234291 638419 234357 638420
rect 234294 637941 234354 638419
rect 234291 637940 234357 637941
rect 234291 637876 234292 637940
rect 234356 637876 234357 637940
rect 234291 637875 234357 637876
rect 234478 529498 234538 639235
rect 234804 632454 235404 667898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 237235 639300 237301 639301
rect 237235 639236 237236 639300
rect 237300 639236 237301 639300
rect 237235 639235 237301 639236
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234478 490738 234538 520422
rect 233558 481898 233618 490502
rect 234804 488454 235404 523898
rect 235582 520658 235642 529262
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234478 394178 234538 481662
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234478 356098 234538 385102
rect 234804 380454 235404 415898
rect 235582 385338 235642 393942
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 233558 346578 233618 355862
rect 234478 341730 234538 346342
rect 234110 341670 234538 341730
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234110 340370 234170 341670
rect 234110 340310 234354 340370
rect 234294 336701 234354 340310
rect 234291 336700 234357 336701
rect 234291 336636 234292 336700
rect 234356 336636 234357 336700
rect 234291 336635 234357 336636
rect 234659 327180 234725 327181
rect 234659 327116 234660 327180
rect 234724 327116 234725 327180
rect 234659 327115 234725 327116
rect 234662 319021 234722 327115
rect 234659 319020 234725 319021
rect 234659 318956 234660 319020
rect 234724 318956 234725 319020
rect 234659 318955 234725 318956
rect 234291 318884 234357 318885
rect 234291 318820 234292 318884
rect 234356 318820 234357 318884
rect 234291 318819 234357 318820
rect 234294 303109 234354 318819
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234291 303108 234357 303109
rect 234291 303044 234292 303108
rect 234356 303044 234357 303108
rect 234291 303043 234357 303044
rect 234291 299572 234357 299573
rect 234291 299508 234292 299572
rect 234356 299508 234357 299572
rect 234291 299507 234357 299508
rect 234294 290461 234354 299507
rect 234291 290460 234357 290461
rect 234291 290396 234292 290460
rect 234356 290396 234357 290460
rect 234291 290395 234357 290396
rect 234659 290460 234725 290461
rect 234659 290396 234660 290460
rect 234724 290396 234725 290460
rect 234659 290395 234725 290396
rect 234662 279170 234722 290395
rect 234478 279110 234722 279170
rect 234478 273461 234538 279110
rect 234475 273460 234541 273461
rect 234475 273396 234476 273460
rect 234540 273396 234541 273460
rect 234475 273395 234541 273396
rect 234107 273324 234173 273325
rect 234107 273260 234108 273324
rect 234172 273260 234173 273324
rect 234107 273259 234173 273260
rect 234110 263805 234170 273259
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234107 263804 234173 263805
rect 234107 263740 234108 263804
rect 234172 263740 234173 263804
rect 234107 263739 234173 263740
rect 233923 263532 233989 263533
rect 233923 263468 233924 263532
rect 233988 263468 233989 263532
rect 233923 263467 233989 263468
rect 233926 262173 233986 263467
rect 233923 262172 233989 262173
rect 233923 262108 233924 262172
rect 233988 262108 233989 262172
rect 233923 262107 233989 262108
rect 234107 252652 234173 252653
rect 234107 252588 234108 252652
rect 234172 252588 234173 252652
rect 234107 252587 234173 252588
rect 234110 247757 234170 252587
rect 234107 247756 234173 247757
rect 234107 247692 234108 247756
rect 234172 247692 234173 247756
rect 234107 247691 234173 247692
rect 234475 247756 234541 247757
rect 234475 247692 234476 247756
rect 234540 247692 234541 247756
rect 234475 247691 234541 247692
rect 234478 225181 234538 247691
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234475 225180 234541 225181
rect 234475 225116 234476 225180
rect 234540 225116 234541 225180
rect 234475 225115 234541 225116
rect 234291 224908 234357 224909
rect 234291 224844 234292 224908
rect 234356 224844 234357 224908
rect 234291 224843 234357 224844
rect 234294 215930 234354 224843
rect 234294 215870 234538 215930
rect 234478 206957 234538 215870
rect 234475 206956 234541 206957
rect 234475 206892 234476 206956
rect 234540 206892 234541 206956
rect 234475 206891 234541 206892
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234291 197436 234357 197437
rect 234291 197372 234292 197436
rect 234356 197372 234357 197436
rect 234291 197371 234357 197372
rect 234294 187781 234354 197371
rect 234291 187780 234357 187781
rect 234291 187716 234292 187780
rect 234356 187716 234357 187780
rect 234291 187715 234357 187716
rect 234475 187780 234541 187781
rect 234475 187716 234476 187780
rect 234540 187716 234541 187780
rect 234475 187715 234541 187716
rect 234478 187509 234538 187715
rect 234475 187508 234541 187509
rect 234475 187444 234476 187508
rect 234540 187444 234541 187508
rect 234475 187443 234541 187444
rect 234659 178124 234725 178125
rect 234659 178060 234660 178124
rect 234724 178060 234725 178124
rect 234659 178059 234725 178060
rect 234662 164253 234722 178059
rect 234804 164454 235404 199898
rect 234291 164252 234357 164253
rect 234291 164188 234292 164252
rect 234356 164188 234357 164252
rect 234291 164187 234357 164188
rect 234659 164252 234725 164253
rect 234659 164188 234660 164252
rect 234724 164188 234725 164252
rect 234659 164187 234725 164188
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234294 154597 234354 164187
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234291 154596 234357 154597
rect 234291 154532 234292 154596
rect 234356 154532 234357 154596
rect 234291 154531 234357 154532
rect 234475 154596 234541 154597
rect 234475 154532 234476 154596
rect 234540 154532 234541 154596
rect 234475 154531 234541 154532
rect 234478 144941 234538 154531
rect 234291 144940 234357 144941
rect 234291 144876 234292 144940
rect 234356 144876 234357 144940
rect 234291 144875 234357 144876
rect 234475 144940 234541 144941
rect 234475 144876 234476 144940
rect 234540 144876 234541 144940
rect 234475 144875 234541 144876
rect 234294 138685 234354 144875
rect 234291 138684 234357 138685
rect 234291 138620 234292 138684
rect 234356 138620 234357 138684
rect 234291 138619 234357 138620
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234475 121684 234541 121685
rect 234475 121620 234476 121684
rect 234540 121620 234541 121684
rect 234475 121619 234541 121620
rect 234478 121410 234538 121619
rect 234659 121412 234725 121413
rect 234659 121410 234660 121412
rect 234478 121350 234660 121410
rect 234659 121348 234660 121350
rect 234724 121348 234725 121412
rect 234659 121347 234725 121348
rect 234659 112980 234725 112981
rect 234659 112916 234660 112980
rect 234724 112916 234725 112980
rect 234659 112915 234725 112916
rect 234662 108490 234722 112915
rect 234294 108430 234722 108490
rect 234294 96661 234354 108430
rect 234291 96660 234357 96661
rect 234291 96596 234292 96660
rect 234356 96596 234357 96660
rect 234291 96595 234357 96596
rect 234475 96660 234541 96661
rect 234475 96596 234476 96660
rect 234540 96596 234541 96660
rect 234475 96595 234541 96596
rect 234478 89861 234538 96595
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234475 89860 234541 89861
rect 234475 89796 234476 89860
rect 234540 89796 234541 89860
rect 234475 89795 234541 89796
rect 234291 89588 234357 89589
rect 234291 89524 234292 89588
rect 234356 89524 234357 89588
rect 234291 89523 234357 89524
rect 234294 80749 234354 89523
rect 234291 80748 234357 80749
rect 234291 80684 234292 80748
rect 234356 80684 234357 80748
rect 234291 80683 234357 80684
rect 234659 80748 234725 80749
rect 234659 80684 234660 80748
rect 234724 80684 234725 80748
rect 234659 80683 234725 80684
rect 234662 75853 234722 80683
rect 234475 75852 234541 75853
rect 234475 75788 234476 75852
rect 234540 75788 234541 75852
rect 234475 75787 234541 75788
rect 234659 75852 234725 75853
rect 234659 75788 234660 75852
rect 234724 75788 234725 75852
rect 234659 75787 234725 75788
rect 234478 51370 234538 75787
rect 234110 51310 234538 51370
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234110 43893 234170 51310
rect 234107 43892 234173 43893
rect 234107 43828 234108 43892
rect 234172 43828 234173 43892
rect 234107 43827 234173 43828
rect 234804 20454 235404 55898
rect 237238 29341 237298 639235
rect 238404 636054 239004 671498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 239995 639300 240061 639301
rect 239995 639236 239996 639300
rect 240060 639236 240061 639300
rect 239995 639235 240061 639236
rect 239443 638484 239509 638485
rect 239443 638420 239444 638484
rect 239508 638420 239509 638484
rect 239443 638419 239509 638420
rect 239446 637941 239506 638419
rect 239443 637940 239509 637941
rect 239443 637876 239444 637940
rect 239508 637876 239509 637940
rect 239443 637875 239509 637876
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 239998 64973 240058 639235
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 242755 639300 242821 639301
rect 242755 639236 242756 639300
rect 242820 639236 242821 639300
rect 242755 639235 242821 639236
rect 244043 639300 244109 639301
rect 244043 639236 244044 639300
rect 244108 639236 244109 639300
rect 244043 639235 244109 639236
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 239995 64972 240061 64973
rect 239995 64908 239996 64972
rect 240060 64908 240061 64972
rect 239995 64907 240061 64908
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 237235 29340 237301 29341
rect 237235 29276 237236 29340
rect 237300 29276 237301 29340
rect 237235 29275 237301 29276
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 231715 16828 231781 16829
rect 231715 16764 231716 16828
rect 231780 16764 231781 16828
rect 231715 16763 231781 16764
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 63654 242604 99098
rect 242758 87141 242818 639235
rect 242755 87140 242821 87141
rect 242755 87076 242756 87140
rect 242820 87076 242821 87140
rect 242755 87075 242821 87076
rect 244046 75989 244106 639235
rect 244227 638484 244293 638485
rect 244227 638420 244228 638484
rect 244292 638420 244293 638484
rect 244227 638419 244293 638420
rect 244230 637941 244290 638419
rect 244227 637940 244293 637941
rect 244227 637876 244228 637940
rect 244292 637876 244293 637940
rect 244227 637875 244293 637876
rect 245604 607254 246204 642698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 247539 639300 247605 639301
rect 247539 639236 247540 639300
rect 247604 639236 247605 639300
rect 247539 639235 247605 639236
rect 249011 639300 249077 639301
rect 249011 639236 249012 639300
rect 249076 639236 249077 639300
rect 249011 639235 249077 639236
rect 252323 639300 252389 639301
rect 252323 639236 252324 639300
rect 252388 639236 252389 639300
rect 252323 639235 252389 639236
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 247542 110669 247602 639235
rect 249014 133925 249074 639235
rect 249011 133924 249077 133925
rect 249011 133860 249012 133924
rect 249076 133860 249077 133924
rect 249011 133859 249077 133860
rect 249931 125900 249997 125901
rect 249931 125836 249932 125900
rect 249996 125836 249997 125900
rect 249931 125835 249997 125836
rect 249934 125629 249994 125835
rect 249931 125628 249997 125629
rect 249931 125564 249932 125628
rect 249996 125564 249997 125628
rect 249931 125563 249997 125564
rect 252326 123181 252386 639235
rect 252804 614454 253404 649898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 255083 639300 255149 639301
rect 255083 639236 255084 639300
rect 255148 639236 255149 639300
rect 255083 639235 255149 639236
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 255086 157589 255146 639235
rect 256404 618054 257004 653498
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 258947 642700 259013 642701
rect 258947 642636 258948 642700
rect 259012 642636 259013 642700
rect 258947 642635 259013 642636
rect 258763 642156 258829 642157
rect 258763 642092 258764 642156
rect 258828 642092 258829 642156
rect 258763 642091 258829 642092
rect 258579 641884 258645 641885
rect 258579 641820 258580 641884
rect 258644 641820 258645 641884
rect 258579 641819 258645 641820
rect 257843 639300 257909 639301
rect 257843 639236 257844 639300
rect 257908 639236 257909 639300
rect 257843 639235 257909 639236
rect 257659 639028 257725 639029
rect 257659 638964 257660 639028
rect 257724 638964 257725 639028
rect 257659 638963 257725 638964
rect 257662 638077 257722 638963
rect 257659 638076 257725 638077
rect 257659 638012 257660 638076
rect 257724 638012 257725 638076
rect 257659 638011 257725 638012
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 255083 157588 255149 157589
rect 255083 157524 255084 157588
rect 255148 157524 255149 157588
rect 255083 157523 255149 157524
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252323 123180 252389 123181
rect 252323 123116 252324 123180
rect 252388 123116 252389 123180
rect 252323 123115 252389 123116
rect 247539 110668 247605 110669
rect 247539 110604 247540 110668
rect 247604 110604 247605 110668
rect 247539 110603 247605 110604
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 244043 75988 244109 75989
rect 244043 75924 244044 75988
rect 244108 75924 244109 75988
rect 244043 75923 244109 75924
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 150054 257004 185498
rect 257846 180981 257906 639235
rect 258027 638484 258093 638485
rect 258027 638420 258028 638484
rect 258092 638420 258093 638484
rect 258027 638419 258093 638420
rect 258030 638077 258090 638419
rect 258027 638076 258093 638077
rect 258027 638012 258028 638076
rect 258092 638012 258093 638076
rect 258027 638011 258093 638012
rect 257843 180980 257909 180981
rect 257843 180916 257844 180980
rect 257908 180916 257909 180980
rect 257843 180915 257909 180916
rect 258582 151741 258642 641819
rect 258766 180709 258826 642091
rect 258950 324325 259010 642635
rect 260004 621654 260604 657098
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 261891 642564 261957 642565
rect 261891 642500 261892 642564
rect 261956 642500 261957 642564
rect 261891 642499 261957 642500
rect 261707 642428 261773 642429
rect 261707 642364 261708 642428
rect 261772 642364 261773 642428
rect 261707 642363 261773 642364
rect 261523 642292 261589 642293
rect 261523 642228 261524 642292
rect 261588 642228 261589 642292
rect 261523 642227 261589 642228
rect 261339 639300 261405 639301
rect 261339 639236 261340 639300
rect 261404 639236 261405 639300
rect 261339 639235 261405 639236
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 258947 324324 259013 324325
rect 258947 324260 258948 324324
rect 259012 324260 259013 324324
rect 258947 324259 259013 324260
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 258763 180708 258829 180709
rect 258763 180644 258764 180708
rect 258828 180644 258829 180708
rect 258763 180643 258829 180644
rect 260004 153654 260604 189098
rect 261342 171325 261402 639235
rect 261526 208317 261586 642227
rect 261710 252517 261770 642363
rect 261894 266253 261954 642499
rect 263363 639300 263429 639301
rect 263363 639236 263364 639300
rect 263428 639236 263429 639300
rect 263363 639235 263429 639236
rect 261891 266252 261957 266253
rect 261891 266188 261892 266252
rect 261956 266188 261957 266252
rect 261891 266187 261957 266188
rect 261707 252516 261773 252517
rect 261707 252452 261708 252516
rect 261772 252452 261773 252516
rect 261707 252451 261773 252452
rect 263366 208589 263426 639235
rect 263604 625254 264204 660698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 267779 638892 267845 638893
rect 267779 638828 267780 638892
rect 267844 638828 267845 638892
rect 267779 638827 267845 638828
rect 267595 638484 267661 638485
rect 267595 638420 267596 638484
rect 267660 638420 267661 638484
rect 267595 638419 267661 638420
rect 267598 638077 267658 638419
rect 267595 638076 267661 638077
rect 267595 638012 267596 638076
rect 267660 638012 267661 638076
rect 267595 638011 267661 638012
rect 267782 637941 267842 638827
rect 267779 637940 267845 637941
rect 267779 637876 267780 637940
rect 267844 637876 267845 637940
rect 267779 637875 267845 637876
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263363 208588 263429 208589
rect 263363 208524 263364 208588
rect 263428 208524 263429 208588
rect 263363 208523 263429 208524
rect 261523 208316 261589 208317
rect 261523 208252 261524 208316
rect 261588 208252 261589 208316
rect 261523 208251 261589 208252
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 261339 171324 261405 171325
rect 261339 171260 261340 171324
rect 261404 171260 261405 171324
rect 261339 171259 261405 171260
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 258579 151740 258645 151741
rect 258579 151676 258580 151740
rect 258644 151676 258645 151740
rect 258579 151675 258645 151676
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 258027 40492 258093 40493
rect 258027 40428 258028 40492
rect 258092 40428 258093 40492
rect 258027 40427 258093 40428
rect 258030 40085 258090 40427
rect 258027 40084 258093 40085
rect 258027 40020 258028 40084
rect 258092 40020 258093 40084
rect 258027 40019 258093 40020
rect 259499 17372 259565 17373
rect 259499 17308 259500 17372
rect 259564 17308 259565 17372
rect 259499 17307 259565 17308
rect 259502 17101 259562 17307
rect 259499 17100 259565 17101
rect 259499 17036 259500 17100
rect 259564 17036 259565 17100
rect 259499 17035 259565 17036
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 157254 264204 192698
rect 270804 632454 271404 667898
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 273115 639300 273181 639301
rect 273115 639236 273116 639300
rect 273180 639236 273181 639300
rect 273115 639235 273181 639236
rect 273118 638077 273178 639235
rect 273115 638076 273181 638077
rect 273115 638012 273116 638076
rect 273180 638012 273181 638076
rect 273115 638011 273181 638012
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 265203 177308 265269 177309
rect 265203 177244 265204 177308
rect 265268 177244 265269 177308
rect 265203 177243 265269 177244
rect 265206 164253 265266 177243
rect 270804 164454 271404 199898
rect 265203 164252 265269 164253
rect 265203 164188 265204 164252
rect 265268 164188 265269 164252
rect 265203 164187 265269 164188
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 268883 17372 268949 17373
rect 268883 17308 268884 17372
rect 268948 17308 268949 17372
rect 268883 17307 268949 17308
rect 268886 16690 268946 17307
rect 268886 16630 269130 16690
rect 269070 16557 269130 16630
rect 269067 16556 269133 16557
rect 269067 16492 269068 16556
rect 269132 16492 269133 16556
rect 269067 16491 269133 16492
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 636054 275004 671498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281211 639300 281277 639301
rect 281211 639236 281212 639300
rect 281276 639236 281277 639300
rect 281211 639235 281277 639236
rect 277163 639028 277229 639029
rect 277163 638964 277164 639028
rect 277228 638964 277229 639028
rect 277163 638963 277229 638964
rect 277531 639028 277597 639029
rect 277531 638964 277532 639028
rect 277596 638964 277597 639028
rect 277531 638963 277597 638964
rect 277166 637941 277226 638963
rect 277347 638892 277413 638893
rect 277347 638828 277348 638892
rect 277412 638828 277413 638892
rect 277347 638827 277413 638828
rect 277163 637940 277229 637941
rect 277163 637876 277164 637940
rect 277228 637876 277229 637940
rect 277163 637875 277229 637876
rect 277350 637805 277410 638827
rect 277534 638485 277594 638963
rect 277531 638484 277597 638485
rect 277531 638420 277532 638484
rect 277596 638420 277597 638484
rect 277531 638419 277597 638420
rect 277347 637804 277413 637805
rect 277347 637740 277348 637804
rect 277412 637740 277413 637804
rect 277347 637739 277413 637740
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 603654 278604 639098
rect 281214 637941 281274 639235
rect 281211 637940 281277 637941
rect 281211 637876 281212 637940
rect 281276 637876 281277 637940
rect 281211 637875 281277 637876
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 607254 282204 642698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 286915 639028 286981 639029
rect 286915 638964 286916 639028
rect 286980 638964 286981 639028
rect 286915 638963 286981 638964
rect 286731 638892 286797 638893
rect 286731 638828 286732 638892
rect 286796 638828 286797 638892
rect 286731 638827 286797 638828
rect 286734 638485 286794 638827
rect 286731 638484 286797 638485
rect 286731 638420 286732 638484
rect 286796 638420 286797 638484
rect 286731 638419 286797 638420
rect 286918 637805 286978 638963
rect 286915 637804 286981 637805
rect 286915 637740 286916 637804
rect 286980 637740 286981 637804
rect 286915 637739 286981 637740
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 285627 133924 285693 133925
rect 285627 133860 285628 133924
rect 285692 133860 285693 133924
rect 285627 133859 285693 133860
rect 285630 133653 285690 133859
rect 285627 133652 285693 133653
rect 285627 133588 285628 133652
rect 285692 133588 285693 133652
rect 285627 133587 285693 133588
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288387 29204 288453 29205
rect 288387 29140 288388 29204
rect 288452 29140 288453 29204
rect 288387 29139 288453 29140
rect 288390 28933 288450 29139
rect 288387 28932 288453 28933
rect 288387 28868 288388 28932
rect 288452 28868 288453 28932
rect 288387 28867 288453 28868
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 296667 638484 296733 638485
rect 296667 638420 296668 638484
rect 296732 638420 296733 638484
rect 296667 638419 296733 638420
rect 296670 637805 296730 638419
rect 296667 637804 296733 637805
rect 296667 637740 296668 637804
rect 296732 637740 296733 637804
rect 296667 637739 296733 637740
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 299604 625254 300204 660698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306603 638484 306669 638485
rect 306603 638420 306604 638484
rect 306668 638420 306669 638484
rect 306603 638419 306669 638420
rect 306606 637805 306666 638419
rect 306603 637804 306669 637805
rect 306603 637740 306604 637804
rect 306668 637740 306669 637804
rect 306603 637739 306669 637740
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299427 157588 299493 157589
rect 299427 157524 299428 157588
rect 299492 157524 299493 157588
rect 299427 157523 299493 157524
rect 299430 157453 299490 157523
rect 299427 157452 299493 157453
rect 299427 157388 299428 157452
rect 299492 157388 299493 157452
rect 299427 157387 299493 157388
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 298139 110668 298205 110669
rect 298139 110604 298140 110668
rect 298204 110604 298205 110668
rect 298139 110603 298205 110604
rect 298142 110533 298202 110603
rect 298139 110532 298205 110533
rect 298139 110468 298140 110532
rect 298204 110468 298205 110532
rect 298139 110467 298205 110468
rect 299427 87412 299493 87413
rect 299427 87348 299428 87412
rect 299492 87348 299493 87412
rect 299427 87347 299493 87348
rect 299430 87141 299490 87347
rect 299427 87140 299493 87141
rect 299427 87076 299428 87140
rect 299492 87076 299493 87140
rect 299427 87075 299493 87076
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 306804 632454 307404 667898
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 307523 639300 307589 639301
rect 307523 639236 307524 639300
rect 307588 639236 307589 639300
rect 307523 639235 307589 639236
rect 307526 637805 307586 639235
rect 307523 637804 307589 637805
rect 307523 637740 307524 637804
rect 307588 637740 307589 637804
rect 307523 637739 307589 637740
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 307707 157860 307773 157861
rect 307707 157796 307708 157860
rect 307772 157796 307773 157860
rect 307707 157795 307773 157796
rect 307710 157453 307770 157795
rect 307707 157452 307773 157453
rect 307707 157388 307708 157452
rect 307772 157388 307773 157452
rect 307707 157387 307773 157388
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 307707 123316 307773 123317
rect 307707 123252 307708 123316
rect 307772 123252 307773 123316
rect 307707 123251 307773 123252
rect 307710 123045 307770 123251
rect 307707 123044 307773 123045
rect 307707 122980 307708 123044
rect 307772 122980 307773 123044
rect 307707 122979 307773 122980
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 309179 63612 309245 63613
rect 309179 63548 309180 63612
rect 309244 63548 309245 63612
rect 309179 63547 309245 63548
rect 309182 63341 309242 63547
rect 309179 63340 309245 63341
rect 309179 63276 309180 63340
rect 309244 63276 309245 63340
rect 309179 63275 309245 63276
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 307707 29204 307773 29205
rect 307707 29140 307708 29204
rect 307772 29140 307773 29204
rect 307707 29139 307773 29140
rect 307710 28933 307770 29139
rect 307707 28932 307773 28933
rect 307707 28868 307708 28932
rect 307772 28868 307773 28932
rect 307707 28867 307773 28868
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306422 17310 306666 17370
rect 306422 16965 306482 17310
rect 306419 16964 306485 16965
rect 306419 16900 306420 16964
rect 306484 16900 306485 16964
rect 306419 16899 306485 16900
rect 306606 16693 306666 17310
rect 306603 16692 306669 16693
rect 306603 16628 306604 16692
rect 306668 16628 306669 16692
rect 306603 16627 306669 16628
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 315987 639164 316053 639165
rect 315987 639100 315988 639164
rect 316052 639100 316053 639164
rect 315987 639099 316053 639100
rect 314004 603654 314604 639098
rect 315990 638485 316050 639099
rect 315987 638484 316053 638485
rect 315987 638420 315988 638484
rect 316052 638420 316053 638484
rect 315987 638419 316053 638420
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 325555 639164 325621 639165
rect 325555 639100 325556 639164
rect 325620 639100 325621 639164
rect 325555 639099 325621 639100
rect 325558 638485 325618 639099
rect 325555 638484 325621 638485
rect 325555 638420 325556 638484
rect 325620 638420 325621 638484
rect 325555 638419 325621 638420
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 318747 181116 318813 181117
rect 318747 181052 318748 181116
rect 318812 181052 318813 181116
rect 318747 181051 318813 181052
rect 318750 180845 318810 181051
rect 318747 180844 318813 180845
rect 318747 180780 318748 180844
rect 318812 180780 318813 180844
rect 318747 180779 318813 180780
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324267 134468 324333 134469
rect 324267 134404 324268 134468
rect 324332 134404 324333 134468
rect 324267 134403 324333 134404
rect 324270 134197 324330 134403
rect 324267 134196 324333 134197
rect 324267 134132 324268 134196
rect 324332 134132 324333 134196
rect 324267 134131 324333 134132
rect 318747 134060 318813 134061
rect 318747 133996 318748 134060
rect 318812 133996 318813 134060
rect 318747 133995 318813 133996
rect 318750 133789 318810 133995
rect 318747 133788 318813 133789
rect 318747 133724 318748 133788
rect 318812 133724 318813 133788
rect 318747 133723 318813 133724
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317459 87412 317525 87413
rect 317459 87348 317460 87412
rect 317524 87348 317525 87412
rect 317459 87347 317525 87348
rect 317462 87141 317522 87347
rect 317459 87140 317525 87141
rect 317459 87076 317460 87140
rect 317524 87076 317525 87140
rect 317459 87075 317525 87076
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 110454 325404 145898
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 327027 111076 327093 111077
rect 327027 111012 327028 111076
rect 327092 111012 327093 111076
rect 327027 111011 327093 111012
rect 327030 110805 327090 111011
rect 327027 110804 327093 110805
rect 327027 110740 327028 110804
rect 327092 110740 327093 110804
rect 327027 110739 327093 110740
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 318747 29340 318813 29341
rect 318747 29276 318748 29340
rect 318812 29276 318813 29340
rect 318747 29275 318813 29276
rect 318750 29069 318810 29275
rect 318747 29068 318813 29069
rect 318747 29004 318748 29068
rect 318812 29004 318813 29068
rect 318747 29003 318813 29004
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 333283 639164 333349 639165
rect 333283 639100 333284 639164
rect 333348 639100 333349 639164
rect 333283 639099 333349 639100
rect 333286 638621 333346 639099
rect 335307 639028 335373 639029
rect 335307 638964 335308 639028
rect 335372 638964 335373 639028
rect 335307 638963 335373 638964
rect 333283 638620 333349 638621
rect 333283 638556 333284 638620
rect 333348 638556 333349 638620
rect 333283 638555 333349 638556
rect 335310 638485 335370 638963
rect 335307 638484 335373 638485
rect 335307 638420 335308 638484
rect 335372 638420 335373 638484
rect 335307 638419 335373 638420
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 335604 625254 336204 660698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342667 639300 342733 639301
rect 342667 639236 342668 639300
rect 342732 639236 342733 639300
rect 342667 639235 342733 639236
rect 336411 639164 336477 639165
rect 336411 639100 336412 639164
rect 336476 639100 336477 639164
rect 336411 639099 336477 639100
rect 342483 639164 342549 639165
rect 342483 639100 342484 639164
rect 342548 639100 342549 639164
rect 342483 639099 342549 639100
rect 336414 638621 336474 639099
rect 342486 638893 342546 639099
rect 342670 638893 342730 639235
rect 342483 638892 342549 638893
rect 342483 638828 342484 638892
rect 342548 638828 342549 638892
rect 342483 638827 342549 638828
rect 342667 638892 342733 638893
rect 342667 638828 342668 638892
rect 342732 638828 342733 638892
rect 342667 638827 342733 638828
rect 336411 638620 336477 638621
rect 336411 638556 336412 638620
rect 336476 638556 336477 638620
rect 336411 638555 336477 638556
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335307 123180 335373 123181
rect 335307 123116 335308 123180
rect 335372 123116 335373 123180
rect 335307 123115 335373 123116
rect 335310 122909 335370 123115
rect 335307 122908 335373 122909
rect 335307 122844 335308 122908
rect 335372 122844 335373 122908
rect 335307 122843 335373 122844
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335307 40084 335373 40085
rect 335307 40020 335308 40084
rect 335372 40020 335373 40084
rect 335307 40019 335373 40020
rect 335310 39813 335370 40019
rect 335307 39812 335373 39813
rect 335307 39748 335308 39812
rect 335372 39748 335373 39812
rect 335307 39747 335373 39748
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 13254 336204 48698
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 343587 181388 343653 181389
rect 343587 181324 343588 181388
rect 343652 181324 343653 181388
rect 343587 181323 343653 181324
rect 343590 181117 343650 181323
rect 343587 181116 343653 181117
rect 343587 181052 343588 181116
rect 343652 181052 343653 181116
rect 343587 181051 343653 181052
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 338067 29612 338133 29613
rect 338067 29548 338068 29612
rect 338132 29548 338133 29612
rect 338067 29547 338133 29548
rect 338070 29341 338130 29547
rect 338067 29340 338133 29341
rect 338067 29276 338068 29340
rect 338132 29276 338133 29340
rect 338067 29275 338133 29276
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 355547 639164 355613 639165
rect 355547 639100 355548 639164
rect 355612 639100 355613 639164
rect 355547 639099 355613 639100
rect 355179 639028 355245 639029
rect 355179 638964 355180 639028
rect 355244 638964 355245 639028
rect 355179 638963 355245 638964
rect 355182 638757 355242 638963
rect 355179 638756 355245 638757
rect 355179 638692 355180 638756
rect 355244 638692 355245 638756
rect 355179 638691 355245 638692
rect 355363 638756 355429 638757
rect 355363 638692 355364 638756
rect 355428 638692 355429 638756
rect 355363 638691 355429 638692
rect 355366 638485 355426 638691
rect 355550 638485 355610 639099
rect 355363 638484 355429 638485
rect 355363 638420 355364 638484
rect 355428 638420 355429 638484
rect 355363 638419 355429 638420
rect 355547 638484 355613 638485
rect 355547 638420 355548 638484
rect 355612 638420 355613 638484
rect 355547 638419 355613 638420
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 360804 614454 361404 649898
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 362171 639300 362237 639301
rect 362171 639236 362172 639300
rect 362236 639236 362237 639300
rect 362171 639235 362237 639236
rect 362174 638757 362234 639235
rect 364195 639164 364261 639165
rect 364195 639100 364196 639164
rect 364260 639100 364261 639164
rect 364195 639099 364261 639100
rect 362355 639028 362421 639029
rect 362355 638964 362356 639028
rect 362420 638964 362421 639028
rect 362355 638963 362421 638964
rect 362358 638757 362418 638963
rect 362171 638756 362237 638757
rect 362171 638692 362172 638756
rect 362236 638692 362237 638756
rect 362171 638691 362237 638692
rect 362355 638756 362421 638757
rect 362355 638692 362356 638756
rect 362420 638692 362421 638756
rect 362355 638691 362421 638692
rect 364198 638485 364258 639099
rect 364195 638484 364261 638485
rect 364195 638420 364196 638484
rect 364260 638420 364261 638484
rect 364195 638419 364261 638420
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 359043 200292 359109 200293
rect 359043 200228 359044 200292
rect 359108 200228 359109 200292
rect 359043 200227 359109 200228
rect 359046 198797 359106 200227
rect 359043 198796 359109 198797
rect 359043 198732 359044 198796
rect 359108 198732 359109 198796
rect 359043 198731 359109 198732
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 360804 182454 361404 217898
rect 364404 618054 365004 653498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 365115 639300 365181 639301
rect 365115 639236 365116 639300
rect 365180 639236 365181 639300
rect 365115 639235 365181 639236
rect 365118 638485 365178 639235
rect 365115 638484 365181 638485
rect 365115 638420 365116 638484
rect 365180 638420 365181 638484
rect 365115 638419 365181 638420
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 362907 204780 362973 204781
rect 362907 204716 362908 204780
rect 362972 204716 362973 204780
rect 362907 204715 362973 204716
rect 362910 204509 362970 204715
rect 362907 204508 362973 204509
rect 362907 204444 362908 204508
rect 362972 204444 362973 204508
rect 362907 204443 362973 204444
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 361619 180980 361685 180981
rect 361619 180916 361620 180980
rect 361684 180916 361685 180980
rect 361619 180915 361685 180916
rect 361622 180709 361682 180915
rect 361619 180708 361685 180709
rect 361619 180644 361620 180708
rect 361684 180644 361685 180708
rect 361619 180643 361685 180644
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 357387 133924 357453 133925
rect 357387 133860 357388 133924
rect 357452 133860 357453 133924
rect 357387 133859 357453 133860
rect 357390 133653 357450 133859
rect 357387 133652 357453 133653
rect 357387 133588 357388 133652
rect 357452 133588 357453 133652
rect 357387 133587 357453 133588
rect 359043 124132 359109 124133
rect 359043 124068 359044 124132
rect 359108 124068 359109 124132
rect 359043 124067 359109 124068
rect 359046 114613 359106 124067
rect 359043 114612 359109 114613
rect 359043 114548 359044 114612
rect 359108 114548 359109 114612
rect 359043 114547 359109 114548
rect 357387 110804 357453 110805
rect 357387 110740 357388 110804
rect 357452 110740 357453 110804
rect 357387 110739 357453 110740
rect 357390 110530 357450 110739
rect 357571 110532 357637 110533
rect 357571 110530 357572 110532
rect 357390 110470 357572 110530
rect 357571 110468 357572 110470
rect 357636 110468 357637 110532
rect 357571 110467 357637 110468
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 357387 76396 357453 76397
rect 357387 76332 357388 76396
rect 357452 76332 357453 76396
rect 357387 76331 357453 76332
rect 357390 76125 357450 76331
rect 357387 76124 357453 76125
rect 357387 76060 357388 76124
rect 357452 76060 357453 76124
rect 357387 76059 357453 76060
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 357387 17236 357453 17237
rect 357387 17172 357388 17236
rect 357452 17172 357453 17236
rect 357387 17171 357453 17172
rect 357390 16965 357450 17171
rect 357387 16964 357453 16965
rect 357387 16900 357388 16964
rect 357452 16900 357453 16964
rect 357387 16899 357453 16900
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 365667 123452 365733 123453
rect 365667 123388 365668 123452
rect 365732 123388 365733 123452
rect 365667 123387 365733 123388
rect 365670 123045 365730 123387
rect 365667 123044 365733 123045
rect 365667 122980 365668 123044
rect 365732 122980 365733 123044
rect 365667 122979 365733 122980
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 367139 17100 367205 17101
rect 367139 17036 367140 17100
rect 367204 17036 367205 17100
rect 367139 17035 367205 17036
rect 367142 16829 367202 17035
rect 367139 16828 367205 16829
rect 367139 16764 367140 16828
rect 367204 16764 367205 16828
rect 367139 16763 367205 16764
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 374867 639164 374933 639165
rect 374867 639100 374868 639164
rect 374932 639100 374933 639164
rect 374867 639099 374933 639100
rect 374499 639028 374565 639029
rect 374499 638964 374500 639028
rect 374564 638964 374565 639028
rect 374499 638963 374565 638964
rect 374502 638757 374562 638963
rect 374499 638756 374565 638757
rect 374499 638692 374500 638756
rect 374564 638692 374565 638756
rect 374499 638691 374565 638692
rect 374683 638756 374749 638757
rect 374683 638692 374684 638756
rect 374748 638692 374749 638756
rect 374683 638691 374749 638692
rect 374686 638485 374746 638691
rect 374870 638485 374930 639099
rect 374683 638484 374749 638485
rect 374683 638420 374684 638484
rect 374748 638420 374749 638484
rect 374683 638419 374749 638420
rect 374867 638484 374933 638485
rect 374867 638420 374868 638484
rect 374932 638420 374933 638484
rect 374867 638419 374933 638420
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 372475 204780 372541 204781
rect 372475 204716 372476 204780
rect 372540 204716 372541 204780
rect 372475 204715 372541 204716
rect 372478 204509 372538 204715
rect 372475 204508 372541 204509
rect 372475 204444 372476 204508
rect 372540 204444 372541 204508
rect 372475 204443 372541 204444
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 375419 87140 375485 87141
rect 375419 87076 375420 87140
rect 375484 87076 375485 87140
rect 375419 87075 375485 87076
rect 375422 86869 375482 87075
rect 375419 86868 375485 86869
rect 375419 86804 375420 86868
rect 375484 86804 375485 86868
rect 375419 86803 375485 86804
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 376707 76124 376773 76125
rect 376707 76060 376708 76124
rect 376772 76060 376773 76124
rect 376707 76059 376773 76060
rect 376891 76124 376957 76125
rect 376891 76060 376892 76124
rect 376956 76060 376957 76124
rect 376891 76059 376957 76060
rect 376710 75850 376770 76059
rect 376894 75850 376954 76059
rect 376710 75790 376954 75850
rect 373947 63748 374013 63749
rect 373947 63684 373948 63748
rect 374012 63684 374013 63748
rect 373947 63683 374013 63684
rect 373950 63477 374010 63683
rect 373947 63476 374013 63477
rect 373947 63412 373948 63476
rect 374012 63412 374013 63476
rect 373947 63411 374013 63412
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 373947 29612 374013 29613
rect 373947 29548 373948 29612
rect 374012 29548 374013 29612
rect 373947 29547 374013 29548
rect 373950 29341 374010 29547
rect 373947 29340 374013 29341
rect 373947 29276 373948 29340
rect 374012 29276 374013 29340
rect 373947 29275 374013 29276
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 384987 639436 385053 639437
rect 384987 639372 384988 639436
rect 385052 639372 385053 639436
rect 384987 639371 385053 639372
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 384067 639164 384133 639165
rect 384067 639100 384068 639164
rect 384132 639100 384133 639164
rect 384067 639099 384133 639100
rect 384070 638485 384130 639099
rect 384990 638893 385050 639371
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 384435 638892 384501 638893
rect 384435 638828 384436 638892
rect 384500 638890 384501 638892
rect 384803 638892 384869 638893
rect 384803 638890 384804 638892
rect 384500 638830 384804 638890
rect 384500 638828 384501 638830
rect 384435 638827 384501 638828
rect 384803 638828 384804 638830
rect 384868 638828 384869 638892
rect 384803 638827 384869 638828
rect 384987 638892 385053 638893
rect 384987 638828 384988 638892
rect 385052 638828 385053 638892
rect 384987 638827 385053 638828
rect 384251 638756 384317 638757
rect 384251 638692 384252 638756
rect 384316 638692 384317 638756
rect 384251 638691 384317 638692
rect 384254 638485 384314 638691
rect 384067 638484 384133 638485
rect 384067 638420 384068 638484
rect 384132 638420 384133 638484
rect 384067 638419 384133 638420
rect 384251 638484 384317 638485
rect 384251 638420 384252 638484
rect 384316 638420 384317 638484
rect 384251 638419 384317 638420
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 384987 157860 385053 157861
rect 384987 157796 384988 157860
rect 385052 157796 385053 157860
rect 384987 157795 385053 157796
rect 384990 157450 385050 157795
rect 384806 157390 385050 157450
rect 384806 157317 384866 157390
rect 384803 157316 384869 157317
rect 384803 157252 384804 157316
rect 384868 157252 384869 157316
rect 384803 157251 384869 157252
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 384990 87350 385234 87410
rect 384990 87277 385050 87350
rect 385174 87277 385234 87350
rect 384987 87276 385053 87277
rect 384987 87212 384988 87276
rect 385052 87212 385053 87276
rect 384987 87211 385053 87212
rect 385171 87276 385237 87277
rect 385171 87212 385172 87276
rect 385236 87212 385237 87276
rect 385171 87211 385237 87212
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 383699 40356 383765 40357
rect 383699 40292 383700 40356
rect 383764 40292 383765 40356
rect 383699 40291 383765 40292
rect 383702 40085 383762 40291
rect 383699 40084 383765 40085
rect 383699 40020 383700 40084
rect 383764 40020 383765 40084
rect 383699 40019 383765 40020
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 398603 639164 398669 639165
rect 398603 639100 398604 639164
rect 398668 639100 398669 639164
rect 398603 639099 398669 639100
rect 398971 639164 399037 639165
rect 398971 639100 398972 639164
rect 399036 639100 399037 639164
rect 398971 639099 399037 639100
rect 398606 638890 398666 639099
rect 398974 638890 399034 639099
rect 398606 638830 399034 638890
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 392163 138276 392229 138277
rect 392163 138212 392164 138276
rect 392228 138212 392229 138276
rect 392163 138211 392229 138212
rect 392166 135285 392226 138211
rect 392163 135284 392229 135285
rect 392163 135220 392164 135284
rect 392228 135220 392229 135284
rect 392163 135219 392229 135220
rect 393267 134196 393333 134197
rect 393267 134132 393268 134196
rect 393332 134132 393333 134196
rect 393267 134131 393333 134132
rect 393270 133925 393330 134131
rect 393267 133924 393333 133925
rect 393267 133860 393268 133924
rect 393332 133860 393333 133924
rect 393267 133859 393333 133860
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 618054 401004 653498
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 402835 639708 402901 639709
rect 402835 639644 402836 639708
rect 402900 639644 402901 639708
rect 402835 639643 402901 639644
rect 402838 639029 402898 639643
rect 402835 639028 402901 639029
rect 402835 638964 402836 639028
rect 402900 638964 402901 639028
rect 402835 638963 402901 638964
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 408539 639300 408605 639301
rect 408539 639236 408540 639300
rect 408604 639236 408605 639300
rect 408539 639235 408605 639236
rect 408723 639300 408789 639301
rect 408723 639236 408724 639300
rect 408788 639236 408789 639300
rect 408723 639235 408789 639236
rect 408542 639029 408602 639235
rect 408539 639028 408605 639029
rect 408539 638964 408540 639028
rect 408604 638964 408605 639028
rect 408539 638963 408605 638964
rect 408355 638892 408421 638893
rect 408355 638828 408356 638892
rect 408420 638890 408421 638892
rect 408539 638892 408605 638893
rect 408539 638890 408540 638892
rect 408420 638830 408540 638890
rect 408420 638828 408421 638830
rect 408355 638827 408421 638828
rect 408539 638828 408540 638830
rect 408604 638828 408605 638892
rect 408539 638827 408605 638828
rect 408726 638757 408786 639235
rect 408723 638756 408789 638757
rect 408723 638692 408724 638756
rect 408788 638692 408789 638756
rect 408723 638691 408789 638692
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 632454 415404 667898
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 417739 639572 417805 639573
rect 417739 639508 417740 639572
rect 417804 639508 417805 639572
rect 417739 639507 417805 639508
rect 417742 638485 417802 639507
rect 417923 638892 417989 638893
rect 417923 638828 417924 638892
rect 417988 638828 417989 638892
rect 417923 638827 417989 638828
rect 417926 638485 417986 638827
rect 417739 638484 417805 638485
rect 417739 638420 417740 638484
rect 417804 638420 417805 638484
rect 417739 638419 417805 638420
rect 417923 638484 417989 638485
rect 417923 638420 417924 638484
rect 417988 638420 417989 638484
rect 417923 638419 417989 638420
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 422707 639572 422773 639573
rect 422707 639508 422708 639572
rect 422772 639508 422773 639572
rect 422707 639507 422773 639508
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422710 638757 422770 639507
rect 422707 638756 422773 638757
rect 422707 638692 422708 638756
rect 422772 638692 422773 638756
rect 422707 638691 422773 638692
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 425099 17100 425165 17101
rect 425099 17036 425100 17100
rect 425164 17036 425165 17100
rect 425099 17035 425165 17036
rect 425102 16829 425162 17035
rect 425099 16828 425165 16829
rect 425099 16764 425100 16828
rect 425164 16764 425165 16828
rect 425099 16763 425165 16764
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 437243 639028 437309 639029
rect 437243 638964 437244 639028
rect 437308 638964 437309 639028
rect 437243 638963 437309 638964
rect 437246 638757 437306 638963
rect 437427 638892 437493 638893
rect 437427 638828 437428 638892
rect 437492 638890 437493 638892
rect 437795 638892 437861 638893
rect 437795 638890 437796 638892
rect 437492 638830 437796 638890
rect 437492 638828 437493 638830
rect 437427 638827 437493 638828
rect 437795 638828 437796 638830
rect 437860 638828 437861 638892
rect 437795 638827 437861 638828
rect 437243 638756 437309 638757
rect 437243 638692 437244 638756
rect 437308 638692 437309 638756
rect 437243 638691 437309 638692
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 456563 639028 456629 639029
rect 456563 638964 456564 639028
rect 456628 638964 456629 639028
rect 456563 638963 456629 638964
rect 456566 638757 456626 638963
rect 456563 638756 456629 638757
rect 456563 638692 456564 638756
rect 456628 638692 456629 638756
rect 456563 638691 456629 638692
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 451595 99516 451661 99517
rect 451595 99452 451596 99516
rect 451660 99452 451661 99516
rect 451595 99451 451661 99452
rect 451598 96661 451658 99451
rect 451595 96660 451661 96661
rect 451595 96596 451596 96660
rect 451660 96596 451661 96660
rect 451595 96595 451661 96596
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 453987 29612 454053 29613
rect 453987 29548 453988 29612
rect 454052 29548 454053 29612
rect 453987 29547 454053 29548
rect 453990 29205 454050 29547
rect 453987 29204 454053 29205
rect 453987 29140 453988 29204
rect 454052 29140 454053 29204
rect 453987 29139 454053 29140
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 462267 639300 462333 639301
rect 462267 639236 462268 639300
rect 462332 639236 462333 639300
rect 462267 639235 462333 639236
rect 462270 638621 462330 639235
rect 462267 638620 462333 638621
rect 462267 638556 462268 638620
rect 462332 638556 462333 638620
rect 462267 638555 462333 638556
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 463371 204780 463437 204781
rect 463371 204716 463372 204780
rect 463436 204716 463437 204780
rect 463371 204715 463437 204716
rect 463374 204370 463434 204715
rect 463555 204372 463621 204373
rect 463555 204370 463556 204372
rect 463374 204310 463556 204370
rect 463555 204308 463556 204310
rect 463620 204308 463621 204372
rect 463555 204307 463621 204308
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 463555 181116 463621 181117
rect 463555 181052 463556 181116
rect 463620 181052 463621 181116
rect 463555 181051 463621 181052
rect 463558 180845 463618 181051
rect 463555 180844 463621 180845
rect 463555 180780 463556 180844
rect 463620 180780 463621 180844
rect 463555 180779 463621 180780
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 463371 110940 463437 110941
rect 463371 110876 463372 110940
rect 463436 110876 463437 110940
rect 463371 110875 463437 110876
rect 463374 110530 463434 110875
rect 463555 110532 463621 110533
rect 463555 110530 463556 110532
rect 463374 110470 463556 110530
rect 463555 110468 463556 110470
rect 463620 110468 463621 110532
rect 463555 110467 463621 110468
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 463555 87276 463621 87277
rect 463555 87212 463556 87276
rect 463620 87212 463621 87276
rect 463555 87211 463621 87212
rect 463558 87005 463618 87211
rect 463555 87004 463621 87005
rect 463555 86940 463556 87004
rect 463620 86940 463621 87004
rect 463555 86939 463621 86940
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 463555 29476 463621 29477
rect 463555 29412 463556 29476
rect 463620 29412 463621 29476
rect 463555 29411 463621 29412
rect 463558 29069 463618 29411
rect 463555 29068 463621 29069
rect 463555 29004 463556 29068
rect 463620 29004 463621 29068
rect 463555 29003 463621 29004
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 473307 134060 473373 134061
rect 473307 133996 473308 134060
rect 473372 133996 473373 134060
rect 473307 133995 473373 133996
rect 473310 133653 473370 133995
rect 473307 133652 473373 133653
rect 473307 133588 473308 133652
rect 473372 133588 473373 133652
rect 473307 133587 473373 133588
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 488579 639300 488645 639301
rect 488579 639236 488580 639300
rect 488644 639236 488645 639300
rect 488579 639235 488645 639236
rect 488582 638485 488642 639235
rect 488579 638484 488645 638485
rect 488579 638420 488580 638484
rect 488644 638420 488645 638484
rect 488579 638419 488645 638420
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 502011 204780 502077 204781
rect 502011 204716 502012 204780
rect 502076 204716 502077 204780
rect 502011 204715 502077 204716
rect 502014 204370 502074 204715
rect 502195 204372 502261 204373
rect 502195 204370 502196 204372
rect 502014 204310 502196 204370
rect 502195 204308 502196 204310
rect 502260 204308 502261 204372
rect 502195 204307 502261 204308
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 502195 181116 502261 181117
rect 502195 181052 502196 181116
rect 502260 181052 502261 181116
rect 502195 181051 502261 181052
rect 502198 180845 502258 181051
rect 502195 180844 502261 180845
rect 502195 180780 502196 180844
rect 502260 180780 502261 180844
rect 502195 180779 502261 180780
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 502011 157860 502077 157861
rect 502011 157796 502012 157860
rect 502076 157796 502077 157860
rect 502011 157795 502077 157796
rect 502014 157450 502074 157795
rect 502195 157452 502261 157453
rect 502195 157450 502196 157452
rect 502014 157390 502196 157450
rect 502195 157388 502196 157390
rect 502260 157388 502261 157452
rect 502195 157387 502261 157388
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 502195 134196 502261 134197
rect 502195 134132 502196 134196
rect 502260 134132 502261 134196
rect 502195 134131 502261 134132
rect 502198 133925 502258 134131
rect 502195 133924 502261 133925
rect 502195 133860 502196 133924
rect 502260 133860 502261 133924
rect 502195 133859 502261 133860
rect 502011 110940 502077 110941
rect 502011 110876 502012 110940
rect 502076 110876 502077 110940
rect 502011 110875 502077 110876
rect 502014 110530 502074 110875
rect 502195 110532 502261 110533
rect 502195 110530 502196 110532
rect 502014 110470 502196 110530
rect 502195 110468 502196 110470
rect 502260 110468 502261 110532
rect 502195 110467 502261 110468
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 502195 87276 502261 87277
rect 502195 87212 502196 87276
rect 502260 87212 502261 87276
rect 502195 87211 502261 87212
rect 502198 87005 502258 87211
rect 502195 87004 502261 87005
rect 502195 86940 502196 87004
rect 502260 86940 502261 87004
rect 502195 86939 502261 86940
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 502011 64020 502077 64021
rect 502011 63956 502012 64020
rect 502076 63956 502077 64020
rect 502011 63955 502077 63956
rect 502014 63610 502074 63955
rect 502195 63612 502261 63613
rect 502195 63610 502196 63612
rect 502014 63550 502196 63610
rect 502195 63548 502196 63550
rect 502260 63548 502261 63612
rect 502195 63547 502261 63548
rect 502195 40356 502261 40357
rect 502195 40292 502196 40356
rect 502260 40292 502261 40356
rect 502195 40291 502261 40292
rect 502198 40085 502258 40291
rect 502195 40084 502261 40085
rect 502195 40020 502196 40084
rect 502260 40020 502261 40084
rect 502195 40019 502261 40020
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 502195 29476 502261 29477
rect 502195 29412 502196 29476
rect 502260 29412 502261 29476
rect 502195 29411 502261 29412
rect 502198 29069 502258 29411
rect 502195 29068 502261 29069
rect 502195 29004 502196 29068
rect 502260 29004 502261 29068
rect 502195 29003 502261 29004
rect 502011 17100 502077 17101
rect 502011 17036 502012 17100
rect 502076 17036 502077 17100
rect 502011 17035 502077 17036
rect 502014 16690 502074 17035
rect 502195 16692 502261 16693
rect 502195 16690 502196 16692
rect 502014 16630 502196 16690
rect 502195 16628 502196 16630
rect 502260 16628 502261 16692
rect 502195 16627 502261 16628
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 509739 639300 509805 639301
rect 509739 639236 509740 639300
rect 509804 639236 509805 639300
rect 509739 639235 509805 639236
rect 509742 638349 509802 639235
rect 509739 638348 509805 638349
rect 509739 638284 509740 638348
rect 509804 638284 509805 638348
rect 509739 638283 509805 638284
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 525379 639300 525445 639301
rect 525379 639236 525380 639300
rect 525444 639236 525445 639300
rect 525379 639235 525445 639236
rect 525195 638484 525261 638485
rect 525195 638420 525196 638484
rect 525260 638420 525261 638484
rect 525195 638419 525261 638420
rect 525198 638077 525258 638419
rect 525382 638213 525442 639235
rect 525563 638348 525629 638349
rect 525563 638284 525564 638348
rect 525628 638284 525629 638348
rect 525563 638283 525629 638284
rect 525379 638212 525445 638213
rect 525379 638148 525380 638212
rect 525444 638148 525445 638212
rect 525379 638147 525445 638148
rect 525195 638076 525261 638077
rect 525195 638012 525196 638076
rect 525260 638012 525261 638076
rect 525195 638011 525261 638012
rect 525566 637805 525626 638283
rect 525563 637804 525629 637805
rect 525563 637740 525564 637804
rect 525628 637740 525629 637804
rect 525563 637739 525629 637740
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 520227 87004 520293 87005
rect 520227 86940 520228 87004
rect 520292 86940 520293 87004
rect 520227 86939 520293 86940
rect 520230 86733 520290 86939
rect 520227 86732 520293 86733
rect 520227 86668 520228 86732
rect 520292 86668 520293 86732
rect 520227 86667 520293 86668
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 521515 29476 521581 29477
rect 521515 29412 521516 29476
rect 521580 29412 521581 29476
rect 521515 29411 521581 29412
rect 521518 29069 521578 29411
rect 521515 29068 521581 29069
rect 521515 29004 521516 29068
rect 521580 29004 521581 29068
rect 521515 29003 521581 29004
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 636054 527004 671498
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 527403 642836 527469 642837
rect 527403 642772 527404 642836
rect 527468 642772 527469 642836
rect 527403 642771 527469 642772
rect 527219 639300 527285 639301
rect 527219 639236 527220 639300
rect 527284 639236 527285 639300
rect 527219 639235 527285 639236
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 527222 570485 527282 639235
rect 527406 637802 527466 642771
rect 527955 642020 528021 642021
rect 527955 641956 527956 642020
rect 528020 641956 528021 642020
rect 527955 641955 528021 641956
rect 527406 637742 527650 637802
rect 527590 637533 527650 637742
rect 527587 637532 527653 637533
rect 527587 637468 527588 637532
rect 527652 637468 527653 637532
rect 527587 637467 527653 637468
rect 527403 628012 527469 628013
rect 527403 627948 527404 628012
rect 527468 627948 527469 628012
rect 527403 627947 527469 627948
rect 527406 621077 527466 627947
rect 527403 621076 527469 621077
rect 527403 621012 527404 621076
rect 527468 621012 527469 621076
rect 527403 621011 527469 621012
rect 527958 611778 528018 641955
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 529059 638484 529125 638485
rect 529059 638420 529060 638484
rect 529124 638420 529125 638484
rect 529059 638419 529125 638420
rect 528139 637396 528205 637397
rect 528139 637332 528140 637396
rect 528204 637332 528205 637396
rect 528139 637331 528205 637332
rect 528142 628149 528202 637331
rect 528139 628148 528205 628149
rect 528139 628084 528140 628148
rect 528204 628084 528205 628148
rect 528139 628083 528205 628084
rect 528323 621076 528389 621077
rect 528323 621012 528324 621076
rect 528388 621012 528389 621076
rect 528323 621011 528389 621012
rect 528326 618221 528386 621011
rect 528323 618220 528389 618221
rect 528323 618156 528324 618220
rect 528388 618156 528389 618220
rect 528323 618155 528389 618156
rect 528875 618084 528941 618085
rect 528875 618020 528876 618084
rect 528940 618020 528941 618084
rect 528875 618019 528941 618020
rect 527587 601764 527653 601765
rect 527587 601700 527588 601764
rect 527652 601700 527653 601764
rect 527587 601699 527653 601700
rect 527590 592245 527650 601699
rect 527587 592244 527653 592245
rect 527587 592180 527588 592244
rect 527652 592180 527653 592244
rect 527587 592179 527653 592180
rect 527587 591972 527653 591973
rect 527587 591908 527588 591972
rect 527652 591908 527653 591972
rect 527587 591907 527653 591908
rect 527590 589525 527650 591907
rect 527403 589524 527469 589525
rect 527403 589460 527404 589524
rect 527468 589460 527469 589524
rect 527403 589459 527469 589460
rect 527587 589524 527653 589525
rect 527587 589460 527588 589524
rect 527652 589460 527653 589524
rect 527587 589459 527653 589460
rect 527406 589250 527466 589459
rect 527406 589190 527834 589250
rect 527774 588570 527834 589190
rect 527590 588510 527834 588570
rect 527590 579730 527650 588510
rect 527590 579670 527834 579730
rect 527774 572930 527834 579670
rect 527590 572870 527834 572930
rect 527219 570484 527285 570485
rect 527219 570420 527220 570484
rect 527284 570420 527285 570484
rect 527219 570419 527285 570420
rect 527590 570213 527650 572870
rect 527587 570212 527653 570213
rect 527587 570148 527588 570212
rect 527652 570148 527653 570212
rect 527587 570147 527653 570148
rect 527219 570076 527285 570077
rect 527219 570012 527220 570076
rect 527284 570012 527285 570076
rect 527219 570011 527285 570012
rect 527403 570076 527469 570077
rect 527403 570012 527404 570076
rect 527468 570012 527469 570076
rect 527403 570011 527469 570012
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 527222 428365 527282 570011
rect 527406 568581 527466 570011
rect 527403 568580 527469 568581
rect 527403 568516 527404 568580
rect 527468 568516 527469 568580
rect 527403 568515 527469 568516
rect 527587 559060 527653 559061
rect 527587 558996 527588 559060
rect 527652 558996 527653 559060
rect 527587 558995 527653 558996
rect 527590 554029 527650 558995
rect 527587 554028 527653 554029
rect 527587 553964 527588 554028
rect 527652 553964 527653 554028
rect 527587 553963 527653 553964
rect 527958 553890 528018 610862
rect 528878 608701 528938 618019
rect 528507 608700 528573 608701
rect 528507 608636 528508 608700
rect 528572 608636 528573 608700
rect 528507 608635 528573 608636
rect 528875 608700 528941 608701
rect 528875 608636 528876 608700
rect 528940 608636 528941 608700
rect 528875 608635 528941 608636
rect 528510 601765 528570 608635
rect 528507 601764 528573 601765
rect 528507 601700 528508 601764
rect 528572 601700 528573 601764
rect 528507 601699 528573 601700
rect 528139 568580 528205 568581
rect 528139 568516 528140 568580
rect 528204 568516 528205 568580
rect 528139 568515 528205 568516
rect 528142 559197 528202 568515
rect 528139 559196 528205 559197
rect 528139 559132 528140 559196
rect 528204 559132 528205 559196
rect 528139 559131 528205 559132
rect 527590 553830 528018 553890
rect 527590 553210 527650 553830
rect 527955 553756 528021 553757
rect 527955 553692 527956 553756
rect 528020 553692 528021 553756
rect 527955 553691 528021 553692
rect 527958 553349 528018 553691
rect 527955 553348 528021 553349
rect 527955 553284 527956 553348
rect 528020 553284 528021 553348
rect 527955 553283 528021 553284
rect 527590 553150 528018 553210
rect 527587 553076 527653 553077
rect 527587 553012 527588 553076
rect 527652 553012 527653 553076
rect 527587 553011 527653 553012
rect 527590 533765 527650 553011
rect 527958 534258 528018 553150
rect 527587 533764 527653 533765
rect 527587 533700 527588 533764
rect 527652 533700 527653 533764
rect 527587 533699 527653 533700
rect 527590 514861 527650 533342
rect 527587 514860 527653 514861
rect 527587 514796 527588 514860
rect 527652 514796 527653 514860
rect 527587 514795 527653 514796
rect 527587 514724 527653 514725
rect 527587 514660 527588 514724
rect 527652 514660 527653 514724
rect 527587 514659 527653 514660
rect 527590 512277 527650 514659
rect 527587 512276 527653 512277
rect 527587 512212 527588 512276
rect 527652 512212 527653 512276
rect 527587 512211 527653 512212
rect 527771 512140 527837 512141
rect 527771 512076 527772 512140
rect 527836 512076 527837 512140
rect 527771 512075 527837 512076
rect 527774 505205 527834 512075
rect 527771 505204 527837 505205
rect 527771 505140 527772 505204
rect 527836 505140 527837 505204
rect 527771 505139 527837 505140
rect 527403 504932 527469 504933
rect 527403 504868 527404 504932
rect 527468 504868 527469 504932
rect 527403 504867 527469 504868
rect 527406 495410 527466 504867
rect 527406 495350 527834 495410
rect 527774 492557 527834 495350
rect 527771 492556 527837 492557
rect 527771 492492 527772 492556
rect 527836 492492 527837 492556
rect 527771 492491 527837 492492
rect 528139 492420 528205 492421
rect 528139 492356 528140 492420
rect 528204 492356 528205 492420
rect 528139 492355 528205 492356
rect 528142 483037 528202 492355
rect 527587 483036 527653 483037
rect 527587 482972 527588 483036
rect 527652 482972 527653 483036
rect 527587 482971 527653 482972
rect 528139 483036 528205 483037
rect 528139 482972 528140 483036
rect 528204 482972 528205 483036
rect 528139 482971 528205 482972
rect 527590 471885 527650 482971
rect 527587 471884 527653 471885
rect 527587 471820 527588 471884
rect 527652 471820 527653 471884
rect 527587 471819 527653 471820
rect 527955 471748 528021 471749
rect 527955 471684 527956 471748
rect 528020 471684 528021 471748
rect 527955 471683 528021 471684
rect 527958 462365 528018 471683
rect 527955 462364 528021 462365
rect 527955 462300 527956 462364
rect 528020 462300 528021 462364
rect 527955 462299 528021 462300
rect 528139 462364 528205 462365
rect 528139 462300 528140 462364
rect 528204 462300 528205 462364
rect 528139 462299 528205 462300
rect 528142 454069 528202 462299
rect 527771 454068 527837 454069
rect 527771 454004 527772 454068
rect 527836 454004 527837 454068
rect 527771 454003 527837 454004
rect 528139 454068 528205 454069
rect 528139 454004 528140 454068
rect 528204 454004 528205 454068
rect 528139 454003 528205 454004
rect 527774 447269 527834 454003
rect 527771 447268 527837 447269
rect 527771 447204 527772 447268
rect 527836 447204 527837 447268
rect 527771 447203 527837 447204
rect 527587 446996 527653 446997
rect 527587 446932 527588 446996
rect 527652 446932 527653 446996
rect 527587 446931 527653 446932
rect 527219 428364 527285 428365
rect 527219 428300 527220 428364
rect 527284 428300 527285 428364
rect 527219 428299 527285 428300
rect 527590 425101 527650 446931
rect 527771 428364 527837 428365
rect 527771 428300 527772 428364
rect 527836 428300 527837 428364
rect 527771 428299 527837 428300
rect 527587 425100 527653 425101
rect 527587 425036 527588 425100
rect 527652 425036 527653 425100
rect 527587 425035 527653 425036
rect 527587 424964 527653 424965
rect 527587 424900 527588 424964
rect 527652 424900 527653 424964
rect 527587 424899 527653 424900
rect 527219 421700 527285 421701
rect 527219 421636 527220 421700
rect 527284 421636 527285 421700
rect 527219 421635 527285 421636
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 527222 21997 527282 421635
rect 527590 389418 527650 424899
rect 527774 421701 527834 428299
rect 527771 421700 527837 421701
rect 527771 421636 527772 421700
rect 527836 421636 527837 421700
rect 527771 421635 527837 421636
rect 527590 368797 527650 388502
rect 527587 368796 527653 368797
rect 527587 368732 527588 368796
rect 527652 368732 527653 368796
rect 527587 368731 527653 368732
rect 529062 274685 529122 638419
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 529059 274684 529125 274685
rect 529059 274620 529060 274684
rect 529124 274620 529125 274684
rect 529059 274619 529125 274620
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 531267 204780 531333 204781
rect 531267 204716 531268 204780
rect 531332 204716 531333 204780
rect 531267 204715 531333 204716
rect 531270 204509 531330 204715
rect 531267 204508 531333 204509
rect 531267 204444 531268 204508
rect 531332 204444 531333 204508
rect 531267 204443 531333 204444
rect 531267 181252 531333 181253
rect 531267 181188 531268 181252
rect 531332 181188 531333 181252
rect 531267 181187 531333 181188
rect 531270 180981 531330 181187
rect 531267 180980 531333 180981
rect 531267 180916 531268 180980
rect 531332 180916 531333 180980
rect 531267 180915 531333 180916
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 531267 170236 531333 170237
rect 531267 170172 531268 170236
rect 531332 170172 531333 170236
rect 531267 170171 531333 170172
rect 531270 169965 531330 170171
rect 531267 169964 531333 169965
rect 531267 169900 531268 169964
rect 531332 169900 531333 169964
rect 531267 169899 531333 169900
rect 531267 157860 531333 157861
rect 531267 157796 531268 157860
rect 531332 157796 531333 157860
rect 531267 157795 531333 157796
rect 531270 157589 531330 157795
rect 531267 157588 531333 157589
rect 531267 157524 531268 157588
rect 531332 157524 531333 157588
rect 531267 157523 531333 157524
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 531267 134332 531333 134333
rect 531267 134268 531268 134332
rect 531332 134268 531333 134332
rect 531267 134267 531333 134268
rect 531270 134061 531330 134267
rect 531267 134060 531333 134061
rect 531267 133996 531268 134060
rect 531332 133996 531333 134060
rect 531267 133995 531333 133996
rect 531267 123316 531333 123317
rect 531267 123252 531268 123316
rect 531332 123252 531333 123316
rect 531267 123251 531333 123252
rect 531270 123045 531330 123251
rect 531267 123044 531333 123045
rect 531267 122980 531268 123044
rect 531332 122980 531333 123044
rect 531267 122979 531333 122980
rect 531267 110940 531333 110941
rect 531267 110876 531268 110940
rect 531332 110876 531333 110940
rect 531267 110875 531333 110876
rect 531270 110669 531330 110875
rect 531267 110668 531333 110669
rect 531267 110604 531268 110668
rect 531332 110604 531333 110668
rect 531267 110603 531333 110604
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 531267 76396 531333 76397
rect 531267 76332 531268 76396
rect 531332 76332 531333 76396
rect 531267 76331 531333 76332
rect 531270 76125 531330 76331
rect 531267 76124 531333 76125
rect 531267 76060 531268 76124
rect 531332 76060 531333 76124
rect 531267 76059 531333 76060
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 531267 64020 531333 64021
rect 531267 63956 531268 64020
rect 531332 63956 531333 64020
rect 531267 63955 531333 63956
rect 531270 63749 531330 63955
rect 531267 63748 531333 63749
rect 531267 63684 531268 63748
rect 531332 63684 531333 63748
rect 531267 63683 531333 63684
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 531267 40492 531333 40493
rect 531267 40428 531268 40492
rect 531332 40428 531333 40492
rect 531267 40427 531333 40428
rect 531270 40221 531330 40427
rect 531267 40220 531333 40221
rect 531267 40156 531268 40220
rect 531332 40156 531333 40220
rect 531267 40155 531333 40156
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 531267 29476 531333 29477
rect 531267 29412 531268 29476
rect 531332 29412 531333 29476
rect 531267 29411 531333 29412
rect 531270 29205 531330 29411
rect 531267 29204 531333 29205
rect 531267 29140 531268 29204
rect 531332 29140 531333 29204
rect 531267 29139 531333 29140
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 527219 21996 527285 21997
rect 527219 21932 527220 21996
rect 527284 21932 527285 21996
rect 527219 21931 527285 21932
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 -4946 530604 27098
rect 531267 17100 531333 17101
rect 531267 17036 531268 17100
rect 531332 17036 531333 17100
rect 531267 17035 531333 17036
rect 531270 16829 531330 17035
rect 531267 16828 531333 16829
rect 531267 16764 531268 16828
rect 531332 16764 531333 16828
rect 531267 16763 531333 16764
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 550587 204508 550653 204509
rect 550587 204444 550588 204508
rect 550652 204444 550653 204508
rect 550587 204443 550653 204444
rect 550590 204237 550650 204443
rect 550587 204236 550653 204237
rect 550587 204172 550588 204236
rect 550652 204172 550653 204236
rect 550587 204171 550653 204172
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 550587 169964 550653 169965
rect 550587 169900 550588 169964
rect 550652 169900 550653 169964
rect 550587 169899 550653 169900
rect 550590 169693 550650 169899
rect 550587 169692 550653 169693
rect 550587 169628 550588 169692
rect 550652 169628 550653 169692
rect 550587 169627 550653 169628
rect 550587 157588 550653 157589
rect 550587 157524 550588 157588
rect 550652 157524 550653 157588
rect 550587 157523 550653 157524
rect 550590 157317 550650 157523
rect 550587 157316 550653 157317
rect 550587 157252 550588 157316
rect 550652 157252 550653 157316
rect 550587 157251 550653 157252
rect 551604 157254 552204 192698
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 550587 134060 550653 134061
rect 550587 133996 550588 134060
rect 550652 133996 550653 134060
rect 550587 133995 550653 133996
rect 550590 133789 550650 133995
rect 550587 133788 550653 133789
rect 550587 133724 550588 133788
rect 550652 133724 550653 133788
rect 550587 133723 550653 133724
rect 550587 123044 550653 123045
rect 550587 122980 550588 123044
rect 550652 122980 550653 123044
rect 550587 122979 550653 122980
rect 550590 122773 550650 122979
rect 550587 122772 550653 122773
rect 550587 122708 550588 122772
rect 550652 122708 550653 122772
rect 550587 122707 550653 122708
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 550587 110668 550653 110669
rect 550587 110604 550588 110668
rect 550652 110604 550653 110668
rect 550587 110603 550653 110604
rect 550590 110397 550650 110603
rect 550587 110396 550653 110397
rect 550587 110332 550588 110396
rect 550652 110332 550653 110396
rect 550587 110331 550653 110332
rect 550587 87548 550653 87549
rect 550587 87484 550588 87548
rect 550652 87484 550653 87548
rect 550587 87483 550653 87484
rect 550590 87141 550650 87483
rect 550587 87140 550653 87141
rect 550587 87076 550588 87140
rect 550652 87076 550653 87140
rect 550587 87075 550653 87076
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 550587 76124 550653 76125
rect 550587 76060 550588 76124
rect 550652 76060 550653 76124
rect 550587 76059 550653 76060
rect 550590 75853 550650 76059
rect 550587 75852 550653 75853
rect 550587 75788 550588 75852
rect 550652 75788 550653 75852
rect 550587 75787 550653 75788
rect 550587 63748 550653 63749
rect 550587 63684 550588 63748
rect 550652 63684 550653 63748
rect 550587 63683 550653 63684
rect 550590 63477 550650 63683
rect 550587 63476 550653 63477
rect 550587 63412 550588 63476
rect 550652 63412 550653 63476
rect 550587 63411 550653 63412
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 550587 40220 550653 40221
rect 550587 40156 550588 40220
rect 550652 40156 550653 40220
rect 550587 40155 550653 40156
rect 550590 39949 550650 40155
rect 550587 39948 550653 39949
rect 550587 39884 550588 39948
rect 550652 39884 550653 39948
rect 550587 39883 550653 39884
rect 550587 29612 550653 29613
rect 550587 29548 550588 29612
rect 550652 29548 550653 29612
rect 550587 29547 550653 29548
rect 550590 29205 550650 29547
rect 550587 29204 550653 29205
rect 550587 29140 550588 29204
rect 550652 29140 550653 29204
rect 550587 29139 550653 29140
rect 550587 16828 550653 16829
rect 550587 16764 550588 16828
rect 550652 16764 550653 16828
rect 550587 16763 550653 16764
rect 550590 16557 550650 16763
rect 550587 16556 550653 16557
rect 550587 16492 550588 16556
rect 550652 16492 550653 16556
rect 550587 16491 550653 16492
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234390 529262 234626 529498
rect 235494 529262 235730 529498
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234390 520422 234626 520658
rect 233470 490502 233706 490738
rect 234390 490502 234626 490738
rect 235494 520422 235730 520658
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 233470 481662 233706 481898
rect 234390 481662 234626 481898
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234390 393942 234626 394178
rect 234390 385102 234626 385338
rect 235494 393942 235730 394178
rect 235494 385102 235730 385338
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 233470 355862 233706 356098
rect 234390 355862 234626 356098
rect 233470 346342 233706 346578
rect 234390 346342 234626 346578
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 242186 639098 242422 639334
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 527870 611542 528106 611778
rect 527870 610862 528106 611098
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 527870 534022 528106 534258
rect 527502 533342 527738 533578
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 527502 389182 527738 389418
rect 527502 388502 527738 388738
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect 526172 611778 528148 611820
rect 526172 611542 527870 611778
rect 528106 611542 528148 611778
rect 526172 611500 528148 611542
rect 526172 611140 526492 611500
rect 526172 611098 528148 611140
rect 526172 610862 527870 611098
rect 528106 610862 528148 611098
rect 526172 610820 528148 610862
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect 525988 534258 528148 534300
rect 525988 534022 527870 534258
rect 528106 534022 528148 534258
rect 525988 533980 528148 534022
rect 525988 533620 526308 533980
rect 525988 533578 527780 533620
rect 525988 533342 527502 533578
rect 527738 533342 527780 533578
rect 525988 533300 527780 533342
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect 234348 529498 235772 529540
rect 234348 529262 234390 529498
rect 234626 529262 235494 529498
rect 235730 529262 235772 529498
rect 234348 529220 235772 529262
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect 234348 520658 235772 520700
rect 234348 520422 234390 520658
rect 234626 520422 235494 520658
rect 235730 520422 235772 520658
rect 234348 520380 235772 520422
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect 233428 490738 234668 490780
rect 233428 490502 233470 490738
rect 233706 490502 234390 490738
rect 234626 490502 234668 490738
rect 233428 490460 234668 490502
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect 233428 481898 234668 481940
rect 233428 481662 233470 481898
rect 233706 481662 234390 481898
rect 234626 481662 234668 481898
rect 233428 481620 234668 481662
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect 234348 394178 235772 394220
rect 234348 393942 234390 394178
rect 234626 393942 235494 394178
rect 235730 393942 235772 394178
rect 234348 393900 235772 393942
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect 525988 389418 527780 389460
rect 525988 389182 527502 389418
rect 527738 389182 527780 389418
rect 525988 389140 527780 389182
rect 525988 388780 526308 389140
rect 525988 388738 527780 388780
rect 525988 388502 527502 388738
rect 527738 388502 527780 388738
rect 525988 388460 527780 388502
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect 234348 385338 235772 385380
rect 234348 385102 234390 385338
rect 234626 385102 235494 385338
rect 235730 385102 235772 385338
rect 234348 385060 235772 385102
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect 233428 356098 234668 356140
rect 233428 355862 233470 356098
rect 233706 355862 234390 356098
rect 234626 355862 234668 356098
rect 233428 355820 234668 355862
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect 233428 346578 234668 346620
rect 233428 346342 233470 346578
rect 233706 346342 234390 346578
rect 234626 346342 234668 346578
rect 233428 346300 234668 346342
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use user_proj_example  mprj
timestamp 1607635834
transform 1 0 230000 0 1 340000
box 0 0 299432 300000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
