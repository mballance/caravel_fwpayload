VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fwpayload
  CLASS BLOCK ;
  FOREIGN fwpayload ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 2000.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 20.440 1500.000 21.040 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1353.240 1500.000 1353.840 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1478.360 1500.000 1478.960 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1603.480 1500.000 1604.080 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1728.600 1500.000 1729.200 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1895.200 1500.000 1895.800 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1473.010 1997.600 1473.290 2000.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1258.650 1997.600 1258.930 2000.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1098.110 1997.600 1098.390 2000.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 937.110 1997.600 937.390 2000.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 776.570 1997.600 776.850 2000.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 144.880 1500.000 145.480 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 616.030 1997.600 616.310 2000.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 455.030 1997.600 455.310 2000.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 294.490 1997.600 294.770 2000.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.490 1997.600 133.770 2000.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1977.480 2.400 1978.080 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1759.880 2.400 1760.480 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1629.320 2.400 1629.920 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1498.760 2.400 1499.360 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1368.200 2.400 1368.800 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1238.320 2.400 1238.920 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 270.000 1500.000 270.600 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1107.760 2.400 1108.360 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 977.200 2.400 977.800 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 759.600 2.400 760.200 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.720 2.400 630.320 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.160 2.400 499.760 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 368.600 2.400 369.200 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 2.400 238.640 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 2.400 108.080 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 395.120 1500.000 395.720 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 520.240 1500.000 520.840 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 645.360 1500.000 645.960 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 769.800 1500.000 770.400 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 978.560 1500.000 979.160 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1103.680 1500.000 1104.280 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1228.120 1500.000 1228.720 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 103.400 1500.000 104.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1436.880 1500.000 1437.480 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1562.000 1500.000 1562.600 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1686.440 1500.000 1687.040 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1811.560 1500.000 1812.160 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1978.160 1500.000 1978.760 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1365.830 1997.600 1366.110 2000.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1151.470 1997.600 1151.750 2000.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 990.930 1997.600 991.210 2000.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 829.930 1997.600 830.210 2000.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 669.390 1997.600 669.670 2000.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 228.520 1500.000 229.120 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 508.850 1997.600 509.130 2000.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.850 1997.600 348.130 2000.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 187.310 1997.600 187.590 2000.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.770 1997.600 27.050 2000.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1890.440 2.400 1891.040 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1672.840 2.400 1673.440 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1542.280 2.400 1542.880 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1411.720 2.400 1412.320 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1281.840 2.400 1282.440 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1151.280 2.400 1151.880 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 353.640 1500.000 354.240 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1020.720 2.400 1021.320 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 890.160 2.400 890.760 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 2.400 673.840 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 2.400 543.280 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 2.400 412.720 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 281.560 2.400 282.160 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 2.400 151.600 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 2.400 21.720 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 478.080 1500.000 478.680 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 603.200 1500.000 603.800 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 728.320 1500.000 728.920 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 853.440 1500.000 854.040 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1061.520 1500.000 1062.120 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1186.640 1500.000 1187.240 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1311.760 1500.000 1312.360 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 61.920 1500.000 62.520 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1394.720 1500.000 1395.320 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1519.840 1500.000 1520.440 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1644.960 1500.000 1645.560 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1770.080 1500.000 1770.680 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1936.680 1500.000 1937.280 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1419.650 1997.600 1419.930 2000.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1205.290 1997.600 1205.570 2000.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1044.290 1997.600 1044.570 2000.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 883.750 1997.600 884.030 2000.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 723.210 1997.600 723.490 2000.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 187.040 1500.000 187.640 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 562.210 1997.600 562.490 2000.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 401.670 1997.600 401.950 2000.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 240.670 1997.600 240.950 2000.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.130 1997.600 80.410 2000.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1933.960 2.400 1934.560 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1716.360 2.400 1716.960 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1585.800 2.400 1586.400 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1455.240 2.400 1455.840 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1325.360 2.400 1325.960 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1194.800 2.400 1195.400 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 311.480 1500.000 312.080 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1064.240 2.400 1064.840 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 933.680 2.400 934.280 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.080 2.400 716.680 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 2.400 586.800 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 2.400 456.240 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 2.400 325.680 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 194.520 2.400 195.120 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 2.400 64.560 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 436.600 1500.000 437.200 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 561.720 1500.000 562.320 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 686.840 1500.000 687.440 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 811.960 1500.000 812.560 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1020.040 1500.000 1020.640 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1145.160 1500.000 1145.760 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1270.280 1500.000 1270.880 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1243.930 0.000 1244.210 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1253.130 0.000 1253.410 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1271.530 0.000 1271.810 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1280.730 0.000 1281.010 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1289.930 0.000 1290.210 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1299.130 0.000 1299.410 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1308.330 0.000 1308.610 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1317.530 0.000 1317.810 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1335.930 0.000 1336.210 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1345.130 0.000 1345.410 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1354.330 0.000 1354.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1363.530 0.000 1363.810 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1372.730 0.000 1373.010 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1381.930 0.000 1382.210 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.330 0.000 1400.610 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1409.530 0.000 1409.810 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.730 0.000 1419.010 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1427.930 0.000 1428.210 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1437.130 0.000 1437.410 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1446.330 0.000 1446.610 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1464.730 0.000 1465.010 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1473.930 0.000 1474.210 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.130 0.000 1483.410 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1492.330 0.000 1492.610 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 573.710 0.000 573.990 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 638.110 0.000 638.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 693.310 0.000 693.590 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.250 0.000 757.530 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 784.850 0.000 785.130 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 794.050 0.000 794.330 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 803.250 0.000 803.530 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 821.650 0.000 821.930 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.050 0.000 840.330 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 849.250 0.000 849.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.450 0.000 858.730 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 867.650 0.000 867.930 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.850 0.000 877.130 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 886.050 0.000 886.330 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 904.450 0.000 904.730 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 913.650 0.000 913.930 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 922.850 0.000 923.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 941.250 0.000 941.530 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 950.450 0.000 950.730 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 968.850 0.000 969.130 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 977.590 0.000 977.870 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 986.790 0.000 987.070 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 995.990 0.000 996.270 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1005.190 0.000 1005.470 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1023.590 0.000 1023.870 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.790 0.000 1033.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1041.990 0.000 1042.270 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1051.190 0.000 1051.470 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1060.390 0.000 1060.670 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1069.590 0.000 1069.870 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1087.990 0.000 1088.270 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1097.190 0.000 1097.470 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1106.390 0.000 1106.670 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1115.590 0.000 1115.870 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1124.790 0.000 1125.070 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1133.990 0.000 1134.270 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1143.190 0.000 1143.470 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1152.390 0.000 1152.670 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1161.590 0.000 1161.870 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1170.790 0.000 1171.070 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.990 0.000 1180.270 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1189.190 0.000 1189.470 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1198.390 0.000 1198.670 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1216.790 0.000 1217.070 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1225.990 0.000 1226.270 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1235.190 0.000 1235.470 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1247.150 0.000 1247.430 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1256.350 0.000 1256.630 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1274.750 0.000 1275.030 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1283.950 0.000 1284.230 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1293.150 0.000 1293.430 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1302.350 0.000 1302.630 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1311.550 0.000 1311.830 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1320.750 0.000 1321.030 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1329.950 0.000 1330.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1339.150 0.000 1339.430 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1348.350 0.000 1348.630 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1357.550 0.000 1357.830 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1366.750 0.000 1367.030 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1375.950 0.000 1376.230 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1394.350 0.000 1394.630 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1403.550 0.000 1403.830 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1412.750 0.000 1413.030 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1421.490 0.000 1421.770 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1430.690 0.000 1430.970 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1439.890 0.000 1440.170 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1458.290 0.000 1458.570 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1467.490 0.000 1467.770 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1476.690 0.000 1476.970 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1485.890 0.000 1486.170 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.090 0.000 1495.370 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.130 0.000 448.410 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 530.930 0.000 531.210 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 613.730 0.000 614.010 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 631.670 0.000 631.950 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 650.070 0.000 650.350 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 659.270 0.000 659.550 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 668.470 0.000 668.750 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 677.670 0.000 677.950 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 696.070 0.000 696.350 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 742.070 0.000 742.350 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 751.270 0.000 751.550 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 760.470 0.000 760.750 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 778.870 0.000 779.150 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 788.070 0.000 788.350 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 797.270 0.000 797.550 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 806.470 0.000 806.750 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 815.670 0.000 815.950 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 824.870 0.000 825.150 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 843.270 0.000 843.550 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.470 0.000 852.750 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 861.670 0.000 861.950 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.870 0.000 871.150 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 880.070 0.000 880.350 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 898.010 0.000 898.290 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 916.410 0.000 916.690 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 925.610 0.000 925.890 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 934.810 0.000 935.090 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 944.010 0.000 944.290 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 962.410 0.000 962.690 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 971.610 0.000 971.890 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 980.810 0.000 981.090 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 990.010 0.000 990.290 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 999.210 0.000 999.490 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1008.410 0.000 1008.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1017.610 0.000 1017.890 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1026.810 0.000 1027.090 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1036.010 0.000 1036.290 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1045.210 0.000 1045.490 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1054.410 0.000 1054.690 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1063.610 0.000 1063.890 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1072.810 0.000 1073.090 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1091.210 0.000 1091.490 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1100.410 0.000 1100.690 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1109.610 0.000 1109.890 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1118.810 0.000 1119.090 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1128.010 0.000 1128.290 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1137.210 0.000 1137.490 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1155.150 0.000 1155.430 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.550 0.000 1173.830 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1182.750 0.000 1183.030 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.950 0.000 1192.230 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1210.350 0.000 1210.630 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1219.550 0.000 1219.830 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1228.750 0.000 1229.030 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1237.950 0.000 1238.230 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1250.370 0.000 1250.650 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1259.570 0.000 1259.850 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1268.770 0.000 1269.050 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1277.970 0.000 1278.250 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.170 0.000 1287.450 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1296.370 0.000 1296.650 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1305.570 0.000 1305.850 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1314.770 0.000 1315.050 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1323.970 0.000 1324.250 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1332.710 0.000 1332.990 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1341.910 0.000 1342.190 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1351.110 0.000 1351.390 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1360.310 0.000 1360.590 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1369.510 0.000 1369.790 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1378.710 0.000 1378.990 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1397.110 0.000 1397.390 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1406.310 0.000 1406.590 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1415.510 0.000 1415.790 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1424.710 0.000 1424.990 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1433.910 0.000 1434.190 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1443.110 0.000 1443.390 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1452.310 0.000 1452.590 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1461.510 0.000 1461.790 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1470.710 0.000 1470.990 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1479.910 0.000 1480.190 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.110 0.000 1489.390 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1498.310 0.000 1498.590 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.890 0.000 681.170 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 726.890 0.000 727.170 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 736.090 0.000 736.370 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 754.490 0.000 754.770 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 791.290 0.000 791.570 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 800.030 0.000 800.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 809.230 0.000 809.510 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 818.430 0.000 818.710 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 836.830 0.000 837.110 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.030 0.000 846.310 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 855.230 0.000 855.510 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.430 0.000 864.710 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 873.630 0.000 873.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.830 0.000 883.110 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 910.430 0.000 910.710 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 919.630 0.000 919.910 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 928.830 0.000 929.110 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.030 0.000 938.310 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 947.230 0.000 947.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.630 0.000 965.910 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 974.830 0.000 975.110 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.030 0.000 984.310 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 993.230 0.000 993.510 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1002.430 0.000 1002.710 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1011.630 0.000 1011.910 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1030.030 0.000 1030.310 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1039.230 0.000 1039.510 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1048.430 0.000 1048.710 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1057.630 0.000 1057.910 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1066.370 0.000 1066.650 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1084.770 0.000 1085.050 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1093.970 0.000 1094.250 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1103.170 0.000 1103.450 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1112.370 0.000 1112.650 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1121.570 0.000 1121.850 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1130.770 0.000 1131.050 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1149.170 0.000 1149.450 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 405.350 0.000 405.630 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1158.370 0.000 1158.650 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1167.570 0.000 1167.850 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1176.770 0.000 1177.050 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.970 0.000 1186.250 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1204.370 0.000 1204.650 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1213.570 0.000 1213.850 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1222.770 0.000 1223.050 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1231.970 0.000 1232.250 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1241.170 0.000 1241.450 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 2.400 ;
    END
  END la_oen[9]
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 1853.040 1500.000 1853.640 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1846.920 2.400 1847.520 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 936.400 1500.000 937.000 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 846.640 2.400 847.240 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1312.470 1997.600 1312.750 2000.000 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1803.400 2.400 1804.000 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 1497.600 894.920 1500.000 895.520 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 803.120 2.400 803.720 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.400 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1988.560 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1988.560 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 1988.405 ;
      LAYER met1 ;
        RECT 3.290 2.760 1498.610 1989.300 ;
      LAYER met2 ;
        RECT 1.470 1997.320 26.490 1998.250 ;
        RECT 27.330 1997.320 79.850 1998.250 ;
        RECT 80.690 1997.320 133.210 1998.250 ;
        RECT 134.050 1997.320 187.030 1998.250 ;
        RECT 187.870 1997.320 240.390 1998.250 ;
        RECT 241.230 1997.320 294.210 1998.250 ;
        RECT 295.050 1997.320 347.570 1998.250 ;
        RECT 348.410 1997.320 401.390 1998.250 ;
        RECT 402.230 1997.320 454.750 1998.250 ;
        RECT 455.590 1997.320 508.570 1998.250 ;
        RECT 509.410 1997.320 561.930 1998.250 ;
        RECT 562.770 1997.320 615.750 1998.250 ;
        RECT 616.590 1997.320 669.110 1998.250 ;
        RECT 669.950 1997.320 722.930 1998.250 ;
        RECT 723.770 1997.320 776.290 1998.250 ;
        RECT 777.130 1997.320 829.650 1998.250 ;
        RECT 830.490 1997.320 883.470 1998.250 ;
        RECT 884.310 1997.320 936.830 1998.250 ;
        RECT 937.670 1997.320 990.650 1998.250 ;
        RECT 991.490 1997.320 1044.010 1998.250 ;
        RECT 1044.850 1997.320 1097.830 1998.250 ;
        RECT 1098.670 1997.320 1151.190 1998.250 ;
        RECT 1152.030 1997.320 1205.010 1998.250 ;
        RECT 1205.850 1997.320 1258.370 1998.250 ;
        RECT 1259.210 1997.320 1312.190 1998.250 ;
        RECT 1313.030 1997.320 1365.550 1998.250 ;
        RECT 1366.390 1997.320 1419.370 1998.250 ;
        RECT 1420.210 1997.320 1472.730 1998.250 ;
        RECT 1473.570 1997.320 1498.580 1998.250 ;
        RECT 1.470 2.680 1498.580 1997.320 ;
        RECT 2.030 2.400 3.950 2.680 ;
        RECT 4.790 2.400 7.170 2.680 ;
        RECT 8.010 2.400 9.930 2.680 ;
        RECT 10.770 2.400 13.150 2.680 ;
        RECT 13.990 2.400 16.370 2.680 ;
        RECT 17.210 2.400 19.130 2.680 ;
        RECT 19.970 2.400 22.350 2.680 ;
        RECT 23.190 2.400 25.570 2.680 ;
        RECT 26.410 2.400 28.330 2.680 ;
        RECT 29.170 2.400 31.550 2.680 ;
        RECT 32.390 2.400 34.770 2.680 ;
        RECT 35.610 2.400 37.530 2.680 ;
        RECT 38.370 2.400 40.750 2.680 ;
        RECT 41.590 2.400 43.970 2.680 ;
        RECT 44.810 2.400 46.730 2.680 ;
        RECT 47.570 2.400 49.950 2.680 ;
        RECT 50.790 2.400 53.170 2.680 ;
        RECT 54.010 2.400 55.930 2.680 ;
        RECT 56.770 2.400 59.150 2.680 ;
        RECT 59.990 2.400 62.370 2.680 ;
        RECT 63.210 2.400 65.130 2.680 ;
        RECT 65.970 2.400 68.350 2.680 ;
        RECT 69.190 2.400 71.570 2.680 ;
        RECT 72.410 2.400 74.330 2.680 ;
        RECT 75.170 2.400 77.550 2.680 ;
        RECT 78.390 2.400 80.770 2.680 ;
        RECT 81.610 2.400 83.530 2.680 ;
        RECT 84.370 2.400 86.750 2.680 ;
        RECT 87.590 2.400 89.510 2.680 ;
        RECT 90.350 2.400 92.730 2.680 ;
        RECT 93.570 2.400 95.950 2.680 ;
        RECT 96.790 2.400 98.710 2.680 ;
        RECT 99.550 2.400 101.930 2.680 ;
        RECT 102.770 2.400 105.150 2.680 ;
        RECT 105.990 2.400 107.910 2.680 ;
        RECT 108.750 2.400 111.130 2.680 ;
        RECT 111.970 2.400 114.350 2.680 ;
        RECT 115.190 2.400 117.110 2.680 ;
        RECT 117.950 2.400 120.330 2.680 ;
        RECT 121.170 2.400 123.550 2.680 ;
        RECT 124.390 2.400 126.310 2.680 ;
        RECT 127.150 2.400 129.530 2.680 ;
        RECT 130.370 2.400 132.750 2.680 ;
        RECT 133.590 2.400 135.510 2.680 ;
        RECT 136.350 2.400 138.730 2.680 ;
        RECT 139.570 2.400 141.950 2.680 ;
        RECT 142.790 2.400 144.710 2.680 ;
        RECT 145.550 2.400 147.930 2.680 ;
        RECT 148.770 2.400 151.150 2.680 ;
        RECT 151.990 2.400 153.910 2.680 ;
        RECT 154.750 2.400 157.130 2.680 ;
        RECT 157.970 2.400 160.350 2.680 ;
        RECT 161.190 2.400 163.110 2.680 ;
        RECT 163.950 2.400 166.330 2.680 ;
        RECT 167.170 2.400 169.550 2.680 ;
        RECT 170.390 2.400 172.310 2.680 ;
        RECT 173.150 2.400 175.530 2.680 ;
        RECT 176.370 2.400 178.290 2.680 ;
        RECT 179.130 2.400 181.510 2.680 ;
        RECT 182.350 2.400 184.730 2.680 ;
        RECT 185.570 2.400 187.490 2.680 ;
        RECT 188.330 2.400 190.710 2.680 ;
        RECT 191.550 2.400 193.930 2.680 ;
        RECT 194.770 2.400 196.690 2.680 ;
        RECT 197.530 2.400 199.910 2.680 ;
        RECT 200.750 2.400 203.130 2.680 ;
        RECT 203.970 2.400 205.890 2.680 ;
        RECT 206.730 2.400 209.110 2.680 ;
        RECT 209.950 2.400 212.330 2.680 ;
        RECT 213.170 2.400 215.090 2.680 ;
        RECT 215.930 2.400 218.310 2.680 ;
        RECT 219.150 2.400 221.530 2.680 ;
        RECT 222.370 2.400 224.290 2.680 ;
        RECT 225.130 2.400 227.510 2.680 ;
        RECT 228.350 2.400 230.730 2.680 ;
        RECT 231.570 2.400 233.490 2.680 ;
        RECT 234.330 2.400 236.710 2.680 ;
        RECT 237.550 2.400 239.930 2.680 ;
        RECT 240.770 2.400 242.690 2.680 ;
        RECT 243.530 2.400 245.910 2.680 ;
        RECT 246.750 2.400 249.130 2.680 ;
        RECT 249.970 2.400 251.890 2.680 ;
        RECT 252.730 2.400 255.110 2.680 ;
        RECT 255.950 2.400 258.330 2.680 ;
        RECT 259.170 2.400 261.090 2.680 ;
        RECT 261.930 2.400 264.310 2.680 ;
        RECT 265.150 2.400 267.070 2.680 ;
        RECT 267.910 2.400 270.290 2.680 ;
        RECT 271.130 2.400 273.510 2.680 ;
        RECT 274.350 2.400 276.270 2.680 ;
        RECT 277.110 2.400 279.490 2.680 ;
        RECT 280.330 2.400 282.710 2.680 ;
        RECT 283.550 2.400 285.470 2.680 ;
        RECT 286.310 2.400 288.690 2.680 ;
        RECT 289.530 2.400 291.910 2.680 ;
        RECT 292.750 2.400 294.670 2.680 ;
        RECT 295.510 2.400 297.890 2.680 ;
        RECT 298.730 2.400 301.110 2.680 ;
        RECT 301.950 2.400 303.870 2.680 ;
        RECT 304.710 2.400 307.090 2.680 ;
        RECT 307.930 2.400 310.310 2.680 ;
        RECT 311.150 2.400 313.070 2.680 ;
        RECT 313.910 2.400 316.290 2.680 ;
        RECT 317.130 2.400 319.510 2.680 ;
        RECT 320.350 2.400 322.270 2.680 ;
        RECT 323.110 2.400 325.490 2.680 ;
        RECT 326.330 2.400 328.710 2.680 ;
        RECT 329.550 2.400 331.470 2.680 ;
        RECT 332.310 2.400 334.690 2.680 ;
        RECT 335.530 2.400 337.910 2.680 ;
        RECT 338.750 2.400 340.670 2.680 ;
        RECT 341.510 2.400 343.890 2.680 ;
        RECT 344.730 2.400 347.110 2.680 ;
        RECT 347.950 2.400 349.870 2.680 ;
        RECT 350.710 2.400 353.090 2.680 ;
        RECT 353.930 2.400 355.850 2.680 ;
        RECT 356.690 2.400 359.070 2.680 ;
        RECT 359.910 2.400 362.290 2.680 ;
        RECT 363.130 2.400 365.050 2.680 ;
        RECT 365.890 2.400 368.270 2.680 ;
        RECT 369.110 2.400 371.490 2.680 ;
        RECT 372.330 2.400 374.250 2.680 ;
        RECT 375.090 2.400 377.470 2.680 ;
        RECT 378.310 2.400 380.690 2.680 ;
        RECT 381.530 2.400 383.450 2.680 ;
        RECT 384.290 2.400 386.670 2.680 ;
        RECT 387.510 2.400 389.890 2.680 ;
        RECT 390.730 2.400 392.650 2.680 ;
        RECT 393.490 2.400 395.870 2.680 ;
        RECT 396.710 2.400 399.090 2.680 ;
        RECT 399.930 2.400 401.850 2.680 ;
        RECT 402.690 2.400 405.070 2.680 ;
        RECT 405.910 2.400 408.290 2.680 ;
        RECT 409.130 2.400 411.050 2.680 ;
        RECT 411.890 2.400 414.270 2.680 ;
        RECT 415.110 2.400 417.490 2.680 ;
        RECT 418.330 2.400 420.250 2.680 ;
        RECT 421.090 2.400 423.470 2.680 ;
        RECT 424.310 2.400 426.690 2.680 ;
        RECT 427.530 2.400 429.450 2.680 ;
        RECT 430.290 2.400 432.670 2.680 ;
        RECT 433.510 2.400 435.890 2.680 ;
        RECT 436.730 2.400 438.650 2.680 ;
        RECT 439.490 2.400 441.870 2.680 ;
        RECT 442.710 2.400 444.630 2.680 ;
        RECT 445.470 2.400 447.850 2.680 ;
        RECT 448.690 2.400 451.070 2.680 ;
        RECT 451.910 2.400 453.830 2.680 ;
        RECT 454.670 2.400 457.050 2.680 ;
        RECT 457.890 2.400 460.270 2.680 ;
        RECT 461.110 2.400 463.030 2.680 ;
        RECT 463.870 2.400 466.250 2.680 ;
        RECT 467.090 2.400 469.470 2.680 ;
        RECT 470.310 2.400 472.230 2.680 ;
        RECT 473.070 2.400 475.450 2.680 ;
        RECT 476.290 2.400 478.670 2.680 ;
        RECT 479.510 2.400 481.430 2.680 ;
        RECT 482.270 2.400 484.650 2.680 ;
        RECT 485.490 2.400 487.870 2.680 ;
        RECT 488.710 2.400 490.630 2.680 ;
        RECT 491.470 2.400 493.850 2.680 ;
        RECT 494.690 2.400 497.070 2.680 ;
        RECT 497.910 2.400 499.830 2.680 ;
        RECT 500.670 2.400 503.050 2.680 ;
        RECT 503.890 2.400 506.270 2.680 ;
        RECT 507.110 2.400 509.030 2.680 ;
        RECT 509.870 2.400 512.250 2.680 ;
        RECT 513.090 2.400 515.470 2.680 ;
        RECT 516.310 2.400 518.230 2.680 ;
        RECT 519.070 2.400 521.450 2.680 ;
        RECT 522.290 2.400 524.670 2.680 ;
        RECT 525.510 2.400 527.430 2.680 ;
        RECT 528.270 2.400 530.650 2.680 ;
        RECT 531.490 2.400 533.410 2.680 ;
        RECT 534.250 2.400 536.630 2.680 ;
        RECT 537.470 2.400 539.850 2.680 ;
        RECT 540.690 2.400 542.610 2.680 ;
        RECT 543.450 2.400 545.830 2.680 ;
        RECT 546.670 2.400 549.050 2.680 ;
        RECT 549.890 2.400 551.810 2.680 ;
        RECT 552.650 2.400 555.030 2.680 ;
        RECT 555.870 2.400 558.250 2.680 ;
        RECT 559.090 2.400 561.010 2.680 ;
        RECT 561.850 2.400 564.230 2.680 ;
        RECT 565.070 2.400 567.450 2.680 ;
        RECT 568.290 2.400 570.210 2.680 ;
        RECT 571.050 2.400 573.430 2.680 ;
        RECT 574.270 2.400 576.650 2.680 ;
        RECT 577.490 2.400 579.410 2.680 ;
        RECT 580.250 2.400 582.630 2.680 ;
        RECT 583.470 2.400 585.850 2.680 ;
        RECT 586.690 2.400 588.610 2.680 ;
        RECT 589.450 2.400 591.830 2.680 ;
        RECT 592.670 2.400 595.050 2.680 ;
        RECT 595.890 2.400 597.810 2.680 ;
        RECT 598.650 2.400 601.030 2.680 ;
        RECT 601.870 2.400 604.250 2.680 ;
        RECT 605.090 2.400 607.010 2.680 ;
        RECT 607.850 2.400 610.230 2.680 ;
        RECT 611.070 2.400 613.450 2.680 ;
        RECT 614.290 2.400 616.210 2.680 ;
        RECT 617.050 2.400 619.430 2.680 ;
        RECT 620.270 2.400 622.190 2.680 ;
        RECT 623.030 2.400 625.410 2.680 ;
        RECT 626.250 2.400 628.630 2.680 ;
        RECT 629.470 2.400 631.390 2.680 ;
        RECT 632.230 2.400 634.610 2.680 ;
        RECT 635.450 2.400 637.830 2.680 ;
        RECT 638.670 2.400 640.590 2.680 ;
        RECT 641.430 2.400 643.810 2.680 ;
        RECT 644.650 2.400 647.030 2.680 ;
        RECT 647.870 2.400 649.790 2.680 ;
        RECT 650.630 2.400 653.010 2.680 ;
        RECT 653.850 2.400 656.230 2.680 ;
        RECT 657.070 2.400 658.990 2.680 ;
        RECT 659.830 2.400 662.210 2.680 ;
        RECT 663.050 2.400 665.430 2.680 ;
        RECT 666.270 2.400 668.190 2.680 ;
        RECT 669.030 2.400 671.410 2.680 ;
        RECT 672.250 2.400 674.630 2.680 ;
        RECT 675.470 2.400 677.390 2.680 ;
        RECT 678.230 2.400 680.610 2.680 ;
        RECT 681.450 2.400 683.830 2.680 ;
        RECT 684.670 2.400 686.590 2.680 ;
        RECT 687.430 2.400 689.810 2.680 ;
        RECT 690.650 2.400 693.030 2.680 ;
        RECT 693.870 2.400 695.790 2.680 ;
        RECT 696.630 2.400 699.010 2.680 ;
        RECT 699.850 2.400 702.230 2.680 ;
        RECT 703.070 2.400 704.990 2.680 ;
        RECT 705.830 2.400 708.210 2.680 ;
        RECT 709.050 2.400 710.970 2.680 ;
        RECT 711.810 2.400 714.190 2.680 ;
        RECT 715.030 2.400 717.410 2.680 ;
        RECT 718.250 2.400 720.170 2.680 ;
        RECT 721.010 2.400 723.390 2.680 ;
        RECT 724.230 2.400 726.610 2.680 ;
        RECT 727.450 2.400 729.370 2.680 ;
        RECT 730.210 2.400 732.590 2.680 ;
        RECT 733.430 2.400 735.810 2.680 ;
        RECT 736.650 2.400 738.570 2.680 ;
        RECT 739.410 2.400 741.790 2.680 ;
        RECT 742.630 2.400 745.010 2.680 ;
        RECT 745.850 2.400 747.770 2.680 ;
        RECT 748.610 2.400 750.990 2.680 ;
        RECT 751.830 2.400 754.210 2.680 ;
        RECT 755.050 2.400 756.970 2.680 ;
        RECT 757.810 2.400 760.190 2.680 ;
        RECT 761.030 2.400 763.410 2.680 ;
        RECT 764.250 2.400 766.170 2.680 ;
        RECT 767.010 2.400 769.390 2.680 ;
        RECT 770.230 2.400 772.610 2.680 ;
        RECT 773.450 2.400 775.370 2.680 ;
        RECT 776.210 2.400 778.590 2.680 ;
        RECT 779.430 2.400 781.810 2.680 ;
        RECT 782.650 2.400 784.570 2.680 ;
        RECT 785.410 2.400 787.790 2.680 ;
        RECT 788.630 2.400 791.010 2.680 ;
        RECT 791.850 2.400 793.770 2.680 ;
        RECT 794.610 2.400 796.990 2.680 ;
        RECT 797.830 2.400 799.750 2.680 ;
        RECT 800.590 2.400 802.970 2.680 ;
        RECT 803.810 2.400 806.190 2.680 ;
        RECT 807.030 2.400 808.950 2.680 ;
        RECT 809.790 2.400 812.170 2.680 ;
        RECT 813.010 2.400 815.390 2.680 ;
        RECT 816.230 2.400 818.150 2.680 ;
        RECT 818.990 2.400 821.370 2.680 ;
        RECT 822.210 2.400 824.590 2.680 ;
        RECT 825.430 2.400 827.350 2.680 ;
        RECT 828.190 2.400 830.570 2.680 ;
        RECT 831.410 2.400 833.790 2.680 ;
        RECT 834.630 2.400 836.550 2.680 ;
        RECT 837.390 2.400 839.770 2.680 ;
        RECT 840.610 2.400 842.990 2.680 ;
        RECT 843.830 2.400 845.750 2.680 ;
        RECT 846.590 2.400 848.970 2.680 ;
        RECT 849.810 2.400 852.190 2.680 ;
        RECT 853.030 2.400 854.950 2.680 ;
        RECT 855.790 2.400 858.170 2.680 ;
        RECT 859.010 2.400 861.390 2.680 ;
        RECT 862.230 2.400 864.150 2.680 ;
        RECT 864.990 2.400 867.370 2.680 ;
        RECT 868.210 2.400 870.590 2.680 ;
        RECT 871.430 2.400 873.350 2.680 ;
        RECT 874.190 2.400 876.570 2.680 ;
        RECT 877.410 2.400 879.790 2.680 ;
        RECT 880.630 2.400 882.550 2.680 ;
        RECT 883.390 2.400 885.770 2.680 ;
        RECT 886.610 2.400 888.530 2.680 ;
        RECT 889.370 2.400 891.750 2.680 ;
        RECT 892.590 2.400 894.970 2.680 ;
        RECT 895.810 2.400 897.730 2.680 ;
        RECT 898.570 2.400 900.950 2.680 ;
        RECT 901.790 2.400 904.170 2.680 ;
        RECT 905.010 2.400 906.930 2.680 ;
        RECT 907.770 2.400 910.150 2.680 ;
        RECT 910.990 2.400 913.370 2.680 ;
        RECT 914.210 2.400 916.130 2.680 ;
        RECT 916.970 2.400 919.350 2.680 ;
        RECT 920.190 2.400 922.570 2.680 ;
        RECT 923.410 2.400 925.330 2.680 ;
        RECT 926.170 2.400 928.550 2.680 ;
        RECT 929.390 2.400 931.770 2.680 ;
        RECT 932.610 2.400 934.530 2.680 ;
        RECT 935.370 2.400 937.750 2.680 ;
        RECT 938.590 2.400 940.970 2.680 ;
        RECT 941.810 2.400 943.730 2.680 ;
        RECT 944.570 2.400 946.950 2.680 ;
        RECT 947.790 2.400 950.170 2.680 ;
        RECT 951.010 2.400 952.930 2.680 ;
        RECT 953.770 2.400 956.150 2.680 ;
        RECT 956.990 2.400 959.370 2.680 ;
        RECT 960.210 2.400 962.130 2.680 ;
        RECT 962.970 2.400 965.350 2.680 ;
        RECT 966.190 2.400 968.570 2.680 ;
        RECT 969.410 2.400 971.330 2.680 ;
        RECT 972.170 2.400 974.550 2.680 ;
        RECT 975.390 2.400 977.310 2.680 ;
        RECT 978.150 2.400 980.530 2.680 ;
        RECT 981.370 2.400 983.750 2.680 ;
        RECT 984.590 2.400 986.510 2.680 ;
        RECT 987.350 2.400 989.730 2.680 ;
        RECT 990.570 2.400 992.950 2.680 ;
        RECT 993.790 2.400 995.710 2.680 ;
        RECT 996.550 2.400 998.930 2.680 ;
        RECT 999.770 2.400 1002.150 2.680 ;
        RECT 1002.990 2.400 1004.910 2.680 ;
        RECT 1005.750 2.400 1008.130 2.680 ;
        RECT 1008.970 2.400 1011.350 2.680 ;
        RECT 1012.190 2.400 1014.110 2.680 ;
        RECT 1014.950 2.400 1017.330 2.680 ;
        RECT 1018.170 2.400 1020.550 2.680 ;
        RECT 1021.390 2.400 1023.310 2.680 ;
        RECT 1024.150 2.400 1026.530 2.680 ;
        RECT 1027.370 2.400 1029.750 2.680 ;
        RECT 1030.590 2.400 1032.510 2.680 ;
        RECT 1033.350 2.400 1035.730 2.680 ;
        RECT 1036.570 2.400 1038.950 2.680 ;
        RECT 1039.790 2.400 1041.710 2.680 ;
        RECT 1042.550 2.400 1044.930 2.680 ;
        RECT 1045.770 2.400 1048.150 2.680 ;
        RECT 1048.990 2.400 1050.910 2.680 ;
        RECT 1051.750 2.400 1054.130 2.680 ;
        RECT 1054.970 2.400 1057.350 2.680 ;
        RECT 1058.190 2.400 1060.110 2.680 ;
        RECT 1060.950 2.400 1063.330 2.680 ;
        RECT 1064.170 2.400 1066.090 2.680 ;
        RECT 1066.930 2.400 1069.310 2.680 ;
        RECT 1070.150 2.400 1072.530 2.680 ;
        RECT 1073.370 2.400 1075.290 2.680 ;
        RECT 1076.130 2.400 1078.510 2.680 ;
        RECT 1079.350 2.400 1081.730 2.680 ;
        RECT 1082.570 2.400 1084.490 2.680 ;
        RECT 1085.330 2.400 1087.710 2.680 ;
        RECT 1088.550 2.400 1090.930 2.680 ;
        RECT 1091.770 2.400 1093.690 2.680 ;
        RECT 1094.530 2.400 1096.910 2.680 ;
        RECT 1097.750 2.400 1100.130 2.680 ;
        RECT 1100.970 2.400 1102.890 2.680 ;
        RECT 1103.730 2.400 1106.110 2.680 ;
        RECT 1106.950 2.400 1109.330 2.680 ;
        RECT 1110.170 2.400 1112.090 2.680 ;
        RECT 1112.930 2.400 1115.310 2.680 ;
        RECT 1116.150 2.400 1118.530 2.680 ;
        RECT 1119.370 2.400 1121.290 2.680 ;
        RECT 1122.130 2.400 1124.510 2.680 ;
        RECT 1125.350 2.400 1127.730 2.680 ;
        RECT 1128.570 2.400 1130.490 2.680 ;
        RECT 1131.330 2.400 1133.710 2.680 ;
        RECT 1134.550 2.400 1136.930 2.680 ;
        RECT 1137.770 2.400 1139.690 2.680 ;
        RECT 1140.530 2.400 1142.910 2.680 ;
        RECT 1143.750 2.400 1146.130 2.680 ;
        RECT 1146.970 2.400 1148.890 2.680 ;
        RECT 1149.730 2.400 1152.110 2.680 ;
        RECT 1152.950 2.400 1154.870 2.680 ;
        RECT 1155.710 2.400 1158.090 2.680 ;
        RECT 1158.930 2.400 1161.310 2.680 ;
        RECT 1162.150 2.400 1164.070 2.680 ;
        RECT 1164.910 2.400 1167.290 2.680 ;
        RECT 1168.130 2.400 1170.510 2.680 ;
        RECT 1171.350 2.400 1173.270 2.680 ;
        RECT 1174.110 2.400 1176.490 2.680 ;
        RECT 1177.330 2.400 1179.710 2.680 ;
        RECT 1180.550 2.400 1182.470 2.680 ;
        RECT 1183.310 2.400 1185.690 2.680 ;
        RECT 1186.530 2.400 1188.910 2.680 ;
        RECT 1189.750 2.400 1191.670 2.680 ;
        RECT 1192.510 2.400 1194.890 2.680 ;
        RECT 1195.730 2.400 1198.110 2.680 ;
        RECT 1198.950 2.400 1200.870 2.680 ;
        RECT 1201.710 2.400 1204.090 2.680 ;
        RECT 1204.930 2.400 1207.310 2.680 ;
        RECT 1208.150 2.400 1210.070 2.680 ;
        RECT 1210.910 2.400 1213.290 2.680 ;
        RECT 1214.130 2.400 1216.510 2.680 ;
        RECT 1217.350 2.400 1219.270 2.680 ;
        RECT 1220.110 2.400 1222.490 2.680 ;
        RECT 1223.330 2.400 1225.710 2.680 ;
        RECT 1226.550 2.400 1228.470 2.680 ;
        RECT 1229.310 2.400 1231.690 2.680 ;
        RECT 1232.530 2.400 1234.910 2.680 ;
        RECT 1235.750 2.400 1237.670 2.680 ;
        RECT 1238.510 2.400 1240.890 2.680 ;
        RECT 1241.730 2.400 1243.650 2.680 ;
        RECT 1244.490 2.400 1246.870 2.680 ;
        RECT 1247.710 2.400 1250.090 2.680 ;
        RECT 1250.930 2.400 1252.850 2.680 ;
        RECT 1253.690 2.400 1256.070 2.680 ;
        RECT 1256.910 2.400 1259.290 2.680 ;
        RECT 1260.130 2.400 1262.050 2.680 ;
        RECT 1262.890 2.400 1265.270 2.680 ;
        RECT 1266.110 2.400 1268.490 2.680 ;
        RECT 1269.330 2.400 1271.250 2.680 ;
        RECT 1272.090 2.400 1274.470 2.680 ;
        RECT 1275.310 2.400 1277.690 2.680 ;
        RECT 1278.530 2.400 1280.450 2.680 ;
        RECT 1281.290 2.400 1283.670 2.680 ;
        RECT 1284.510 2.400 1286.890 2.680 ;
        RECT 1287.730 2.400 1289.650 2.680 ;
        RECT 1290.490 2.400 1292.870 2.680 ;
        RECT 1293.710 2.400 1296.090 2.680 ;
        RECT 1296.930 2.400 1298.850 2.680 ;
        RECT 1299.690 2.400 1302.070 2.680 ;
        RECT 1302.910 2.400 1305.290 2.680 ;
        RECT 1306.130 2.400 1308.050 2.680 ;
        RECT 1308.890 2.400 1311.270 2.680 ;
        RECT 1312.110 2.400 1314.490 2.680 ;
        RECT 1315.330 2.400 1317.250 2.680 ;
        RECT 1318.090 2.400 1320.470 2.680 ;
        RECT 1321.310 2.400 1323.690 2.680 ;
        RECT 1324.530 2.400 1326.450 2.680 ;
        RECT 1327.290 2.400 1329.670 2.680 ;
        RECT 1330.510 2.400 1332.430 2.680 ;
        RECT 1333.270 2.400 1335.650 2.680 ;
        RECT 1336.490 2.400 1338.870 2.680 ;
        RECT 1339.710 2.400 1341.630 2.680 ;
        RECT 1342.470 2.400 1344.850 2.680 ;
        RECT 1345.690 2.400 1348.070 2.680 ;
        RECT 1348.910 2.400 1350.830 2.680 ;
        RECT 1351.670 2.400 1354.050 2.680 ;
        RECT 1354.890 2.400 1357.270 2.680 ;
        RECT 1358.110 2.400 1360.030 2.680 ;
        RECT 1360.870 2.400 1363.250 2.680 ;
        RECT 1364.090 2.400 1366.470 2.680 ;
        RECT 1367.310 2.400 1369.230 2.680 ;
        RECT 1370.070 2.400 1372.450 2.680 ;
        RECT 1373.290 2.400 1375.670 2.680 ;
        RECT 1376.510 2.400 1378.430 2.680 ;
        RECT 1379.270 2.400 1381.650 2.680 ;
        RECT 1382.490 2.400 1384.870 2.680 ;
        RECT 1385.710 2.400 1387.630 2.680 ;
        RECT 1388.470 2.400 1390.850 2.680 ;
        RECT 1391.690 2.400 1394.070 2.680 ;
        RECT 1394.910 2.400 1396.830 2.680 ;
        RECT 1397.670 2.400 1400.050 2.680 ;
        RECT 1400.890 2.400 1403.270 2.680 ;
        RECT 1404.110 2.400 1406.030 2.680 ;
        RECT 1406.870 2.400 1409.250 2.680 ;
        RECT 1410.090 2.400 1412.470 2.680 ;
        RECT 1413.310 2.400 1415.230 2.680 ;
        RECT 1416.070 2.400 1418.450 2.680 ;
        RECT 1419.290 2.400 1421.210 2.680 ;
        RECT 1422.050 2.400 1424.430 2.680 ;
        RECT 1425.270 2.400 1427.650 2.680 ;
        RECT 1428.490 2.400 1430.410 2.680 ;
        RECT 1431.250 2.400 1433.630 2.680 ;
        RECT 1434.470 2.400 1436.850 2.680 ;
        RECT 1437.690 2.400 1439.610 2.680 ;
        RECT 1440.450 2.400 1442.830 2.680 ;
        RECT 1443.670 2.400 1446.050 2.680 ;
        RECT 1446.890 2.400 1448.810 2.680 ;
        RECT 1449.650 2.400 1452.030 2.680 ;
        RECT 1452.870 2.400 1455.250 2.680 ;
        RECT 1456.090 2.400 1458.010 2.680 ;
        RECT 1458.850 2.400 1461.230 2.680 ;
        RECT 1462.070 2.400 1464.450 2.680 ;
        RECT 1465.290 2.400 1467.210 2.680 ;
        RECT 1468.050 2.400 1470.430 2.680 ;
        RECT 1471.270 2.400 1473.650 2.680 ;
        RECT 1474.490 2.400 1476.410 2.680 ;
        RECT 1477.250 2.400 1479.630 2.680 ;
        RECT 1480.470 2.400 1482.850 2.680 ;
        RECT 1483.690 2.400 1485.610 2.680 ;
        RECT 1486.450 2.400 1488.830 2.680 ;
        RECT 1489.670 2.400 1492.050 2.680 ;
        RECT 1492.890 2.400 1494.810 2.680 ;
        RECT 1495.650 2.400 1498.030 2.680 ;
      LAYER met3 ;
        RECT 1.445 1979.160 1497.600 1988.485 ;
        RECT 1.445 1978.480 1497.200 1979.160 ;
        RECT 2.800 1977.760 1497.200 1978.480 ;
        RECT 2.800 1977.080 1497.600 1977.760 ;
        RECT 1.445 1937.680 1497.600 1977.080 ;
        RECT 1.445 1936.280 1497.200 1937.680 ;
        RECT 1.445 1934.960 1497.600 1936.280 ;
        RECT 2.800 1933.560 1497.600 1934.960 ;
        RECT 1.445 1896.200 1497.600 1933.560 ;
        RECT 1.445 1894.800 1497.200 1896.200 ;
        RECT 1.445 1891.440 1497.600 1894.800 ;
        RECT 2.800 1890.040 1497.600 1891.440 ;
        RECT 1.445 1854.040 1497.600 1890.040 ;
        RECT 1.445 1852.640 1497.200 1854.040 ;
        RECT 1.445 1847.920 1497.600 1852.640 ;
        RECT 2.800 1846.520 1497.600 1847.920 ;
        RECT 1.445 1812.560 1497.600 1846.520 ;
        RECT 1.445 1811.160 1497.200 1812.560 ;
        RECT 1.445 1804.400 1497.600 1811.160 ;
        RECT 2.800 1803.000 1497.600 1804.400 ;
        RECT 1.445 1771.080 1497.600 1803.000 ;
        RECT 1.445 1769.680 1497.200 1771.080 ;
        RECT 1.445 1760.880 1497.600 1769.680 ;
        RECT 2.800 1759.480 1497.600 1760.880 ;
        RECT 1.445 1729.600 1497.600 1759.480 ;
        RECT 1.445 1728.200 1497.200 1729.600 ;
        RECT 1.445 1717.360 1497.600 1728.200 ;
        RECT 2.800 1715.960 1497.600 1717.360 ;
        RECT 1.445 1687.440 1497.600 1715.960 ;
        RECT 1.445 1686.040 1497.200 1687.440 ;
        RECT 1.445 1673.840 1497.600 1686.040 ;
        RECT 2.800 1672.440 1497.600 1673.840 ;
        RECT 1.445 1645.960 1497.600 1672.440 ;
        RECT 1.445 1644.560 1497.200 1645.960 ;
        RECT 1.445 1630.320 1497.600 1644.560 ;
        RECT 2.800 1628.920 1497.600 1630.320 ;
        RECT 1.445 1604.480 1497.600 1628.920 ;
        RECT 1.445 1603.080 1497.200 1604.480 ;
        RECT 1.445 1586.800 1497.600 1603.080 ;
        RECT 2.800 1585.400 1497.600 1586.800 ;
        RECT 1.445 1563.000 1497.600 1585.400 ;
        RECT 1.445 1561.600 1497.200 1563.000 ;
        RECT 1.445 1543.280 1497.600 1561.600 ;
        RECT 2.800 1541.880 1497.600 1543.280 ;
        RECT 1.445 1520.840 1497.600 1541.880 ;
        RECT 1.445 1519.440 1497.200 1520.840 ;
        RECT 1.445 1499.760 1497.600 1519.440 ;
        RECT 2.800 1498.360 1497.600 1499.760 ;
        RECT 1.445 1479.360 1497.600 1498.360 ;
        RECT 1.445 1477.960 1497.200 1479.360 ;
        RECT 1.445 1456.240 1497.600 1477.960 ;
        RECT 2.800 1454.840 1497.600 1456.240 ;
        RECT 1.445 1437.880 1497.600 1454.840 ;
        RECT 1.445 1436.480 1497.200 1437.880 ;
        RECT 1.445 1412.720 1497.600 1436.480 ;
        RECT 2.800 1411.320 1497.600 1412.720 ;
        RECT 1.445 1395.720 1497.600 1411.320 ;
        RECT 1.445 1394.320 1497.200 1395.720 ;
        RECT 1.445 1369.200 1497.600 1394.320 ;
        RECT 2.800 1367.800 1497.600 1369.200 ;
        RECT 1.445 1354.240 1497.600 1367.800 ;
        RECT 1.445 1352.840 1497.200 1354.240 ;
        RECT 1.445 1326.360 1497.600 1352.840 ;
        RECT 2.800 1324.960 1497.600 1326.360 ;
        RECT 1.445 1312.760 1497.600 1324.960 ;
        RECT 1.445 1311.360 1497.200 1312.760 ;
        RECT 1.445 1282.840 1497.600 1311.360 ;
        RECT 2.800 1281.440 1497.600 1282.840 ;
        RECT 1.445 1271.280 1497.600 1281.440 ;
        RECT 1.445 1269.880 1497.200 1271.280 ;
        RECT 1.445 1239.320 1497.600 1269.880 ;
        RECT 2.800 1237.920 1497.600 1239.320 ;
        RECT 1.445 1229.120 1497.600 1237.920 ;
        RECT 1.445 1227.720 1497.200 1229.120 ;
        RECT 1.445 1195.800 1497.600 1227.720 ;
        RECT 2.800 1194.400 1497.600 1195.800 ;
        RECT 1.445 1187.640 1497.600 1194.400 ;
        RECT 1.445 1186.240 1497.200 1187.640 ;
        RECT 1.445 1152.280 1497.600 1186.240 ;
        RECT 2.800 1150.880 1497.600 1152.280 ;
        RECT 1.445 1146.160 1497.600 1150.880 ;
        RECT 1.445 1144.760 1497.200 1146.160 ;
        RECT 1.445 1108.760 1497.600 1144.760 ;
        RECT 2.800 1107.360 1497.600 1108.760 ;
        RECT 1.445 1104.680 1497.600 1107.360 ;
        RECT 1.445 1103.280 1497.200 1104.680 ;
        RECT 1.445 1065.240 1497.600 1103.280 ;
        RECT 2.800 1063.840 1497.600 1065.240 ;
        RECT 1.445 1062.520 1497.600 1063.840 ;
        RECT 1.445 1061.120 1497.200 1062.520 ;
        RECT 1.445 1021.720 1497.600 1061.120 ;
        RECT 2.800 1021.040 1497.600 1021.720 ;
        RECT 2.800 1020.320 1497.200 1021.040 ;
        RECT 1.445 1019.640 1497.200 1020.320 ;
        RECT 1.445 979.560 1497.600 1019.640 ;
        RECT 1.445 978.200 1497.200 979.560 ;
        RECT 2.800 978.160 1497.200 978.200 ;
        RECT 2.800 976.800 1497.600 978.160 ;
        RECT 1.445 937.400 1497.600 976.800 ;
        RECT 1.445 936.000 1497.200 937.400 ;
        RECT 1.445 934.680 1497.600 936.000 ;
        RECT 2.800 933.280 1497.600 934.680 ;
        RECT 1.445 895.920 1497.600 933.280 ;
        RECT 1.445 894.520 1497.200 895.920 ;
        RECT 1.445 891.160 1497.600 894.520 ;
        RECT 2.800 889.760 1497.600 891.160 ;
        RECT 1.445 854.440 1497.600 889.760 ;
        RECT 1.445 853.040 1497.200 854.440 ;
        RECT 1.445 847.640 1497.600 853.040 ;
        RECT 2.800 846.240 1497.600 847.640 ;
        RECT 1.445 812.960 1497.600 846.240 ;
        RECT 1.445 811.560 1497.200 812.960 ;
        RECT 1.445 804.120 1497.600 811.560 ;
        RECT 2.800 802.720 1497.600 804.120 ;
        RECT 1.445 770.800 1497.600 802.720 ;
        RECT 1.445 769.400 1497.200 770.800 ;
        RECT 1.445 760.600 1497.600 769.400 ;
        RECT 2.800 759.200 1497.600 760.600 ;
        RECT 1.445 729.320 1497.600 759.200 ;
        RECT 1.445 727.920 1497.200 729.320 ;
        RECT 1.445 717.080 1497.600 727.920 ;
        RECT 2.800 715.680 1497.600 717.080 ;
        RECT 1.445 687.840 1497.600 715.680 ;
        RECT 1.445 686.440 1497.200 687.840 ;
        RECT 1.445 674.240 1497.600 686.440 ;
        RECT 2.800 672.840 1497.600 674.240 ;
        RECT 1.445 646.360 1497.600 672.840 ;
        RECT 1.445 644.960 1497.200 646.360 ;
        RECT 1.445 630.720 1497.600 644.960 ;
        RECT 2.800 629.320 1497.600 630.720 ;
        RECT 1.445 604.200 1497.600 629.320 ;
        RECT 1.445 602.800 1497.200 604.200 ;
        RECT 1.445 587.200 1497.600 602.800 ;
        RECT 2.800 585.800 1497.600 587.200 ;
        RECT 1.445 562.720 1497.600 585.800 ;
        RECT 1.445 561.320 1497.200 562.720 ;
        RECT 1.445 543.680 1497.600 561.320 ;
        RECT 2.800 542.280 1497.600 543.680 ;
        RECT 1.445 521.240 1497.600 542.280 ;
        RECT 1.445 519.840 1497.200 521.240 ;
        RECT 1.445 500.160 1497.600 519.840 ;
        RECT 2.800 498.760 1497.600 500.160 ;
        RECT 1.445 479.080 1497.600 498.760 ;
        RECT 1.445 477.680 1497.200 479.080 ;
        RECT 1.445 456.640 1497.600 477.680 ;
        RECT 2.800 455.240 1497.600 456.640 ;
        RECT 1.445 437.600 1497.600 455.240 ;
        RECT 1.445 436.200 1497.200 437.600 ;
        RECT 1.445 413.120 1497.600 436.200 ;
        RECT 2.800 411.720 1497.600 413.120 ;
        RECT 1.445 396.120 1497.600 411.720 ;
        RECT 1.445 394.720 1497.200 396.120 ;
        RECT 1.445 369.600 1497.600 394.720 ;
        RECT 2.800 368.200 1497.600 369.600 ;
        RECT 1.445 354.640 1497.600 368.200 ;
        RECT 1.445 353.240 1497.200 354.640 ;
        RECT 1.445 326.080 1497.600 353.240 ;
        RECT 2.800 324.680 1497.600 326.080 ;
        RECT 1.445 312.480 1497.600 324.680 ;
        RECT 1.445 311.080 1497.200 312.480 ;
        RECT 1.445 282.560 1497.600 311.080 ;
        RECT 2.800 281.160 1497.600 282.560 ;
        RECT 1.445 271.000 1497.600 281.160 ;
        RECT 1.445 269.600 1497.200 271.000 ;
        RECT 1.445 239.040 1497.600 269.600 ;
        RECT 2.800 237.640 1497.600 239.040 ;
        RECT 1.445 229.520 1497.600 237.640 ;
        RECT 1.445 228.120 1497.200 229.520 ;
        RECT 1.445 195.520 1497.600 228.120 ;
        RECT 2.800 194.120 1497.600 195.520 ;
        RECT 1.445 188.040 1497.600 194.120 ;
        RECT 1.445 186.640 1497.200 188.040 ;
        RECT 1.445 152.000 1497.600 186.640 ;
        RECT 2.800 150.600 1497.600 152.000 ;
        RECT 1.445 145.880 1497.600 150.600 ;
        RECT 1.445 144.480 1497.200 145.880 ;
        RECT 1.445 108.480 1497.600 144.480 ;
        RECT 2.800 107.080 1497.600 108.480 ;
        RECT 1.445 104.400 1497.600 107.080 ;
        RECT 1.445 103.000 1497.200 104.400 ;
        RECT 1.445 64.960 1497.600 103.000 ;
        RECT 2.800 63.560 1497.600 64.960 ;
        RECT 1.445 62.920 1497.600 63.560 ;
        RECT 1.445 61.520 1497.200 62.920 ;
        RECT 1.445 22.120 1497.600 61.520 ;
        RECT 2.800 21.440 1497.600 22.120 ;
        RECT 2.800 20.720 1497.200 21.440 ;
        RECT 1.445 20.040 1497.200 20.720 ;
        RECT 1.445 10.715 1497.600 20.040 ;
      LAYER met4 ;
        RECT 81.255 10.640 97.440 1988.560 ;
        RECT 99.840 10.640 1481.840 1988.560 ;
  END
END fwpayload
END LIBRARY

