
`include "fwrisc_formal_opcode_defines.svh"

`utype_auipc(idata, $anyconst, $anyconst);