VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2700.000 BY 3700.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 2.400 571.840 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 2.400 437.200 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3463.960 2700.000 3464.560 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 2.400 369.880 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 2.400 302.560 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3531.280 2700.000 3531.880 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2675.450 0.000 2675.730 2.400 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 2.400 235.240 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 337.270 3697.600 337.550 3700.000 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3598.600 2700.000 3599.200 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2680.510 0.000 2680.790 2.400 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3262.000 2700.000 3262.600 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 2.400 167.920 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2686.030 0.000 2686.310 2.400 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 2.400 100.600 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3665.920 2700.000 3666.520 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 262.290 3697.600 262.570 3700.000 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 187.310 3697.600 187.590 3700.000 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2691.550 0.000 2691.830 2.400 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 112.330 3697.600 112.610 3700.000 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2697.070 0.000 2697.350 2.400 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 2.400 33.960 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 562.210 3697.600 562.490 3700.000 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 37.350 3697.600 37.630 3700.000 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 487.230 3697.600 487.510 3700.000 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2664.410 0.000 2664.690 2.400 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.920 2.400 504.520 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3329.320 2700.000 3329.920 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 412.250 3697.600 412.530 3700.000 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2669.930 0.000 2670.210 2.400 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3396.640 2700.000 3397.240 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 33.360 2700.000 33.960 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2185.560 2700.000 2186.160 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2387.520 2700.000 2388.120 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2589.480 2700.000 2590.080 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2791.440 2700.000 2792.040 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3060.040 2700.000 3060.640 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2662.110 3697.600 2662.390 3700.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2362.190 3697.600 2362.470 3700.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2137.250 3697.600 2137.530 3700.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1912.310 3697.600 1912.590 3700.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1687.370 3697.600 1687.650 3700.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 234.640 2700.000 235.240 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1462.430 3697.600 1462.710 3700.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1237.030 3697.600 1237.310 3700.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1012.090 3697.600 1012.370 3700.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.150 3697.600 787.430 3700.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3665.920 2.400 3666.520 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3329.320 2.400 3329.920 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3127.360 2.400 3127.960 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2925.400 2.400 2926.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2724.120 2.400 2724.720 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2522.160 2.400 2522.760 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 436.600 2700.000 437.200 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2320.200 2.400 2320.800 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 2118.240 2.400 2118.840 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1782.320 2.400 1782.920 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1580.360 2.400 1580.960 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1378.400 2.400 1379.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1176.440 2.400 1177.040 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 974.480 2.400 975.080 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 2.400 773.800 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 638.560 2700.000 639.160 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 840.520 2700.000 841.120 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1041.800 2700.000 1042.400 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1243.760 2700.000 1244.360 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1580.360 2700.000 1580.960 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1782.320 2700.000 1782.920 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1983.600 2700.000 1984.200 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 167.320 2700.000 167.920 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2320.200 2700.000 2320.800 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2522.160 2700.000 2522.760 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2724.120 2700.000 2724.720 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2925.400 2700.000 2926.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3194.680 2700.000 3195.280 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2512.150 3697.600 2512.430 3700.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2212.230 3697.600 2212.510 3700.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1987.290 3697.600 1987.570 3700.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1762.350 3697.600 1762.630 3700.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1537.410 3697.600 1537.690 3700.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 369.280 2700.000 369.880 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1312.010 3697.600 1312.290 3700.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1087.070 3697.600 1087.350 3700.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 862.130 3697.600 862.410 3700.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 637.190 3697.600 637.470 3700.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3531.280 2.400 3531.880 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3194.680 2.400 3195.280 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2992.720 2.400 2993.320 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2791.440 2.400 2792.040 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2589.480 2.400 2590.080 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2387.520 2.400 2388.120 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 571.240 2700.000 571.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2185.560 2.400 2186.160 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1983.600 2.400 1984.200 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1647.680 2.400 1648.280 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1445.720 2.400 1446.320 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1243.760 2.400 1244.360 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1041.800 2.400 1042.400 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 840.520 2.400 841.120 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 2.400 639.160 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 773.200 2700.000 773.800 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 974.480 2700.000 975.080 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1176.440 2700.000 1177.040 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1378.400 2700.000 1379.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1715.000 2700.000 1715.600 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1916.280 2700.000 1916.880 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2118.240 2700.000 2118.840 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 100.000 2700.000 100.600 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2252.880 2700.000 2253.480 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2454.840 2700.000 2455.440 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2656.800 2700.000 2657.400 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2858.080 2700.000 2858.680 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 3127.360 2700.000 3127.960 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2587.130 3697.600 2587.410 3700.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2287.210 3697.600 2287.490 3700.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2062.270 3697.600 2062.550 3700.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1837.330 3697.600 1837.610 3700.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1612.390 3697.600 1612.670 3700.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 301.960 2700.000 302.560 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1387.450 3697.600 1387.730 3700.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1162.050 3697.600 1162.330 3700.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 937.110 3697.600 937.390 3700.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 712.170 3697.600 712.450 3700.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3598.600 2.400 3599.200 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3262.000 2.400 3262.600 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 3060.040 2.400 3060.640 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2858.080 2.400 2858.680 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2656.800 2.400 2657.400 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2454.840 2.400 2455.440 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 503.920 2700.000 504.520 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2252.880 2.400 2253.480 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2050.920 2.400 2051.520 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1715.000 2.400 1715.600 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1513.040 2.400 1513.640 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1311.080 2.400 1311.680 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 1109.120 2.400 1109.720 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 907.840 2.400 908.440 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 2.400 706.480 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 705.880 2700.000 706.480 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 907.840 2700.000 908.440 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1109.120 2700.000 1109.720 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1311.080 2700.000 1311.680 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1647.680 2700.000 1648.280 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1849.640 2700.000 1850.240 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2050.920 2700.000 2051.520 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2203.490 0.000 2203.770 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2219.590 0.000 2219.870 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2236.150 0.000 2236.430 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2252.250 0.000 2252.530 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2268.810 0.000 2269.090 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2284.910 0.000 2285.190 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2301.010 0.000 2301.290 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2317.570 0.000 2317.850 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2333.670 0.000 2333.950 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2349.770 0.000 2350.050 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 739.770 0.000 740.050 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2366.330 0.000 2366.610 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2382.430 0.000 2382.710 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2398.530 0.000 2398.810 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2415.090 0.000 2415.370 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2431.190 0.000 2431.470 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2447.750 0.000 2448.030 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2463.850 0.000 2464.130 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2479.950 0.000 2480.230 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2496.510 0.000 2496.790 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2512.610 0.000 2512.890 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 755.870 0.000 756.150 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2528.710 0.000 2528.990 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2545.270 0.000 2545.550 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2561.370 0.000 2561.650 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2577.470 0.000 2577.750 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2594.030 0.000 2594.310 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2610.130 0.000 2610.410 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2626.230 0.000 2626.510 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2642.790 0.000 2643.070 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 771.970 0.000 772.250 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 788.530 0.000 788.810 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 804.630 0.000 804.910 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 820.730 0.000 821.010 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 837.290 0.000 837.570 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 869.490 0.000 869.770 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 886.050 0.000 886.330 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 593.030 0.000 593.310 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 902.150 0.000 902.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 918.710 0.000 918.990 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 934.810 0.000 935.090 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 950.910 0.000 951.190 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 967.470 0.000 967.750 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.570 0.000 983.850 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 999.670 0.000 999.950 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1016.230 0.000 1016.510 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.330 0.000 1032.610 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1048.430 0.000 1048.710 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1064.990 0.000 1065.270 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1081.090 0.000 1081.370 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1097.650 0.000 1097.930 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1113.750 0.000 1114.030 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1129.850 0.000 1130.130 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.510 0.000 1162.790 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1178.610 0.000 1178.890 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1211.270 0.000 1211.550 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1227.370 0.000 1227.650 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1243.930 0.000 1244.210 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1260.030 0.000 1260.310 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1276.130 0.000 1276.410 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1292.690 0.000 1292.970 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1308.790 0.000 1309.070 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1325.350 0.000 1325.630 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1341.450 0.000 1341.730 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1357.550 0.000 1357.830 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1374.110 0.000 1374.390 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 641.790 0.000 642.070 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1390.210 0.000 1390.490 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1406.310 0.000 1406.590 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1422.870 0.000 1423.150 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1438.970 0.000 1439.250 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1455.070 0.000 1455.350 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1471.630 0.000 1471.910 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1487.730 0.000 1488.010 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1504.290 0.000 1504.570 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1520.390 0.000 1520.670 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1536.490 0.000 1536.770 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 658.350 0.000 658.630 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1553.050 0.000 1553.330 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1569.150 0.000 1569.430 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1585.250 0.000 1585.530 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1601.810 0.000 1602.090 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1617.910 0.000 1618.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1634.010 0.000 1634.290 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1650.570 0.000 1650.850 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1666.670 0.000 1666.950 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1683.230 0.000 1683.510 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1699.330 0.000 1699.610 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 674.450 0.000 674.730 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1715.430 0.000 1715.710 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1731.990 0.000 1732.270 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1748.090 0.000 1748.370 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1764.190 0.000 1764.470 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1780.750 0.000 1781.030 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1796.850 0.000 1797.130 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1812.950 0.000 1813.230 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1829.510 0.000 1829.790 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1845.610 0.000 1845.890 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1861.710 0.000 1861.990 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 690.550 0.000 690.830 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1878.270 0.000 1878.550 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1894.370 0.000 1894.650 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1910.930 0.000 1911.210 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1927.030 0.000 1927.310 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1943.130 0.000 1943.410 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1959.690 0.000 1959.970 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1975.790 0.000 1976.070 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1991.890 0.000 1992.170 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2008.450 0.000 2008.730 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2024.550 0.000 2024.830 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 707.110 0.000 707.390 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2040.650 0.000 2040.930 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2057.210 0.000 2057.490 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2073.310 0.000 2073.590 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2089.870 0.000 2090.150 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2105.970 0.000 2106.250 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2122.070 0.000 2122.350 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2138.630 0.000 2138.910 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2154.730 0.000 2155.010 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2170.830 0.000 2171.110 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2187.390 0.000 2187.670 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 723.210 0.000 723.490 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 582.450 0.000 582.730 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2209.010 0.000 2209.290 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2225.110 0.000 2225.390 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2241.670 0.000 2241.950 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2257.770 0.000 2258.050 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2273.870 0.000 2274.150 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2290.430 0.000 2290.710 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2306.530 0.000 2306.810 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2322.630 0.000 2322.910 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2339.190 0.000 2339.470 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2355.290 0.000 2355.570 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 744.830 0.000 745.110 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2371.390 0.000 2371.670 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2387.950 0.000 2388.230 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2404.050 0.000 2404.330 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2420.610 0.000 2420.890 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2436.710 0.000 2436.990 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2452.810 0.000 2453.090 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2469.370 0.000 2469.650 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2485.470 0.000 2485.750 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2501.570 0.000 2501.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2518.130 0.000 2518.410 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 761.390 0.000 761.670 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2534.230 0.000 2534.510 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2550.330 0.000 2550.610 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2566.890 0.000 2567.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2582.990 0.000 2583.270 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2599.550 0.000 2599.830 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2615.650 0.000 2615.930 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2631.750 0.000 2632.030 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2648.310 0.000 2648.590 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 777.490 0.000 777.770 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 810.150 0.000 810.430 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 826.250 0.000 826.530 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 842.810 0.000 843.090 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 858.910 0.000 859.190 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 875.010 0.000 875.290 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 891.570 0.000 891.850 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 598.550 0.000 598.830 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 907.670 0.000 907.950 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 923.770 0.000 924.050 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 940.330 0.000 940.610 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 972.530 0.000 972.810 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 989.090 0.000 989.370 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1005.190 0.000 1005.470 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1021.290 0.000 1021.570 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1037.850 0.000 1038.130 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1053.950 0.000 1054.230 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1070.510 0.000 1070.790 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1086.610 0.000 1086.890 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1102.710 0.000 1102.990 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1119.270 0.000 1119.550 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1135.370 0.000 1135.650 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1151.470 0.000 1151.750 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1168.030 0.000 1168.310 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1184.130 0.000 1184.410 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1200.230 0.000 1200.510 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1216.790 0.000 1217.070 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1232.890 0.000 1233.170 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1249.450 0.000 1249.730 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1281.650 0.000 1281.930 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1298.210 0.000 1298.490 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1314.310 0.000 1314.590 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1330.410 0.000 1330.690 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1346.970 0.000 1347.250 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1363.070 0.000 1363.350 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1379.170 0.000 1379.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1395.730 0.000 1396.010 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1411.830 0.000 1412.110 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1428.390 0.000 1428.670 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1444.490 0.000 1444.770 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1460.590 0.000 1460.870 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1477.150 0.000 1477.430 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1493.250 0.000 1493.530 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1509.350 0.000 1509.630 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1525.910 0.000 1526.190 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1542.010 0.000 1542.290 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 663.870 0.000 664.150 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1558.110 0.000 1558.390 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1574.670 0.000 1574.950 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1590.770 0.000 1591.050 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1606.870 0.000 1607.150 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1623.430 0.000 1623.710 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1639.530 0.000 1639.810 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1656.090 0.000 1656.370 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1672.190 0.000 1672.470 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1688.290 0.000 1688.570 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1704.850 0.000 1705.130 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 679.970 0.000 680.250 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1720.950 0.000 1721.230 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1737.050 0.000 1737.330 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1753.610 0.000 1753.890 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1769.710 0.000 1769.990 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1785.810 0.000 1786.090 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1802.370 0.000 1802.650 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1818.470 0.000 1818.750 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1835.030 0.000 1835.310 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1851.130 0.000 1851.410 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1867.230 0.000 1867.510 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 696.070 0.000 696.350 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1883.790 0.000 1884.070 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1899.890 0.000 1900.170 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1915.990 0.000 1916.270 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1932.550 0.000 1932.830 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1948.650 0.000 1948.930 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1964.750 0.000 1965.030 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1981.310 0.000 1981.590 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1997.410 0.000 1997.690 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2013.970 0.000 2014.250 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2030.070 0.000 2030.350 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 712.630 0.000 712.910 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2046.170 0.000 2046.450 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2062.730 0.000 2063.010 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2078.830 0.000 2079.110 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2094.930 0.000 2095.210 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2111.490 0.000 2111.770 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2127.590 0.000 2127.870 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2143.690 0.000 2143.970 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2160.250 0.000 2160.530 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2176.350 0.000 2176.630 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2192.910 0.000 2193.190 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 728.730 0.000 729.010 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.970 0.000 588.250 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2214.530 0.000 2214.810 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2230.630 0.000 2230.910 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2246.730 0.000 2247.010 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2263.290 0.000 2263.570 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2279.390 0.000 2279.670 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2295.490 0.000 2295.770 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2312.050 0.000 2312.330 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2328.150 0.000 2328.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2344.710 0.000 2344.990 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2360.810 0.000 2361.090 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 750.350 0.000 750.630 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2376.910 0.000 2377.190 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2393.470 0.000 2393.750 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2409.570 0.000 2409.850 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2425.670 0.000 2425.950 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2442.230 0.000 2442.510 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2458.330 0.000 2458.610 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2474.430 0.000 2474.710 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2490.990 0.000 2491.270 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2507.090 0.000 2507.370 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2523.650 0.000 2523.930 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2539.750 0.000 2540.030 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2555.850 0.000 2556.130 2.400 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2572.410 0.000 2572.690 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2588.510 0.000 2588.790 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2604.610 0.000 2604.890 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2621.170 0.000 2621.450 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2637.270 0.000 2637.550 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2653.370 0.000 2653.650 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.010 0.000 783.290 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 799.110 0.000 799.390 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 815.670 0.000 815.950 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 831.770 0.000 832.050 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 847.870 0.000 848.150 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.430 0.000 864.710 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 880.530 0.000 880.810 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.630 0.000 896.910 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 913.190 0.000 913.470 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.290 0.000 929.570 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 945.390 0.000 945.670 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 961.950 0.000 962.230 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 978.050 0.000 978.330 2.400 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 994.610 0.000 994.890 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1010.710 0.000 1010.990 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1026.810 0.000 1027.090 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.370 0.000 1043.650 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1059.470 0.000 1059.750 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 620.170 0.000 620.450 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1092.130 0.000 1092.410 2.400 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1108.230 0.000 1108.510 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1124.330 0.000 1124.610 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1140.890 0.000 1141.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1156.990 0.000 1157.270 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1173.550 0.000 1173.830 2.400 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1189.650 0.000 1189.930 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1205.750 0.000 1206.030 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1222.310 0.000 1222.590 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 636.730 0.000 637.010 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1238.410 0.000 1238.690 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1254.510 0.000 1254.790 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1271.070 0.000 1271.350 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.170 0.000 1287.450 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1303.270 0.000 1303.550 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1319.830 0.000 1320.110 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1335.930 0.000 1336.210 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1352.490 0.000 1352.770 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1368.590 0.000 1368.870 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1384.690 0.000 1384.970 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 652.830 0.000 653.110 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1401.250 0.000 1401.530 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1417.350 0.000 1417.630 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1433.450 0.000 1433.730 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1450.010 0.000 1450.290 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1466.110 0.000 1466.390 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1482.210 0.000 1482.490 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1498.770 0.000 1499.050 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1514.870 0.000 1515.150 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1530.970 0.000 1531.250 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1547.530 0.000 1547.810 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.930 0.000 669.210 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1563.630 0.000 1563.910 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1580.190 0.000 1580.470 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1596.290 0.000 1596.570 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1612.390 0.000 1612.670 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1628.950 0.000 1629.230 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1645.050 0.000 1645.330 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1661.150 0.000 1661.430 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1677.710 0.000 1677.990 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1693.810 0.000 1694.090 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1709.910 0.000 1710.190 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 685.490 0.000 685.770 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1726.470 0.000 1726.750 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1742.570 0.000 1742.850 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1759.130 0.000 1759.410 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1775.230 0.000 1775.510 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1791.330 0.000 1791.610 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1807.890 0.000 1808.170 2.400 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1823.990 0.000 1824.270 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1840.090 0.000 1840.370 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1856.650 0.000 1856.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1872.750 0.000 1873.030 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 701.590 0.000 701.870 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1888.850 0.000 1889.130 2.400 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1905.410 0.000 1905.690 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1921.510 0.000 1921.790 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1938.070 0.000 1938.350 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1954.170 0.000 1954.450 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1970.270 0.000 1970.550 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1986.830 0.000 1987.110 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2002.930 0.000 2003.210 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2019.030 0.000 2019.310 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2035.590 0.000 2035.870 2.400 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2051.690 0.000 2051.970 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2067.790 0.000 2068.070 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2084.350 0.000 2084.630 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2100.450 0.000 2100.730 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2116.550 0.000 2116.830 2.400 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2133.110 0.000 2133.390 2.400 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2149.210 0.000 2149.490 2.400 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2165.770 0.000 2166.050 2.400 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2181.870 0.000 2182.150 2.400 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2197.970 0.000 2198.250 2.400 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2658.890 0.000 2659.170 2.400 ;
    END
  END user_clock2
  PIN vccd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 2992.720 2700.000 2993.320 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3463.960 2.400 3464.560 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1513.040 2700.000 1513.640 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1916.280 2.400 1916.880 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2437.170 3697.600 2437.450 3700.000 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3396.640 2.400 3397.240 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2697.600 1445.720 2700.000 1446.320 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 1849.640 2.400 1850.240 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 251.710 0.000 251.990 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 283.910 0.000 284.190 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 349.230 0.000 349.510 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 381.890 0.000 382.170 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 397.990 0.000 398.270 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.090 0.000 414.370 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 446.750 0.000 447.030 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 462.850 0.000 463.130 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.290 0.000 78.570 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 544.270 0.000 544.550 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 560.830 0.000 561.110 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 137.630 0.000 137.910 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 0.000 170.570 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 273.330 0.000 273.610 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 305.990 0.000 306.270 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 354.750 0.000 355.030 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 370.850 0.000 371.130 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 0.000 62.010 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.510 0.000 403.790 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 435.710 0.000 435.990 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 468.370 0.000 468.650 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 501.030 0.000 501.310 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 517.130 0.000 517.410 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 549.790 0.000 550.070 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 565.890 0.000 566.170 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.150 0.000 143.430 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 376.370 0.000 376.650 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.250 0.000 67.530 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.470 0.000 392.750 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 473.890 0.000 474.170 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 522.650 0.000 522.930 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 538.750 0.000 539.030 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 148.670 0.000 148.950 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 72.770 0.000 73.050 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.400 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 2694.220 28.090 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 2694.220 104.680 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2694.220 3688.405 ;
      LAYER met1 ;
        RECT 2.370 2.760 2694.220 3688.560 ;
      LAYER met2 ;
        RECT 2.400 3697.320 37.070 3697.600 ;
        RECT 37.910 3697.320 112.050 3697.600 ;
        RECT 112.890 3697.320 187.030 3697.600 ;
        RECT 187.870 3697.320 262.010 3697.600 ;
        RECT 262.850 3697.320 336.990 3697.600 ;
        RECT 337.830 3697.320 411.970 3697.600 ;
        RECT 412.810 3697.320 486.950 3697.600 ;
        RECT 487.790 3697.320 561.930 3697.600 ;
        RECT 562.770 3697.320 636.910 3697.600 ;
        RECT 637.750 3697.320 711.890 3697.600 ;
        RECT 712.730 3697.320 786.870 3697.600 ;
        RECT 787.710 3697.320 861.850 3697.600 ;
        RECT 862.690 3697.320 936.830 3697.600 ;
        RECT 937.670 3697.320 1011.810 3697.600 ;
        RECT 1012.650 3697.320 1086.790 3697.600 ;
        RECT 1087.630 3697.320 1161.770 3697.600 ;
        RECT 1162.610 3697.320 1236.750 3697.600 ;
        RECT 1237.590 3697.320 1311.730 3697.600 ;
        RECT 1312.570 3697.320 1387.170 3697.600 ;
        RECT 1388.010 3697.320 1462.150 3697.600 ;
        RECT 1462.990 3697.320 1537.130 3697.600 ;
        RECT 1537.970 3697.320 1612.110 3697.600 ;
        RECT 1612.950 3697.320 1687.090 3697.600 ;
        RECT 1687.930 3697.320 1762.070 3697.600 ;
        RECT 1762.910 3697.320 1837.050 3697.600 ;
        RECT 1837.890 3697.320 1912.030 3697.600 ;
        RECT 1912.870 3697.320 1987.010 3697.600 ;
        RECT 1987.850 3697.320 2061.990 3697.600 ;
        RECT 2062.830 3697.320 2136.970 3697.600 ;
        RECT 2137.810 3697.320 2211.950 3697.600 ;
        RECT 2212.790 3697.320 2286.930 3697.600 ;
        RECT 2287.770 3697.320 2361.910 3697.600 ;
        RECT 2362.750 3697.320 2436.890 3697.600 ;
        RECT 2437.730 3697.320 2511.870 3697.600 ;
        RECT 2512.710 3697.320 2586.850 3697.600 ;
        RECT 2587.690 3697.320 2661.830 3697.600 ;
        RECT 2662.670 3697.320 2689.070 3697.600 ;
        RECT 2.400 2.680 2689.070 3697.320 ;
        RECT 2.950 2.400 7.170 2.680 ;
        RECT 8.010 2.400 12.690 2.680 ;
        RECT 13.530 2.400 18.210 2.680 ;
        RECT 19.050 2.400 23.730 2.680 ;
        RECT 24.570 2.400 28.790 2.680 ;
        RECT 29.630 2.400 34.310 2.680 ;
        RECT 35.150 2.400 39.830 2.680 ;
        RECT 40.670 2.400 45.350 2.680 ;
        RECT 46.190 2.400 50.870 2.680 ;
        RECT 51.710 2.400 55.930 2.680 ;
        RECT 56.770 2.400 61.450 2.680 ;
        RECT 62.290 2.400 66.970 2.680 ;
        RECT 67.810 2.400 72.490 2.680 ;
        RECT 73.330 2.400 78.010 2.680 ;
        RECT 78.850 2.400 83.070 2.680 ;
        RECT 83.910 2.400 88.590 2.680 ;
        RECT 89.430 2.400 94.110 2.680 ;
        RECT 94.950 2.400 99.630 2.680 ;
        RECT 100.470 2.400 104.690 2.680 ;
        RECT 105.530 2.400 110.210 2.680 ;
        RECT 111.050 2.400 115.730 2.680 ;
        RECT 116.570 2.400 121.250 2.680 ;
        RECT 122.090 2.400 126.770 2.680 ;
        RECT 127.610 2.400 131.830 2.680 ;
        RECT 132.670 2.400 137.350 2.680 ;
        RECT 138.190 2.400 142.870 2.680 ;
        RECT 143.710 2.400 148.390 2.680 ;
        RECT 149.230 2.400 153.910 2.680 ;
        RECT 154.750 2.400 158.970 2.680 ;
        RECT 159.810 2.400 164.490 2.680 ;
        RECT 165.330 2.400 170.010 2.680 ;
        RECT 170.850 2.400 175.530 2.680 ;
        RECT 176.370 2.400 180.590 2.680 ;
        RECT 181.430 2.400 186.110 2.680 ;
        RECT 186.950 2.400 191.630 2.680 ;
        RECT 192.470 2.400 197.150 2.680 ;
        RECT 197.990 2.400 202.670 2.680 ;
        RECT 203.510 2.400 207.730 2.680 ;
        RECT 208.570 2.400 213.250 2.680 ;
        RECT 214.090 2.400 218.770 2.680 ;
        RECT 219.610 2.400 224.290 2.680 ;
        RECT 225.130 2.400 229.810 2.680 ;
        RECT 230.650 2.400 234.870 2.680 ;
        RECT 235.710 2.400 240.390 2.680 ;
        RECT 241.230 2.400 245.910 2.680 ;
        RECT 246.750 2.400 251.430 2.680 ;
        RECT 252.270 2.400 256.490 2.680 ;
        RECT 257.330 2.400 262.010 2.680 ;
        RECT 262.850 2.400 267.530 2.680 ;
        RECT 268.370 2.400 273.050 2.680 ;
        RECT 273.890 2.400 278.570 2.680 ;
        RECT 279.410 2.400 283.630 2.680 ;
        RECT 284.470 2.400 289.150 2.680 ;
        RECT 289.990 2.400 294.670 2.680 ;
        RECT 295.510 2.400 300.190 2.680 ;
        RECT 301.030 2.400 305.710 2.680 ;
        RECT 306.550 2.400 310.770 2.680 ;
        RECT 311.610 2.400 316.290 2.680 ;
        RECT 317.130 2.400 321.810 2.680 ;
        RECT 322.650 2.400 327.330 2.680 ;
        RECT 328.170 2.400 332.850 2.680 ;
        RECT 333.690 2.400 337.910 2.680 ;
        RECT 338.750 2.400 343.430 2.680 ;
        RECT 344.270 2.400 348.950 2.680 ;
        RECT 349.790 2.400 354.470 2.680 ;
        RECT 355.310 2.400 359.530 2.680 ;
        RECT 360.370 2.400 365.050 2.680 ;
        RECT 365.890 2.400 370.570 2.680 ;
        RECT 371.410 2.400 376.090 2.680 ;
        RECT 376.930 2.400 381.610 2.680 ;
        RECT 382.450 2.400 386.670 2.680 ;
        RECT 387.510 2.400 392.190 2.680 ;
        RECT 393.030 2.400 397.710 2.680 ;
        RECT 398.550 2.400 403.230 2.680 ;
        RECT 404.070 2.400 408.750 2.680 ;
        RECT 409.590 2.400 413.810 2.680 ;
        RECT 414.650 2.400 419.330 2.680 ;
        RECT 420.170 2.400 424.850 2.680 ;
        RECT 425.690 2.400 430.370 2.680 ;
        RECT 431.210 2.400 435.430 2.680 ;
        RECT 436.270 2.400 440.950 2.680 ;
        RECT 441.790 2.400 446.470 2.680 ;
        RECT 447.310 2.400 451.990 2.680 ;
        RECT 452.830 2.400 457.510 2.680 ;
        RECT 458.350 2.400 462.570 2.680 ;
        RECT 463.410 2.400 468.090 2.680 ;
        RECT 468.930 2.400 473.610 2.680 ;
        RECT 474.450 2.400 479.130 2.680 ;
        RECT 479.970 2.400 484.650 2.680 ;
        RECT 485.490 2.400 489.710 2.680 ;
        RECT 490.550 2.400 495.230 2.680 ;
        RECT 496.070 2.400 500.750 2.680 ;
        RECT 501.590 2.400 506.270 2.680 ;
        RECT 507.110 2.400 511.330 2.680 ;
        RECT 512.170 2.400 516.850 2.680 ;
        RECT 517.690 2.400 522.370 2.680 ;
        RECT 523.210 2.400 527.890 2.680 ;
        RECT 528.730 2.400 533.410 2.680 ;
        RECT 534.250 2.400 538.470 2.680 ;
        RECT 539.310 2.400 543.990 2.680 ;
        RECT 544.830 2.400 549.510 2.680 ;
        RECT 550.350 2.400 555.030 2.680 ;
        RECT 555.870 2.400 560.550 2.680 ;
        RECT 561.390 2.400 565.610 2.680 ;
        RECT 566.450 2.400 571.130 2.680 ;
        RECT 571.970 2.400 576.650 2.680 ;
        RECT 577.490 2.400 582.170 2.680 ;
        RECT 583.010 2.400 587.690 2.680 ;
        RECT 588.530 2.400 592.750 2.680 ;
        RECT 593.590 2.400 598.270 2.680 ;
        RECT 599.110 2.400 603.790 2.680 ;
        RECT 604.630 2.400 609.310 2.680 ;
        RECT 610.150 2.400 614.370 2.680 ;
        RECT 615.210 2.400 619.890 2.680 ;
        RECT 620.730 2.400 625.410 2.680 ;
        RECT 626.250 2.400 630.930 2.680 ;
        RECT 631.770 2.400 636.450 2.680 ;
        RECT 637.290 2.400 641.510 2.680 ;
        RECT 642.350 2.400 647.030 2.680 ;
        RECT 647.870 2.400 652.550 2.680 ;
        RECT 653.390 2.400 658.070 2.680 ;
        RECT 658.910 2.400 663.590 2.680 ;
        RECT 664.430 2.400 668.650 2.680 ;
        RECT 669.490 2.400 674.170 2.680 ;
        RECT 675.010 2.400 679.690 2.680 ;
        RECT 680.530 2.400 685.210 2.680 ;
        RECT 686.050 2.400 690.270 2.680 ;
        RECT 691.110 2.400 695.790 2.680 ;
        RECT 696.630 2.400 701.310 2.680 ;
        RECT 702.150 2.400 706.830 2.680 ;
        RECT 707.670 2.400 712.350 2.680 ;
        RECT 713.190 2.400 717.410 2.680 ;
        RECT 718.250 2.400 722.930 2.680 ;
        RECT 723.770 2.400 728.450 2.680 ;
        RECT 729.290 2.400 733.970 2.680 ;
        RECT 734.810 2.400 739.490 2.680 ;
        RECT 740.330 2.400 744.550 2.680 ;
        RECT 745.390 2.400 750.070 2.680 ;
        RECT 750.910 2.400 755.590 2.680 ;
        RECT 756.430 2.400 761.110 2.680 ;
        RECT 761.950 2.400 766.170 2.680 ;
        RECT 767.010 2.400 771.690 2.680 ;
        RECT 772.530 2.400 777.210 2.680 ;
        RECT 778.050 2.400 782.730 2.680 ;
        RECT 783.570 2.400 788.250 2.680 ;
        RECT 789.090 2.400 793.310 2.680 ;
        RECT 794.150 2.400 798.830 2.680 ;
        RECT 799.670 2.400 804.350 2.680 ;
        RECT 805.190 2.400 809.870 2.680 ;
        RECT 810.710 2.400 815.390 2.680 ;
        RECT 816.230 2.400 820.450 2.680 ;
        RECT 821.290 2.400 825.970 2.680 ;
        RECT 826.810 2.400 831.490 2.680 ;
        RECT 832.330 2.400 837.010 2.680 ;
        RECT 837.850 2.400 842.530 2.680 ;
        RECT 843.370 2.400 847.590 2.680 ;
        RECT 848.430 2.400 853.110 2.680 ;
        RECT 853.950 2.400 858.630 2.680 ;
        RECT 859.470 2.400 864.150 2.680 ;
        RECT 864.990 2.400 869.210 2.680 ;
        RECT 870.050 2.400 874.730 2.680 ;
        RECT 875.570 2.400 880.250 2.680 ;
        RECT 881.090 2.400 885.770 2.680 ;
        RECT 886.610 2.400 891.290 2.680 ;
        RECT 892.130 2.400 896.350 2.680 ;
        RECT 897.190 2.400 901.870 2.680 ;
        RECT 902.710 2.400 907.390 2.680 ;
        RECT 908.230 2.400 912.910 2.680 ;
        RECT 913.750 2.400 918.430 2.680 ;
        RECT 919.270 2.400 923.490 2.680 ;
        RECT 924.330 2.400 929.010 2.680 ;
        RECT 929.850 2.400 934.530 2.680 ;
        RECT 935.370 2.400 940.050 2.680 ;
        RECT 940.890 2.400 945.110 2.680 ;
        RECT 945.950 2.400 950.630 2.680 ;
        RECT 951.470 2.400 956.150 2.680 ;
        RECT 956.990 2.400 961.670 2.680 ;
        RECT 962.510 2.400 967.190 2.680 ;
        RECT 968.030 2.400 972.250 2.680 ;
        RECT 973.090 2.400 977.770 2.680 ;
        RECT 978.610 2.400 983.290 2.680 ;
        RECT 984.130 2.400 988.810 2.680 ;
        RECT 989.650 2.400 994.330 2.680 ;
        RECT 995.170 2.400 999.390 2.680 ;
        RECT 1000.230 2.400 1004.910 2.680 ;
        RECT 1005.750 2.400 1010.430 2.680 ;
        RECT 1011.270 2.400 1015.950 2.680 ;
        RECT 1016.790 2.400 1021.010 2.680 ;
        RECT 1021.850 2.400 1026.530 2.680 ;
        RECT 1027.370 2.400 1032.050 2.680 ;
        RECT 1032.890 2.400 1037.570 2.680 ;
        RECT 1038.410 2.400 1043.090 2.680 ;
        RECT 1043.930 2.400 1048.150 2.680 ;
        RECT 1048.990 2.400 1053.670 2.680 ;
        RECT 1054.510 2.400 1059.190 2.680 ;
        RECT 1060.030 2.400 1064.710 2.680 ;
        RECT 1065.550 2.400 1070.230 2.680 ;
        RECT 1071.070 2.400 1075.290 2.680 ;
        RECT 1076.130 2.400 1080.810 2.680 ;
        RECT 1081.650 2.400 1086.330 2.680 ;
        RECT 1087.170 2.400 1091.850 2.680 ;
        RECT 1092.690 2.400 1097.370 2.680 ;
        RECT 1098.210 2.400 1102.430 2.680 ;
        RECT 1103.270 2.400 1107.950 2.680 ;
        RECT 1108.790 2.400 1113.470 2.680 ;
        RECT 1114.310 2.400 1118.990 2.680 ;
        RECT 1119.830 2.400 1124.050 2.680 ;
        RECT 1124.890 2.400 1129.570 2.680 ;
        RECT 1130.410 2.400 1135.090 2.680 ;
        RECT 1135.930 2.400 1140.610 2.680 ;
        RECT 1141.450 2.400 1146.130 2.680 ;
        RECT 1146.970 2.400 1151.190 2.680 ;
        RECT 1152.030 2.400 1156.710 2.680 ;
        RECT 1157.550 2.400 1162.230 2.680 ;
        RECT 1163.070 2.400 1167.750 2.680 ;
        RECT 1168.590 2.400 1173.270 2.680 ;
        RECT 1174.110 2.400 1178.330 2.680 ;
        RECT 1179.170 2.400 1183.850 2.680 ;
        RECT 1184.690 2.400 1189.370 2.680 ;
        RECT 1190.210 2.400 1194.890 2.680 ;
        RECT 1195.730 2.400 1199.950 2.680 ;
        RECT 1200.790 2.400 1205.470 2.680 ;
        RECT 1206.310 2.400 1210.990 2.680 ;
        RECT 1211.830 2.400 1216.510 2.680 ;
        RECT 1217.350 2.400 1222.030 2.680 ;
        RECT 1222.870 2.400 1227.090 2.680 ;
        RECT 1227.930 2.400 1232.610 2.680 ;
        RECT 1233.450 2.400 1238.130 2.680 ;
        RECT 1238.970 2.400 1243.650 2.680 ;
        RECT 1244.490 2.400 1249.170 2.680 ;
        RECT 1250.010 2.400 1254.230 2.680 ;
        RECT 1255.070 2.400 1259.750 2.680 ;
        RECT 1260.590 2.400 1265.270 2.680 ;
        RECT 1266.110 2.400 1270.790 2.680 ;
        RECT 1271.630 2.400 1275.850 2.680 ;
        RECT 1276.690 2.400 1281.370 2.680 ;
        RECT 1282.210 2.400 1286.890 2.680 ;
        RECT 1287.730 2.400 1292.410 2.680 ;
        RECT 1293.250 2.400 1297.930 2.680 ;
        RECT 1298.770 2.400 1302.990 2.680 ;
        RECT 1303.830 2.400 1308.510 2.680 ;
        RECT 1309.350 2.400 1314.030 2.680 ;
        RECT 1314.870 2.400 1319.550 2.680 ;
        RECT 1320.390 2.400 1325.070 2.680 ;
        RECT 1325.910 2.400 1330.130 2.680 ;
        RECT 1330.970 2.400 1335.650 2.680 ;
        RECT 1336.490 2.400 1341.170 2.680 ;
        RECT 1342.010 2.400 1346.690 2.680 ;
        RECT 1347.530 2.400 1352.210 2.680 ;
        RECT 1353.050 2.400 1357.270 2.680 ;
        RECT 1358.110 2.400 1362.790 2.680 ;
        RECT 1363.630 2.400 1368.310 2.680 ;
        RECT 1369.150 2.400 1373.830 2.680 ;
        RECT 1374.670 2.400 1378.890 2.680 ;
        RECT 1379.730 2.400 1384.410 2.680 ;
        RECT 1385.250 2.400 1389.930 2.680 ;
        RECT 1390.770 2.400 1395.450 2.680 ;
        RECT 1396.290 2.400 1400.970 2.680 ;
        RECT 1401.810 2.400 1406.030 2.680 ;
        RECT 1406.870 2.400 1411.550 2.680 ;
        RECT 1412.390 2.400 1417.070 2.680 ;
        RECT 1417.910 2.400 1422.590 2.680 ;
        RECT 1423.430 2.400 1428.110 2.680 ;
        RECT 1428.950 2.400 1433.170 2.680 ;
        RECT 1434.010 2.400 1438.690 2.680 ;
        RECT 1439.530 2.400 1444.210 2.680 ;
        RECT 1445.050 2.400 1449.730 2.680 ;
        RECT 1450.570 2.400 1454.790 2.680 ;
        RECT 1455.630 2.400 1460.310 2.680 ;
        RECT 1461.150 2.400 1465.830 2.680 ;
        RECT 1466.670 2.400 1471.350 2.680 ;
        RECT 1472.190 2.400 1476.870 2.680 ;
        RECT 1477.710 2.400 1481.930 2.680 ;
        RECT 1482.770 2.400 1487.450 2.680 ;
        RECT 1488.290 2.400 1492.970 2.680 ;
        RECT 1493.810 2.400 1498.490 2.680 ;
        RECT 1499.330 2.400 1504.010 2.680 ;
        RECT 1504.850 2.400 1509.070 2.680 ;
        RECT 1509.910 2.400 1514.590 2.680 ;
        RECT 1515.430 2.400 1520.110 2.680 ;
        RECT 1520.950 2.400 1525.630 2.680 ;
        RECT 1526.470 2.400 1530.690 2.680 ;
        RECT 1531.530 2.400 1536.210 2.680 ;
        RECT 1537.050 2.400 1541.730 2.680 ;
        RECT 1542.570 2.400 1547.250 2.680 ;
        RECT 1548.090 2.400 1552.770 2.680 ;
        RECT 1553.610 2.400 1557.830 2.680 ;
        RECT 1558.670 2.400 1563.350 2.680 ;
        RECT 1564.190 2.400 1568.870 2.680 ;
        RECT 1569.710 2.400 1574.390 2.680 ;
        RECT 1575.230 2.400 1579.910 2.680 ;
        RECT 1580.750 2.400 1584.970 2.680 ;
        RECT 1585.810 2.400 1590.490 2.680 ;
        RECT 1591.330 2.400 1596.010 2.680 ;
        RECT 1596.850 2.400 1601.530 2.680 ;
        RECT 1602.370 2.400 1606.590 2.680 ;
        RECT 1607.430 2.400 1612.110 2.680 ;
        RECT 1612.950 2.400 1617.630 2.680 ;
        RECT 1618.470 2.400 1623.150 2.680 ;
        RECT 1623.990 2.400 1628.670 2.680 ;
        RECT 1629.510 2.400 1633.730 2.680 ;
        RECT 1634.570 2.400 1639.250 2.680 ;
        RECT 1640.090 2.400 1644.770 2.680 ;
        RECT 1645.610 2.400 1650.290 2.680 ;
        RECT 1651.130 2.400 1655.810 2.680 ;
        RECT 1656.650 2.400 1660.870 2.680 ;
        RECT 1661.710 2.400 1666.390 2.680 ;
        RECT 1667.230 2.400 1671.910 2.680 ;
        RECT 1672.750 2.400 1677.430 2.680 ;
        RECT 1678.270 2.400 1682.950 2.680 ;
        RECT 1683.790 2.400 1688.010 2.680 ;
        RECT 1688.850 2.400 1693.530 2.680 ;
        RECT 1694.370 2.400 1699.050 2.680 ;
        RECT 1699.890 2.400 1704.570 2.680 ;
        RECT 1705.410 2.400 1709.630 2.680 ;
        RECT 1710.470 2.400 1715.150 2.680 ;
        RECT 1715.990 2.400 1720.670 2.680 ;
        RECT 1721.510 2.400 1726.190 2.680 ;
        RECT 1727.030 2.400 1731.710 2.680 ;
        RECT 1732.550 2.400 1736.770 2.680 ;
        RECT 1737.610 2.400 1742.290 2.680 ;
        RECT 1743.130 2.400 1747.810 2.680 ;
        RECT 1748.650 2.400 1753.330 2.680 ;
        RECT 1754.170 2.400 1758.850 2.680 ;
        RECT 1759.690 2.400 1763.910 2.680 ;
        RECT 1764.750 2.400 1769.430 2.680 ;
        RECT 1770.270 2.400 1774.950 2.680 ;
        RECT 1775.790 2.400 1780.470 2.680 ;
        RECT 1781.310 2.400 1785.530 2.680 ;
        RECT 1786.370 2.400 1791.050 2.680 ;
        RECT 1791.890 2.400 1796.570 2.680 ;
        RECT 1797.410 2.400 1802.090 2.680 ;
        RECT 1802.930 2.400 1807.610 2.680 ;
        RECT 1808.450 2.400 1812.670 2.680 ;
        RECT 1813.510 2.400 1818.190 2.680 ;
        RECT 1819.030 2.400 1823.710 2.680 ;
        RECT 1824.550 2.400 1829.230 2.680 ;
        RECT 1830.070 2.400 1834.750 2.680 ;
        RECT 1835.590 2.400 1839.810 2.680 ;
        RECT 1840.650 2.400 1845.330 2.680 ;
        RECT 1846.170 2.400 1850.850 2.680 ;
        RECT 1851.690 2.400 1856.370 2.680 ;
        RECT 1857.210 2.400 1861.430 2.680 ;
        RECT 1862.270 2.400 1866.950 2.680 ;
        RECT 1867.790 2.400 1872.470 2.680 ;
        RECT 1873.310 2.400 1877.990 2.680 ;
        RECT 1878.830 2.400 1883.510 2.680 ;
        RECT 1884.350 2.400 1888.570 2.680 ;
        RECT 1889.410 2.400 1894.090 2.680 ;
        RECT 1894.930 2.400 1899.610 2.680 ;
        RECT 1900.450 2.400 1905.130 2.680 ;
        RECT 1905.970 2.400 1910.650 2.680 ;
        RECT 1911.490 2.400 1915.710 2.680 ;
        RECT 1916.550 2.400 1921.230 2.680 ;
        RECT 1922.070 2.400 1926.750 2.680 ;
        RECT 1927.590 2.400 1932.270 2.680 ;
        RECT 1933.110 2.400 1937.790 2.680 ;
        RECT 1938.630 2.400 1942.850 2.680 ;
        RECT 1943.690 2.400 1948.370 2.680 ;
        RECT 1949.210 2.400 1953.890 2.680 ;
        RECT 1954.730 2.400 1959.410 2.680 ;
        RECT 1960.250 2.400 1964.470 2.680 ;
        RECT 1965.310 2.400 1969.990 2.680 ;
        RECT 1970.830 2.400 1975.510 2.680 ;
        RECT 1976.350 2.400 1981.030 2.680 ;
        RECT 1981.870 2.400 1986.550 2.680 ;
        RECT 1987.390 2.400 1991.610 2.680 ;
        RECT 1992.450 2.400 1997.130 2.680 ;
        RECT 1997.970 2.400 2002.650 2.680 ;
        RECT 2003.490 2.400 2008.170 2.680 ;
        RECT 2009.010 2.400 2013.690 2.680 ;
        RECT 2014.530 2.400 2018.750 2.680 ;
        RECT 2019.590 2.400 2024.270 2.680 ;
        RECT 2025.110 2.400 2029.790 2.680 ;
        RECT 2030.630 2.400 2035.310 2.680 ;
        RECT 2036.150 2.400 2040.370 2.680 ;
        RECT 2041.210 2.400 2045.890 2.680 ;
        RECT 2046.730 2.400 2051.410 2.680 ;
        RECT 2052.250 2.400 2056.930 2.680 ;
        RECT 2057.770 2.400 2062.450 2.680 ;
        RECT 2063.290 2.400 2067.510 2.680 ;
        RECT 2068.350 2.400 2073.030 2.680 ;
        RECT 2073.870 2.400 2078.550 2.680 ;
        RECT 2079.390 2.400 2084.070 2.680 ;
        RECT 2084.910 2.400 2089.590 2.680 ;
        RECT 2090.430 2.400 2094.650 2.680 ;
        RECT 2095.490 2.400 2100.170 2.680 ;
        RECT 2101.010 2.400 2105.690 2.680 ;
        RECT 2106.530 2.400 2111.210 2.680 ;
        RECT 2112.050 2.400 2116.270 2.680 ;
        RECT 2117.110 2.400 2121.790 2.680 ;
        RECT 2122.630 2.400 2127.310 2.680 ;
        RECT 2128.150 2.400 2132.830 2.680 ;
        RECT 2133.670 2.400 2138.350 2.680 ;
        RECT 2139.190 2.400 2143.410 2.680 ;
        RECT 2144.250 2.400 2148.930 2.680 ;
        RECT 2149.770 2.400 2154.450 2.680 ;
        RECT 2155.290 2.400 2159.970 2.680 ;
        RECT 2160.810 2.400 2165.490 2.680 ;
        RECT 2166.330 2.400 2170.550 2.680 ;
        RECT 2171.390 2.400 2176.070 2.680 ;
        RECT 2176.910 2.400 2181.590 2.680 ;
        RECT 2182.430 2.400 2187.110 2.680 ;
        RECT 2187.950 2.400 2192.630 2.680 ;
        RECT 2193.470 2.400 2197.690 2.680 ;
        RECT 2198.530 2.400 2203.210 2.680 ;
        RECT 2204.050 2.400 2208.730 2.680 ;
        RECT 2209.570 2.400 2214.250 2.680 ;
        RECT 2215.090 2.400 2219.310 2.680 ;
        RECT 2220.150 2.400 2224.830 2.680 ;
        RECT 2225.670 2.400 2230.350 2.680 ;
        RECT 2231.190 2.400 2235.870 2.680 ;
        RECT 2236.710 2.400 2241.390 2.680 ;
        RECT 2242.230 2.400 2246.450 2.680 ;
        RECT 2247.290 2.400 2251.970 2.680 ;
        RECT 2252.810 2.400 2257.490 2.680 ;
        RECT 2258.330 2.400 2263.010 2.680 ;
        RECT 2263.850 2.400 2268.530 2.680 ;
        RECT 2269.370 2.400 2273.590 2.680 ;
        RECT 2274.430 2.400 2279.110 2.680 ;
        RECT 2279.950 2.400 2284.630 2.680 ;
        RECT 2285.470 2.400 2290.150 2.680 ;
        RECT 2290.990 2.400 2295.210 2.680 ;
        RECT 2296.050 2.400 2300.730 2.680 ;
        RECT 2301.570 2.400 2306.250 2.680 ;
        RECT 2307.090 2.400 2311.770 2.680 ;
        RECT 2312.610 2.400 2317.290 2.680 ;
        RECT 2318.130 2.400 2322.350 2.680 ;
        RECT 2323.190 2.400 2327.870 2.680 ;
        RECT 2328.710 2.400 2333.390 2.680 ;
        RECT 2334.230 2.400 2338.910 2.680 ;
        RECT 2339.750 2.400 2344.430 2.680 ;
        RECT 2345.270 2.400 2349.490 2.680 ;
        RECT 2350.330 2.400 2355.010 2.680 ;
        RECT 2355.850 2.400 2360.530 2.680 ;
        RECT 2361.370 2.400 2366.050 2.680 ;
        RECT 2366.890 2.400 2371.110 2.680 ;
        RECT 2371.950 2.400 2376.630 2.680 ;
        RECT 2377.470 2.400 2382.150 2.680 ;
        RECT 2382.990 2.400 2387.670 2.680 ;
        RECT 2388.510 2.400 2393.190 2.680 ;
        RECT 2394.030 2.400 2398.250 2.680 ;
        RECT 2399.090 2.400 2403.770 2.680 ;
        RECT 2404.610 2.400 2409.290 2.680 ;
        RECT 2410.130 2.400 2414.810 2.680 ;
        RECT 2415.650 2.400 2420.330 2.680 ;
        RECT 2421.170 2.400 2425.390 2.680 ;
        RECT 2426.230 2.400 2430.910 2.680 ;
        RECT 2431.750 2.400 2436.430 2.680 ;
        RECT 2437.270 2.400 2441.950 2.680 ;
        RECT 2442.790 2.400 2447.470 2.680 ;
        RECT 2448.310 2.400 2452.530 2.680 ;
        RECT 2453.370 2.400 2458.050 2.680 ;
        RECT 2458.890 2.400 2463.570 2.680 ;
        RECT 2464.410 2.400 2469.090 2.680 ;
        RECT 2469.930 2.400 2474.150 2.680 ;
        RECT 2474.990 2.400 2479.670 2.680 ;
        RECT 2480.510 2.400 2485.190 2.680 ;
        RECT 2486.030 2.400 2490.710 2.680 ;
        RECT 2491.550 2.400 2496.230 2.680 ;
        RECT 2497.070 2.400 2501.290 2.680 ;
        RECT 2502.130 2.400 2506.810 2.680 ;
        RECT 2507.650 2.400 2512.330 2.680 ;
        RECT 2513.170 2.400 2517.850 2.680 ;
        RECT 2518.690 2.400 2523.370 2.680 ;
        RECT 2524.210 2.400 2528.430 2.680 ;
        RECT 2529.270 2.400 2533.950 2.680 ;
        RECT 2534.790 2.400 2539.470 2.680 ;
        RECT 2540.310 2.400 2544.990 2.680 ;
        RECT 2545.830 2.400 2550.050 2.680 ;
        RECT 2550.890 2.400 2555.570 2.680 ;
        RECT 2556.410 2.400 2561.090 2.680 ;
        RECT 2561.930 2.400 2566.610 2.680 ;
        RECT 2567.450 2.400 2572.130 2.680 ;
        RECT 2572.970 2.400 2577.190 2.680 ;
        RECT 2578.030 2.400 2582.710 2.680 ;
        RECT 2583.550 2.400 2588.230 2.680 ;
        RECT 2589.070 2.400 2593.750 2.680 ;
        RECT 2594.590 2.400 2599.270 2.680 ;
        RECT 2600.110 2.400 2604.330 2.680 ;
        RECT 2605.170 2.400 2609.850 2.680 ;
        RECT 2610.690 2.400 2615.370 2.680 ;
        RECT 2616.210 2.400 2620.890 2.680 ;
        RECT 2621.730 2.400 2625.950 2.680 ;
        RECT 2626.790 2.400 2631.470 2.680 ;
        RECT 2632.310 2.400 2636.990 2.680 ;
        RECT 2637.830 2.400 2642.510 2.680 ;
        RECT 2643.350 2.400 2648.030 2.680 ;
        RECT 2648.870 2.400 2653.090 2.680 ;
        RECT 2653.930 2.400 2658.610 2.680 ;
        RECT 2659.450 2.400 2664.130 2.680 ;
        RECT 2664.970 2.400 2669.650 2.680 ;
        RECT 2670.490 2.400 2675.170 2.680 ;
        RECT 2676.010 2.400 2680.230 2.680 ;
        RECT 2681.070 2.400 2685.750 2.680 ;
        RECT 2686.590 2.400 2689.070 2.680 ;
      LAYER met3 ;
        RECT 2.400 3666.920 2697.600 3688.485 ;
        RECT 2.800 3665.520 2697.200 3666.920 ;
        RECT 2.400 3599.600 2697.600 3665.520 ;
        RECT 2.800 3598.200 2697.200 3599.600 ;
        RECT 2.400 3532.280 2697.600 3598.200 ;
        RECT 2.800 3530.880 2697.200 3532.280 ;
        RECT 2.400 3464.960 2697.600 3530.880 ;
        RECT 2.800 3463.560 2697.200 3464.960 ;
        RECT 2.400 3397.640 2697.600 3463.560 ;
        RECT 2.800 3396.240 2697.200 3397.640 ;
        RECT 2.400 3330.320 2697.600 3396.240 ;
        RECT 2.800 3328.920 2697.200 3330.320 ;
        RECT 2.400 3263.000 2697.600 3328.920 ;
        RECT 2.800 3261.600 2697.200 3263.000 ;
        RECT 2.400 3195.680 2697.600 3261.600 ;
        RECT 2.800 3194.280 2697.200 3195.680 ;
        RECT 2.400 3128.360 2697.600 3194.280 ;
        RECT 2.800 3126.960 2697.200 3128.360 ;
        RECT 2.400 3061.040 2697.600 3126.960 ;
        RECT 2.800 3059.640 2697.200 3061.040 ;
        RECT 2.400 2993.720 2697.600 3059.640 ;
        RECT 2.800 2992.320 2697.200 2993.720 ;
        RECT 2.400 2926.400 2697.600 2992.320 ;
        RECT 2.800 2925.000 2697.200 2926.400 ;
        RECT 2.400 2859.080 2697.600 2925.000 ;
        RECT 2.800 2857.680 2697.200 2859.080 ;
        RECT 2.400 2792.440 2697.600 2857.680 ;
        RECT 2.800 2791.040 2697.200 2792.440 ;
        RECT 2.400 2725.120 2697.600 2791.040 ;
        RECT 2.800 2723.720 2697.200 2725.120 ;
        RECT 2.400 2657.800 2697.600 2723.720 ;
        RECT 2.800 2656.400 2697.200 2657.800 ;
        RECT 2.400 2590.480 2697.600 2656.400 ;
        RECT 2.800 2589.080 2697.200 2590.480 ;
        RECT 2.400 2523.160 2697.600 2589.080 ;
        RECT 2.800 2521.760 2697.200 2523.160 ;
        RECT 2.400 2455.840 2697.600 2521.760 ;
        RECT 2.800 2454.440 2697.200 2455.840 ;
        RECT 2.400 2388.520 2697.600 2454.440 ;
        RECT 2.800 2387.120 2697.200 2388.520 ;
        RECT 2.400 2321.200 2697.600 2387.120 ;
        RECT 2.800 2319.800 2697.200 2321.200 ;
        RECT 2.400 2253.880 2697.600 2319.800 ;
        RECT 2.800 2252.480 2697.200 2253.880 ;
        RECT 2.400 2186.560 2697.600 2252.480 ;
        RECT 2.800 2185.160 2697.200 2186.560 ;
        RECT 2.400 2119.240 2697.600 2185.160 ;
        RECT 2.800 2117.840 2697.200 2119.240 ;
        RECT 2.400 2051.920 2697.600 2117.840 ;
        RECT 2.800 2050.520 2697.200 2051.920 ;
        RECT 2.400 1984.600 2697.600 2050.520 ;
        RECT 2.800 1983.200 2697.200 1984.600 ;
        RECT 2.400 1917.280 2697.600 1983.200 ;
        RECT 2.800 1915.880 2697.200 1917.280 ;
        RECT 2.400 1850.640 2697.600 1915.880 ;
        RECT 2.800 1849.240 2697.200 1850.640 ;
        RECT 2.400 1783.320 2697.600 1849.240 ;
        RECT 2.800 1781.920 2697.200 1783.320 ;
        RECT 2.400 1716.000 2697.600 1781.920 ;
        RECT 2.800 1714.600 2697.200 1716.000 ;
        RECT 2.400 1648.680 2697.600 1714.600 ;
        RECT 2.800 1647.280 2697.200 1648.680 ;
        RECT 2.400 1581.360 2697.600 1647.280 ;
        RECT 2.800 1579.960 2697.200 1581.360 ;
        RECT 2.400 1514.040 2697.600 1579.960 ;
        RECT 2.800 1512.640 2697.200 1514.040 ;
        RECT 2.400 1446.720 2697.600 1512.640 ;
        RECT 2.800 1445.320 2697.200 1446.720 ;
        RECT 2.400 1379.400 2697.600 1445.320 ;
        RECT 2.800 1378.000 2697.200 1379.400 ;
        RECT 2.400 1312.080 2697.600 1378.000 ;
        RECT 2.800 1310.680 2697.200 1312.080 ;
        RECT 2.400 1244.760 2697.600 1310.680 ;
        RECT 2.800 1243.360 2697.200 1244.760 ;
        RECT 2.400 1177.440 2697.600 1243.360 ;
        RECT 2.800 1176.040 2697.200 1177.440 ;
        RECT 2.400 1110.120 2697.600 1176.040 ;
        RECT 2.800 1108.720 2697.200 1110.120 ;
        RECT 2.400 1042.800 2697.600 1108.720 ;
        RECT 2.800 1041.400 2697.200 1042.800 ;
        RECT 2.400 975.480 2697.600 1041.400 ;
        RECT 2.800 974.080 2697.200 975.480 ;
        RECT 2.400 908.840 2697.600 974.080 ;
        RECT 2.800 907.440 2697.200 908.840 ;
        RECT 2.400 841.520 2697.600 907.440 ;
        RECT 2.800 840.120 2697.200 841.520 ;
        RECT 2.400 774.200 2697.600 840.120 ;
        RECT 2.800 772.800 2697.200 774.200 ;
        RECT 2.400 706.880 2697.600 772.800 ;
        RECT 2.800 705.480 2697.200 706.880 ;
        RECT 2.400 639.560 2697.600 705.480 ;
        RECT 2.800 638.160 2697.200 639.560 ;
        RECT 2.400 572.240 2697.600 638.160 ;
        RECT 2.800 570.840 2697.200 572.240 ;
        RECT 2.400 504.920 2697.600 570.840 ;
        RECT 2.800 503.520 2697.200 504.920 ;
        RECT 2.400 437.600 2697.600 503.520 ;
        RECT 2.800 436.200 2697.200 437.600 ;
        RECT 2.400 370.280 2697.600 436.200 ;
        RECT 2.800 368.880 2697.200 370.280 ;
        RECT 2.400 302.960 2697.600 368.880 ;
        RECT 2.800 301.560 2697.200 302.960 ;
        RECT 2.400 235.640 2697.600 301.560 ;
        RECT 2.800 234.240 2697.200 235.640 ;
        RECT 2.400 168.320 2697.600 234.240 ;
        RECT 2.800 166.920 2697.200 168.320 ;
        RECT 2.400 101.000 2697.600 166.920 ;
        RECT 2.800 99.600 2697.200 101.000 ;
        RECT 2.400 34.360 2697.600 99.600 ;
        RECT 2.800 32.960 2697.200 34.360 ;
        RECT 2.400 10.715 2697.600 32.960 ;
      LAYER met4 ;
        RECT 16.855 10.640 2633.840 3688.560 ;
      LAYER met5 ;
        RECT 5.520 179.670 2694.220 3627.820 ;
  END
END user_project_wrapper
END LIBRARY

