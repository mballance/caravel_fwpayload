VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN -0.005 0.000 ;
  SIZE 1097.885 BY 1100.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 3.710 1096.000 3.990 1100.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 293.050 1096.000 293.330 1100.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.030 1096.000 322.310 1100.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 351.010 1096.000 351.290 1100.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 379.530 1096.000 379.810 1100.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.510 1096.000 408.790 1100.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 437.490 1096.000 437.770 1100.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 466.470 1096.000 466.750 1100.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 495.450 1096.000 495.730 1100.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 524.430 1096.000 524.710 1100.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 553.410 1096.000 553.690 1100.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 32.230 1096.000 32.510 1100.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 582.390 1096.000 582.670 1100.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 611.370 1096.000 611.650 1100.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 640.350 1096.000 640.630 1100.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 669.330 1096.000 669.610 1100.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.310 1096.000 698.590 1100.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 727.290 1096.000 727.570 1100.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 755.810 1096.000 756.090 1100.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 784.790 1096.000 785.070 1100.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 813.770 1096.000 814.050 1100.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 842.750 1096.000 843.030 1100.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.210 1096.000 61.490 1100.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 871.730 1096.000 872.010 1100.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 900.710 1096.000 900.990 1100.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.690 1096.000 929.970 1100.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 958.670 1096.000 958.950 1100.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 987.650 1096.000 987.930 1100.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1016.630 1096.000 1016.910 1100.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1045.610 1096.000 1045.890 1100.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1074.590 1096.000 1074.870 1100.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 90.190 1096.000 90.470 1100.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.170 1096.000 119.450 1100.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.150 1096.000 148.430 1100.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 177.130 1096.000 177.410 1100.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.110 1096.000 206.390 1100.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 235.090 1096.000 235.370 1100.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.070 1096.000 264.350 1100.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 12.910 1096.000 13.190 1100.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 302.710 1096.000 302.990 1100.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 331.690 1096.000 331.970 1100.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 360.670 1096.000 360.950 1100.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 389.190 1096.000 389.470 1100.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 418.170 1096.000 418.450 1100.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 447.150 1096.000 447.430 1100.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 476.130 1096.000 476.410 1100.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 505.110 1096.000 505.390 1100.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 534.090 1096.000 534.370 1100.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 563.070 1096.000 563.350 1100.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.890 1096.000 42.170 1100.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 592.050 1096.000 592.330 1100.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 621.030 1096.000 621.310 1100.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 650.010 1096.000 650.290 1100.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 678.990 1096.000 679.270 1100.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 707.970 1096.000 708.250 1100.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 736.950 1096.000 737.230 1100.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 765.470 1096.000 765.750 1100.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 794.450 1096.000 794.730 1100.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 823.430 1096.000 823.710 1100.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.410 1096.000 852.690 1100.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 70.870 1096.000 71.150 1100.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 881.390 1096.000 881.670 1100.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 910.370 1096.000 910.650 1100.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 939.350 1096.000 939.630 1100.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 968.330 1096.000 968.610 1100.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 997.310 1096.000 997.590 1100.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1026.290 1096.000 1026.570 1100.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1055.270 1096.000 1055.550 1100.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1084.250 1096.000 1084.530 1100.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 99.850 1096.000 100.130 1100.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.830 1096.000 129.110 1100.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 157.810 1096.000 158.090 1100.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 186.790 1096.000 187.070 1100.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 215.770 1096.000 216.050 1100.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 244.750 1096.000 245.030 1100.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 273.730 1096.000 274.010 1100.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 22.570 1096.000 22.850 1100.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 312.370 1096.000 312.650 1100.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 341.350 1096.000 341.630 1100.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 370.330 1096.000 370.610 1100.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 398.850 1096.000 399.130 1100.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 427.830 1096.000 428.110 1100.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 456.810 1096.000 457.090 1100.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 485.790 1096.000 486.070 1100.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 514.770 1096.000 515.050 1100.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 543.750 1096.000 544.030 1100.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 572.730 1096.000 573.010 1100.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 51.550 1096.000 51.830 1100.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 601.710 1096.000 601.990 1100.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 630.690 1096.000 630.970 1100.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 659.670 1096.000 659.950 1100.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 688.650 1096.000 688.930 1100.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 717.630 1096.000 717.910 1100.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 746.150 1096.000 746.430 1100.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 775.130 1096.000 775.410 1100.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 804.110 1096.000 804.390 1100.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 833.090 1096.000 833.370 1100.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 862.070 1096.000 862.350 1100.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.530 1096.000 80.810 1100.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 891.050 1096.000 891.330 1100.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 920.030 1096.000 920.310 1100.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 949.010 1096.000 949.290 1100.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 977.990 1096.000 978.270 1100.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1006.970 1096.000 1007.250 1100.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1035.950 1096.000 1036.230 1100.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1064.930 1096.000 1065.210 1100.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1093.910 1096.000 1094.190 1100.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.510 1096.000 109.790 1100.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.490 1096.000 138.770 1100.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.470 1096.000 167.750 1100.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.450 1096.000 196.730 1100.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 225.430 1096.000 225.710 1100.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 254.410 1096.000 254.690 1100.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 283.390 1096.000 283.670 1100.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 237.850 0.000 238.130 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 911.290 0.000 911.570 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 917.730 0.000 918.010 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 924.630 0.000 924.910 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 931.530 0.000 931.810 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 937.970 0.000 938.250 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 944.870 0.000 945.150 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 951.310 0.000 951.590 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 958.210 0.000 958.490 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.110 0.000 965.390 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 971.550 0.000 971.830 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 305.010 0.000 305.290 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 978.450 0.000 978.730 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 985.350 0.000 985.630 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 991.790 0.000 992.070 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 998.690 0.000 998.970 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1005.590 0.000 1005.870 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1012.030 0.000 1012.310 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1018.930 0.000 1019.210 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1025.370 0.000 1025.650 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.270 0.000 1032.550 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1039.170 0.000 1039.450 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.910 0.000 312.190 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1045.610 0.000 1045.890 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1052.510 0.000 1052.790 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1059.410 0.000 1059.690 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1065.850 0.000 1066.130 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1072.750 0.000 1073.030 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.650 0.000 1079.930 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1086.090 0.000 1086.370 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1092.990 0.000 1093.270 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 318.350 0.000 318.630 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 325.250 0.000 325.530 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 332.150 0.000 332.430 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 338.590 0.000 338.870 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 345.490 0.000 345.770 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 352.390 0.000 352.670 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 358.830 0.000 359.110 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.730 0.000 366.010 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 244.290 0.000 244.570 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 372.630 0.000 372.910 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 379.070 0.000 379.350 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 385.970 0.000 386.250 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.410 0.000 392.690 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 399.310 0.000 399.590 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 406.210 0.000 406.490 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 412.650 0.000 412.930 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 419.550 0.000 419.830 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.450 0.000 426.730 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.890 0.000 433.170 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 251.190 0.000 251.470 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 439.790 0.000 440.070 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 446.690 0.000 446.970 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 453.130 0.000 453.410 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.030 0.000 460.310 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 466.470 0.000 466.750 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 473.370 0.000 473.650 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 480.270 0.000 480.550 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 486.710 0.000 486.990 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 493.610 0.000 493.890 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 500.510 0.000 500.790 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.090 0.000 258.370 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 506.950 0.000 507.230 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 513.850 0.000 514.130 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 520.750 0.000 521.030 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.190 0.000 527.470 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 534.090 0.000 534.370 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 540.530 0.000 540.810 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 547.430 0.000 547.710 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 554.330 0.000 554.610 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 560.770 0.000 561.050 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 567.670 0.000 567.950 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.530 0.000 264.810 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 574.570 0.000 574.850 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 581.010 0.000 581.290 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.910 0.000 588.190 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 594.810 0.000 595.090 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 601.250 0.000 601.530 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 608.150 0.000 608.430 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 615.050 0.000 615.330 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 621.490 0.000 621.770 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 628.390 0.000 628.670 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 634.830 0.000 635.110 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 271.430 0.000 271.710 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 641.730 0.000 642.010 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 648.630 0.000 648.910 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 655.070 0.000 655.350 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 661.970 0.000 662.250 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 668.870 0.000 669.150 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 675.310 0.000 675.590 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 682.210 0.000 682.490 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 689.110 0.000 689.390 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 695.550 0.000 695.830 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 702.450 0.000 702.730 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 278.330 0.000 278.610 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 708.890 0.000 709.170 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 715.790 0.000 716.070 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.690 0.000 722.970 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 729.130 0.000 729.410 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 736.030 0.000 736.310 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 742.930 0.000 743.210 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 749.370 0.000 749.650 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 756.270 0.000 756.550 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 763.170 0.000 763.450 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 769.610 0.000 769.890 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 284.770 0.000 285.050 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 776.510 0.000 776.790 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 782.950 0.000 783.230 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 789.850 0.000 790.130 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 796.750 0.000 797.030 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 803.190 0.000 803.470 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 810.090 0.000 810.370 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 816.990 0.000 817.270 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 823.430 0.000 823.710 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 830.330 0.000 830.610 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 837.230 0.000 837.510 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 291.670 0.000 291.950 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 843.670 0.000 843.950 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 850.570 0.000 850.850 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 857.470 0.000 857.750 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 863.910 0.000 864.190 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 870.810 0.000 871.090 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 877.250 0.000 877.530 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 884.150 0.000 884.430 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 891.050 0.000 891.330 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 897.490 0.000 897.770 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 904.390 0.000 904.670 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 298.110 0.000 298.390 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 240.150 0.000 240.430 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 913.130 0.000 913.410 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 920.030 0.000 920.310 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 926.930 0.000 927.210 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 933.370 0.000 933.650 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 940.270 0.000 940.550 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 947.170 0.000 947.450 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 953.610 0.000 953.890 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 960.510 0.000 960.790 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 967.410 0.000 967.690 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 973.850 0.000 974.130 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 307.310 0.000 307.590 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 980.750 0.000 981.030 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 987.650 0.000 987.930 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 994.090 0.000 994.370 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1000.990 0.000 1001.270 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1007.430 0.000 1007.710 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1014.330 0.000 1014.610 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1021.230 0.000 1021.510 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1027.670 0.000 1027.950 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1034.570 0.000 1034.850 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1041.470 0.000 1041.750 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 314.210 0.000 314.490 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1047.910 0.000 1048.190 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1054.810 0.000 1055.090 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1061.710 0.000 1061.990 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1068.150 0.000 1068.430 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1075.050 0.000 1075.330 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1081.490 0.000 1081.770 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1088.390 0.000 1088.670 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1095.290 0.000 1095.570 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 320.650 0.000 320.930 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 327.550 0.000 327.830 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 334.450 0.000 334.730 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 340.890 0.000 341.170 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.790 0.000 348.070 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.230 0.000 354.510 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 361.130 0.000 361.410 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.030 0.000 368.310 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 246.590 0.000 246.870 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 374.470 0.000 374.750 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 381.370 0.000 381.650 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 388.270 0.000 388.550 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 394.710 0.000 394.990 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 401.610 0.000 401.890 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 408.510 0.000 408.790 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 414.950 0.000 415.230 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 421.850 0.000 422.130 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 428.750 0.000 429.030 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 435.190 0.000 435.470 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 253.490 0.000 253.770 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 442.090 0.000 442.370 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.530 0.000 448.810 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 455.430 0.000 455.710 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 462.330 0.000 462.610 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 468.770 0.000 469.050 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 475.670 0.000 475.950 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 482.570 0.000 482.850 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.010 0.000 489.290 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 495.910 0.000 496.190 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.810 0.000 503.090 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 260.390 0.000 260.670 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 509.250 0.000 509.530 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 516.150 0.000 516.430 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 522.590 0.000 522.870 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 529.490 0.000 529.770 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 536.390 0.000 536.670 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 542.830 0.000 543.110 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 549.730 0.000 550.010 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 556.630 0.000 556.910 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 563.070 0.000 563.350 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 569.970 0.000 570.250 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 266.830 0.000 267.110 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 576.870 0.000 577.150 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 583.310 0.000 583.590 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 590.210 0.000 590.490 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 596.650 0.000 596.930 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 603.550 0.000 603.830 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 610.450 0.000 610.730 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 616.890 0.000 617.170 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 623.790 0.000 624.070 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 630.690 0.000 630.970 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 637.130 0.000 637.410 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 273.730 0.000 274.010 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 644.030 0.000 644.310 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 650.930 0.000 651.210 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 657.370 0.000 657.650 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 664.270 0.000 664.550 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 670.710 0.000 670.990 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 677.610 0.000 677.890 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 684.510 0.000 684.790 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 690.950 0.000 691.230 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 697.850 0.000 698.130 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 704.750 0.000 705.030 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 280.170 0.000 280.450 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 711.190 0.000 711.470 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 718.090 0.000 718.370 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 724.990 0.000 725.270 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 731.430 0.000 731.710 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 738.330 0.000 738.610 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 745.230 0.000 745.510 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 751.670 0.000 751.950 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 758.570 0.000 758.850 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 765.010 0.000 765.290 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 771.910 0.000 772.190 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.070 0.000 287.350 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 778.810 0.000 779.090 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 785.250 0.000 785.530 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 792.150 0.000 792.430 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 799.050 0.000 799.330 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 805.490 0.000 805.770 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 812.390 0.000 812.670 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 819.290 0.000 819.570 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 825.730 0.000 826.010 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 832.630 0.000 832.910 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 839.070 0.000 839.350 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 293.970 0.000 294.250 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 845.970 0.000 846.250 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.870 0.000 853.150 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 859.310 0.000 859.590 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 866.210 0.000 866.490 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 873.110 0.000 873.390 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 879.550 0.000 879.830 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 886.450 0.000 886.730 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 893.350 0.000 893.630 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 899.790 0.000 900.070 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 906.690 0.000 906.970 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 300.410 0.000 300.690 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 241.990 0.000 242.270 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 915.430 0.000 915.710 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 922.330 0.000 922.610 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.230 0.000 929.510 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 935.670 0.000 935.950 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 942.570 0.000 942.850 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 949.470 0.000 949.750 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 955.910 0.000 956.190 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 962.810 0.000 963.090 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 969.250 0.000 969.530 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 976.150 0.000 976.430 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 309.610 0.000 309.890 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 983.050 0.000 983.330 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 989.490 0.000 989.770 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 996.390 0.000 996.670 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1003.290 0.000 1003.570 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1009.730 0.000 1010.010 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1016.630 0.000 1016.910 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1023.530 0.000 1023.810 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1029.970 0.000 1030.250 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1036.870 0.000 1037.150 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1043.770 0.000 1044.050 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.510 0.000 316.790 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1050.210 0.000 1050.490 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1057.110 0.000 1057.390 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1063.550 0.000 1063.830 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1070.450 0.000 1070.730 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1077.350 0.000 1077.630 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.790 0.000 1084.070 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1090.690 0.000 1090.970 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1097.590 0.000 1097.870 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.950 0.000 323.230 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.850 0.000 330.130 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 336.290 0.000 336.570 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 343.190 0.000 343.470 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 350.090 0.000 350.370 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 356.530 0.000 356.810 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 363.430 0.000 363.710 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 370.330 0.000 370.610 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 248.890 0.000 249.170 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 376.770 0.000 377.050 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.670 0.000 383.950 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.570 0.000 390.850 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 397.010 0.000 397.290 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 403.910 0.000 404.190 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 410.350 0.000 410.630 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 417.250 0.000 417.530 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 424.150 0.000 424.430 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 430.590 0.000 430.870 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 437.490 0.000 437.770 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 255.790 0.000 256.070 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 444.390 0.000 444.670 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 450.830 0.000 451.110 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 457.730 0.000 458.010 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 464.630 0.000 464.910 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 471.070 0.000 471.350 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 477.970 0.000 478.250 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 484.410 0.000 484.690 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 491.310 0.000 491.590 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 498.210 0.000 498.490 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 504.650 0.000 504.930 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 262.230 0.000 262.510 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 511.550 0.000 511.830 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 518.450 0.000 518.730 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 524.890 0.000 525.170 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.790 0.000 532.070 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 538.690 0.000 538.970 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 545.130 0.000 545.410 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 552.030 0.000 552.310 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 558.930 0.000 559.210 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 565.370 0.000 565.650 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 572.270 0.000 572.550 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 269.130 0.000 269.410 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 578.710 0.000 578.990 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 585.610 0.000 585.890 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 592.510 0.000 592.790 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 598.950 0.000 599.230 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 605.850 0.000 606.130 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 612.750 0.000 613.030 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 619.190 0.000 619.470 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 626.090 0.000 626.370 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 632.990 0.000 633.270 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 639.430 0.000 639.710 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 276.030 0.000 276.310 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 646.330 0.000 646.610 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 652.770 0.000 653.050 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 659.670 0.000 659.950 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 666.570 0.000 666.850 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 673.010 0.000 673.290 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 679.910 0.000 680.190 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 686.810 0.000 687.090 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 693.250 0.000 693.530 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 700.150 0.000 700.430 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 707.050 0.000 707.330 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.470 0.000 282.750 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 713.490 0.000 713.770 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 720.390 0.000 720.670 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 726.830 0.000 727.110 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 733.730 0.000 734.010 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 740.630 0.000 740.910 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 747.070 0.000 747.350 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 753.970 0.000 754.250 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 760.870 0.000 761.150 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 767.310 0.000 767.590 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 774.210 0.000 774.490 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 289.370 0.000 289.650 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 781.110 0.000 781.390 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 787.550 0.000 787.830 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 794.450 0.000 794.730 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 801.350 0.000 801.630 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 807.790 0.000 808.070 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 814.690 0.000 814.970 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 821.130 0.000 821.410 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 828.030 0.000 828.310 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 834.930 0.000 835.210 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 841.370 0.000 841.650 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 296.270 0.000 296.550 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 848.270 0.000 848.550 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 855.170 0.000 855.450 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 861.610 0.000 861.890 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 868.510 0.000 868.790 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 875.410 0.000 875.690 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 881.850 0.000 882.130 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 888.750 0.000 889.030 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 895.190 0.000 895.470 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 902.090 0.000 902.370 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 908.990 0.000 909.270 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.710 0.000 302.990 4.000 ;
    END
  END la_oen[9]
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 0.030 0.000 0.310 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.870 0.000 2.150 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.170 0.000 4.450 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.370 0.000 13.650 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.730 0.000 90.010 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.170 0.000 96.450 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.070 0.000 103.350 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.970 0.000 110.250 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.410 0.000 116.690 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.310 0.000 123.590 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.210 0.000 130.490 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 136.650 0.000 136.930 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 143.550 0.000 143.830 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 149.990 0.000 150.270 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.110 0.000 22.390 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 156.890 0.000 157.170 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 163.790 0.000 164.070 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.230 0.000 170.510 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 177.130 0.000 177.410 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.030 0.000 184.310 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.470 0.000 190.750 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 197.370 0.000 197.650 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 204.270 0.000 204.550 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 210.710 0.000 210.990 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 217.610 0.000 217.890 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.310 0.000 31.590 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.050 0.000 224.330 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 230.950 0.000 231.230 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.050 0.000 40.330 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 49.250 0.000 49.530 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.690 0.000 55.970 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.590 0.000 62.870 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 69.490 0.000 69.770 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 75.930 0.000 76.210 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 82.830 0.000 83.110 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.470 0.000 6.750 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 15.670 0.000 15.950 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.030 0.000 92.310 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.470 0.000 98.750 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.370 0.000 105.650 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 111.810 0.000 112.090 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.710 0.000 118.990 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 125.610 0.000 125.890 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 132.050 0.000 132.330 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 138.950 0.000 139.230 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 145.850 0.000 146.130 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 152.290 0.000 152.570 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 24.410 0.000 24.690 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.190 0.000 159.470 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.090 0.000 166.370 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.530 0.000 172.810 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 179.430 0.000 179.710 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 186.330 0.000 186.610 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 192.770 0.000 193.050 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 199.670 0.000 199.950 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.110 0.000 206.390 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 213.010 0.000 213.290 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 219.910 0.000 220.190 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 33.610 0.000 33.890 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 226.350 0.000 226.630 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 233.250 0.000 233.530 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 42.350 0.000 42.630 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 51.550 0.000 51.830 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.990 0.000 58.270 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 64.890 0.000 65.170 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.790 0.000 72.070 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 78.230 0.000 78.510 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 85.130 0.000 85.410 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 17.970 0.000 18.250 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.870 0.000 94.150 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 100.770 0.000 101.050 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.670 0.000 107.950 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 114.110 0.000 114.390 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 121.010 0.000 121.290 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 127.910 0.000 128.190 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 134.350 0.000 134.630 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 141.250 0.000 141.530 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 148.150 0.000 148.430 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 154.590 0.000 154.870 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 26.710 0.000 26.990 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 161.490 0.000 161.770 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.930 0.000 168.210 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.830 0.000 175.110 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 181.730 0.000 182.010 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 188.170 0.000 188.450 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 195.070 0.000 195.350 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 201.970 0.000 202.250 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 208.410 0.000 208.690 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 215.310 0.000 215.590 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.210 0.000 222.490 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 35.910 0.000 36.190 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 228.650 0.000 228.930 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 235.550 0.000 235.830 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 44.650 0.000 44.930 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 53.850 0.000 54.130 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 60.290 0.000 60.570 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.190 0.000 67.470 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.090 0.000 74.370 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.530 0.000 80.810 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.430 0.000 87.710 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.810 0.000 20.090 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 29.010 0.000 29.290 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 37.750 0.000 38.030 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.950 0.000 47.230 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 8.770 0.000 9.050 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 11.070 0.000 11.350 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.060 10.640 21.660 1088.240 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.860 10.640 98.460 1088.240 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 4.540 10.795 1093.360 1088.085 ;
      LAYER met1 ;
        RECT 4.150 7.860 1097.890 1096.120 ;
      LAYER met2 ;
        RECT 0.030 1095.720 3.430 1096.150 ;
        RECT 4.270 1095.720 12.630 1096.150 ;
        RECT 13.470 1095.720 22.290 1096.150 ;
        RECT 23.130 1095.720 31.950 1096.150 ;
        RECT 32.790 1095.720 41.610 1096.150 ;
        RECT 42.450 1095.720 51.270 1096.150 ;
        RECT 52.110 1095.720 60.930 1096.150 ;
        RECT 61.770 1095.720 70.590 1096.150 ;
        RECT 71.430 1095.720 80.250 1096.150 ;
        RECT 81.090 1095.720 89.910 1096.150 ;
        RECT 90.750 1095.720 99.570 1096.150 ;
        RECT 100.410 1095.720 109.230 1096.150 ;
        RECT 110.070 1095.720 118.890 1096.150 ;
        RECT 119.730 1095.720 128.550 1096.150 ;
        RECT 129.390 1095.720 138.210 1096.150 ;
        RECT 139.050 1095.720 147.870 1096.150 ;
        RECT 148.710 1095.720 157.530 1096.150 ;
        RECT 158.370 1095.720 167.190 1096.150 ;
        RECT 168.030 1095.720 176.850 1096.150 ;
        RECT 177.690 1095.720 186.510 1096.150 ;
        RECT 187.350 1095.720 196.170 1096.150 ;
        RECT 197.010 1095.720 205.830 1096.150 ;
        RECT 206.670 1095.720 215.490 1096.150 ;
        RECT 216.330 1095.720 225.150 1096.150 ;
        RECT 225.990 1095.720 234.810 1096.150 ;
        RECT 235.650 1095.720 244.470 1096.150 ;
        RECT 245.310 1095.720 254.130 1096.150 ;
        RECT 254.970 1095.720 263.790 1096.150 ;
        RECT 264.630 1095.720 273.450 1096.150 ;
        RECT 274.290 1095.720 283.110 1096.150 ;
        RECT 283.950 1095.720 292.770 1096.150 ;
        RECT 293.610 1095.720 302.430 1096.150 ;
        RECT 303.270 1095.720 312.090 1096.150 ;
        RECT 312.930 1095.720 321.750 1096.150 ;
        RECT 322.590 1095.720 331.410 1096.150 ;
        RECT 332.250 1095.720 341.070 1096.150 ;
        RECT 341.910 1095.720 350.730 1096.150 ;
        RECT 351.570 1095.720 360.390 1096.150 ;
        RECT 361.230 1095.720 370.050 1096.150 ;
        RECT 370.890 1095.720 379.250 1096.150 ;
        RECT 380.090 1095.720 388.910 1096.150 ;
        RECT 389.750 1095.720 398.570 1096.150 ;
        RECT 399.410 1095.720 408.230 1096.150 ;
        RECT 409.070 1095.720 417.890 1096.150 ;
        RECT 418.730 1095.720 427.550 1096.150 ;
        RECT 428.390 1095.720 437.210 1096.150 ;
        RECT 438.050 1095.720 446.870 1096.150 ;
        RECT 447.710 1095.720 456.530 1096.150 ;
        RECT 457.370 1095.720 466.190 1096.150 ;
        RECT 467.030 1095.720 475.850 1096.150 ;
        RECT 476.690 1095.720 485.510 1096.150 ;
        RECT 486.350 1095.720 495.170 1096.150 ;
        RECT 496.010 1095.720 504.830 1096.150 ;
        RECT 505.670 1095.720 514.490 1096.150 ;
        RECT 515.330 1095.720 524.150 1096.150 ;
        RECT 524.990 1095.720 533.810 1096.150 ;
        RECT 534.650 1095.720 543.470 1096.150 ;
        RECT 544.310 1095.720 553.130 1096.150 ;
        RECT 553.970 1095.720 562.790 1096.150 ;
        RECT 563.630 1095.720 572.450 1096.150 ;
        RECT 573.290 1095.720 582.110 1096.150 ;
        RECT 582.950 1095.720 591.770 1096.150 ;
        RECT 592.610 1095.720 601.430 1096.150 ;
        RECT 602.270 1095.720 611.090 1096.150 ;
        RECT 611.930 1095.720 620.750 1096.150 ;
        RECT 621.590 1095.720 630.410 1096.150 ;
        RECT 631.250 1095.720 640.070 1096.150 ;
        RECT 640.910 1095.720 649.730 1096.150 ;
        RECT 650.570 1095.720 659.390 1096.150 ;
        RECT 660.230 1095.720 669.050 1096.150 ;
        RECT 669.890 1095.720 678.710 1096.150 ;
        RECT 679.550 1095.720 688.370 1096.150 ;
        RECT 689.210 1095.720 698.030 1096.150 ;
        RECT 698.870 1095.720 707.690 1096.150 ;
        RECT 708.530 1095.720 717.350 1096.150 ;
        RECT 718.190 1095.720 727.010 1096.150 ;
        RECT 727.850 1095.720 736.670 1096.150 ;
        RECT 737.510 1095.720 745.870 1096.150 ;
        RECT 746.710 1095.720 755.530 1096.150 ;
        RECT 756.370 1095.720 765.190 1096.150 ;
        RECT 766.030 1095.720 774.850 1096.150 ;
        RECT 775.690 1095.720 784.510 1096.150 ;
        RECT 785.350 1095.720 794.170 1096.150 ;
        RECT 795.010 1095.720 803.830 1096.150 ;
        RECT 804.670 1095.720 813.490 1096.150 ;
        RECT 814.330 1095.720 823.150 1096.150 ;
        RECT 823.990 1095.720 832.810 1096.150 ;
        RECT 833.650 1095.720 842.470 1096.150 ;
        RECT 843.310 1095.720 852.130 1096.150 ;
        RECT 852.970 1095.720 861.790 1096.150 ;
        RECT 862.630 1095.720 871.450 1096.150 ;
        RECT 872.290 1095.720 881.110 1096.150 ;
        RECT 881.950 1095.720 890.770 1096.150 ;
        RECT 891.610 1095.720 900.430 1096.150 ;
        RECT 901.270 1095.720 910.090 1096.150 ;
        RECT 910.930 1095.720 919.750 1096.150 ;
        RECT 920.590 1095.720 929.410 1096.150 ;
        RECT 930.250 1095.720 939.070 1096.150 ;
        RECT 939.910 1095.720 948.730 1096.150 ;
        RECT 949.570 1095.720 958.390 1096.150 ;
        RECT 959.230 1095.720 968.050 1096.150 ;
        RECT 968.890 1095.720 977.710 1096.150 ;
        RECT 978.550 1095.720 987.370 1096.150 ;
        RECT 988.210 1095.720 997.030 1096.150 ;
        RECT 997.870 1095.720 1006.690 1096.150 ;
        RECT 1007.530 1095.720 1016.350 1096.150 ;
        RECT 1017.190 1095.720 1026.010 1096.150 ;
        RECT 1026.850 1095.720 1035.670 1096.150 ;
        RECT 1036.510 1095.720 1045.330 1096.150 ;
        RECT 1046.170 1095.720 1054.990 1096.150 ;
        RECT 1055.830 1095.720 1064.650 1096.150 ;
        RECT 1065.490 1095.720 1074.310 1096.150 ;
        RECT 1075.150 1095.720 1083.970 1096.150 ;
        RECT 1084.810 1095.720 1093.630 1096.150 ;
        RECT 1094.470 1095.720 1097.860 1096.150 ;
        RECT 0.030 4.280 1097.860 1095.720 ;
        RECT 0.590 4.000 1.590 4.280 ;
        RECT 2.430 4.000 3.890 4.280 ;
        RECT 4.730 4.000 6.190 4.280 ;
        RECT 7.030 4.000 8.490 4.280 ;
        RECT 9.330 4.000 10.790 4.280 ;
        RECT 11.630 4.000 13.090 4.280 ;
        RECT 13.930 4.000 15.390 4.280 ;
        RECT 16.230 4.000 17.690 4.280 ;
        RECT 18.530 4.000 19.530 4.280 ;
        RECT 20.370 4.000 21.830 4.280 ;
        RECT 22.670 4.000 24.130 4.280 ;
        RECT 24.970 4.000 26.430 4.280 ;
        RECT 27.270 4.000 28.730 4.280 ;
        RECT 29.570 4.000 31.030 4.280 ;
        RECT 31.870 4.000 33.330 4.280 ;
        RECT 34.170 4.000 35.630 4.280 ;
        RECT 36.470 4.000 37.470 4.280 ;
        RECT 38.310 4.000 39.770 4.280 ;
        RECT 40.610 4.000 42.070 4.280 ;
        RECT 42.910 4.000 44.370 4.280 ;
        RECT 45.210 4.000 46.670 4.280 ;
        RECT 47.510 4.000 48.970 4.280 ;
        RECT 49.810 4.000 51.270 4.280 ;
        RECT 52.110 4.000 53.570 4.280 ;
        RECT 54.410 4.000 55.410 4.280 ;
        RECT 56.250 4.000 57.710 4.280 ;
        RECT 58.550 4.000 60.010 4.280 ;
        RECT 60.850 4.000 62.310 4.280 ;
        RECT 63.150 4.000 64.610 4.280 ;
        RECT 65.450 4.000 66.910 4.280 ;
        RECT 67.750 4.000 69.210 4.280 ;
        RECT 70.050 4.000 71.510 4.280 ;
        RECT 72.350 4.000 73.810 4.280 ;
        RECT 74.650 4.000 75.650 4.280 ;
        RECT 76.490 4.000 77.950 4.280 ;
        RECT 78.790 4.000 80.250 4.280 ;
        RECT 81.090 4.000 82.550 4.280 ;
        RECT 83.390 4.000 84.850 4.280 ;
        RECT 85.690 4.000 87.150 4.280 ;
        RECT 87.990 4.000 89.450 4.280 ;
        RECT 90.290 4.000 91.750 4.280 ;
        RECT 92.590 4.000 93.590 4.280 ;
        RECT 94.430 4.000 95.890 4.280 ;
        RECT 96.730 4.000 98.190 4.280 ;
        RECT 99.030 4.000 100.490 4.280 ;
        RECT 101.330 4.000 102.790 4.280 ;
        RECT 103.630 4.000 105.090 4.280 ;
        RECT 105.930 4.000 107.390 4.280 ;
        RECT 108.230 4.000 109.690 4.280 ;
        RECT 110.530 4.000 111.530 4.280 ;
        RECT 112.370 4.000 113.830 4.280 ;
        RECT 114.670 4.000 116.130 4.280 ;
        RECT 116.970 4.000 118.430 4.280 ;
        RECT 119.270 4.000 120.730 4.280 ;
        RECT 121.570 4.000 123.030 4.280 ;
        RECT 123.870 4.000 125.330 4.280 ;
        RECT 126.170 4.000 127.630 4.280 ;
        RECT 128.470 4.000 129.930 4.280 ;
        RECT 130.770 4.000 131.770 4.280 ;
        RECT 132.610 4.000 134.070 4.280 ;
        RECT 134.910 4.000 136.370 4.280 ;
        RECT 137.210 4.000 138.670 4.280 ;
        RECT 139.510 4.000 140.970 4.280 ;
        RECT 141.810 4.000 143.270 4.280 ;
        RECT 144.110 4.000 145.570 4.280 ;
        RECT 146.410 4.000 147.870 4.280 ;
        RECT 148.710 4.000 149.710 4.280 ;
        RECT 150.550 4.000 152.010 4.280 ;
        RECT 152.850 4.000 154.310 4.280 ;
        RECT 155.150 4.000 156.610 4.280 ;
        RECT 157.450 4.000 158.910 4.280 ;
        RECT 159.750 4.000 161.210 4.280 ;
        RECT 162.050 4.000 163.510 4.280 ;
        RECT 164.350 4.000 165.810 4.280 ;
        RECT 166.650 4.000 167.650 4.280 ;
        RECT 168.490 4.000 169.950 4.280 ;
        RECT 170.790 4.000 172.250 4.280 ;
        RECT 173.090 4.000 174.550 4.280 ;
        RECT 175.390 4.000 176.850 4.280 ;
        RECT 177.690 4.000 179.150 4.280 ;
        RECT 179.990 4.000 181.450 4.280 ;
        RECT 182.290 4.000 183.750 4.280 ;
        RECT 184.590 4.000 186.050 4.280 ;
        RECT 186.890 4.000 187.890 4.280 ;
        RECT 188.730 4.000 190.190 4.280 ;
        RECT 191.030 4.000 192.490 4.280 ;
        RECT 193.330 4.000 194.790 4.280 ;
        RECT 195.630 4.000 197.090 4.280 ;
        RECT 197.930 4.000 199.390 4.280 ;
        RECT 200.230 4.000 201.690 4.280 ;
        RECT 202.530 4.000 203.990 4.280 ;
        RECT 204.830 4.000 205.830 4.280 ;
        RECT 206.670 4.000 208.130 4.280 ;
        RECT 208.970 4.000 210.430 4.280 ;
        RECT 211.270 4.000 212.730 4.280 ;
        RECT 213.570 4.000 215.030 4.280 ;
        RECT 215.870 4.000 217.330 4.280 ;
        RECT 218.170 4.000 219.630 4.280 ;
        RECT 220.470 4.000 221.930 4.280 ;
        RECT 222.770 4.000 223.770 4.280 ;
        RECT 224.610 4.000 226.070 4.280 ;
        RECT 226.910 4.000 228.370 4.280 ;
        RECT 229.210 4.000 230.670 4.280 ;
        RECT 231.510 4.000 232.970 4.280 ;
        RECT 233.810 4.000 235.270 4.280 ;
        RECT 236.110 4.000 237.570 4.280 ;
        RECT 238.410 4.000 239.870 4.280 ;
        RECT 240.710 4.000 241.710 4.280 ;
        RECT 242.550 4.000 244.010 4.280 ;
        RECT 244.850 4.000 246.310 4.280 ;
        RECT 247.150 4.000 248.610 4.280 ;
        RECT 249.450 4.000 250.910 4.280 ;
        RECT 251.750 4.000 253.210 4.280 ;
        RECT 254.050 4.000 255.510 4.280 ;
        RECT 256.350 4.000 257.810 4.280 ;
        RECT 258.650 4.000 260.110 4.280 ;
        RECT 260.950 4.000 261.950 4.280 ;
        RECT 262.790 4.000 264.250 4.280 ;
        RECT 265.090 4.000 266.550 4.280 ;
        RECT 267.390 4.000 268.850 4.280 ;
        RECT 269.690 4.000 271.150 4.280 ;
        RECT 271.990 4.000 273.450 4.280 ;
        RECT 274.290 4.000 275.750 4.280 ;
        RECT 276.590 4.000 278.050 4.280 ;
        RECT 278.890 4.000 279.890 4.280 ;
        RECT 280.730 4.000 282.190 4.280 ;
        RECT 283.030 4.000 284.490 4.280 ;
        RECT 285.330 4.000 286.790 4.280 ;
        RECT 287.630 4.000 289.090 4.280 ;
        RECT 289.930 4.000 291.390 4.280 ;
        RECT 292.230 4.000 293.690 4.280 ;
        RECT 294.530 4.000 295.990 4.280 ;
        RECT 296.830 4.000 297.830 4.280 ;
        RECT 298.670 4.000 300.130 4.280 ;
        RECT 300.970 4.000 302.430 4.280 ;
        RECT 303.270 4.000 304.730 4.280 ;
        RECT 305.570 4.000 307.030 4.280 ;
        RECT 307.870 4.000 309.330 4.280 ;
        RECT 310.170 4.000 311.630 4.280 ;
        RECT 312.470 4.000 313.930 4.280 ;
        RECT 314.770 4.000 316.230 4.280 ;
        RECT 317.070 4.000 318.070 4.280 ;
        RECT 318.910 4.000 320.370 4.280 ;
        RECT 321.210 4.000 322.670 4.280 ;
        RECT 323.510 4.000 324.970 4.280 ;
        RECT 325.810 4.000 327.270 4.280 ;
        RECT 328.110 4.000 329.570 4.280 ;
        RECT 330.410 4.000 331.870 4.280 ;
        RECT 332.710 4.000 334.170 4.280 ;
        RECT 335.010 4.000 336.010 4.280 ;
        RECT 336.850 4.000 338.310 4.280 ;
        RECT 339.150 4.000 340.610 4.280 ;
        RECT 341.450 4.000 342.910 4.280 ;
        RECT 343.750 4.000 345.210 4.280 ;
        RECT 346.050 4.000 347.510 4.280 ;
        RECT 348.350 4.000 349.810 4.280 ;
        RECT 350.650 4.000 352.110 4.280 ;
        RECT 352.950 4.000 353.950 4.280 ;
        RECT 354.790 4.000 356.250 4.280 ;
        RECT 357.090 4.000 358.550 4.280 ;
        RECT 359.390 4.000 360.850 4.280 ;
        RECT 361.690 4.000 363.150 4.280 ;
        RECT 363.990 4.000 365.450 4.280 ;
        RECT 366.290 4.000 367.750 4.280 ;
        RECT 368.590 4.000 370.050 4.280 ;
        RECT 370.890 4.000 372.350 4.280 ;
        RECT 373.190 4.000 374.190 4.280 ;
        RECT 375.030 4.000 376.490 4.280 ;
        RECT 377.330 4.000 378.790 4.280 ;
        RECT 379.630 4.000 381.090 4.280 ;
        RECT 381.930 4.000 383.390 4.280 ;
        RECT 384.230 4.000 385.690 4.280 ;
        RECT 386.530 4.000 387.990 4.280 ;
        RECT 388.830 4.000 390.290 4.280 ;
        RECT 391.130 4.000 392.130 4.280 ;
        RECT 392.970 4.000 394.430 4.280 ;
        RECT 395.270 4.000 396.730 4.280 ;
        RECT 397.570 4.000 399.030 4.280 ;
        RECT 399.870 4.000 401.330 4.280 ;
        RECT 402.170 4.000 403.630 4.280 ;
        RECT 404.470 4.000 405.930 4.280 ;
        RECT 406.770 4.000 408.230 4.280 ;
        RECT 409.070 4.000 410.070 4.280 ;
        RECT 410.910 4.000 412.370 4.280 ;
        RECT 413.210 4.000 414.670 4.280 ;
        RECT 415.510 4.000 416.970 4.280 ;
        RECT 417.810 4.000 419.270 4.280 ;
        RECT 420.110 4.000 421.570 4.280 ;
        RECT 422.410 4.000 423.870 4.280 ;
        RECT 424.710 4.000 426.170 4.280 ;
        RECT 427.010 4.000 428.470 4.280 ;
        RECT 429.310 4.000 430.310 4.280 ;
        RECT 431.150 4.000 432.610 4.280 ;
        RECT 433.450 4.000 434.910 4.280 ;
        RECT 435.750 4.000 437.210 4.280 ;
        RECT 438.050 4.000 439.510 4.280 ;
        RECT 440.350 4.000 441.810 4.280 ;
        RECT 442.650 4.000 444.110 4.280 ;
        RECT 444.950 4.000 446.410 4.280 ;
        RECT 447.250 4.000 448.250 4.280 ;
        RECT 449.090 4.000 450.550 4.280 ;
        RECT 451.390 4.000 452.850 4.280 ;
        RECT 453.690 4.000 455.150 4.280 ;
        RECT 455.990 4.000 457.450 4.280 ;
        RECT 458.290 4.000 459.750 4.280 ;
        RECT 460.590 4.000 462.050 4.280 ;
        RECT 462.890 4.000 464.350 4.280 ;
        RECT 465.190 4.000 466.190 4.280 ;
        RECT 467.030 4.000 468.490 4.280 ;
        RECT 469.330 4.000 470.790 4.280 ;
        RECT 471.630 4.000 473.090 4.280 ;
        RECT 473.930 4.000 475.390 4.280 ;
        RECT 476.230 4.000 477.690 4.280 ;
        RECT 478.530 4.000 479.990 4.280 ;
        RECT 480.830 4.000 482.290 4.280 ;
        RECT 483.130 4.000 484.130 4.280 ;
        RECT 484.970 4.000 486.430 4.280 ;
        RECT 487.270 4.000 488.730 4.280 ;
        RECT 489.570 4.000 491.030 4.280 ;
        RECT 491.870 4.000 493.330 4.280 ;
        RECT 494.170 4.000 495.630 4.280 ;
        RECT 496.470 4.000 497.930 4.280 ;
        RECT 498.770 4.000 500.230 4.280 ;
        RECT 501.070 4.000 502.530 4.280 ;
        RECT 503.370 4.000 504.370 4.280 ;
        RECT 505.210 4.000 506.670 4.280 ;
        RECT 507.510 4.000 508.970 4.280 ;
        RECT 509.810 4.000 511.270 4.280 ;
        RECT 512.110 4.000 513.570 4.280 ;
        RECT 514.410 4.000 515.870 4.280 ;
        RECT 516.710 4.000 518.170 4.280 ;
        RECT 519.010 4.000 520.470 4.280 ;
        RECT 521.310 4.000 522.310 4.280 ;
        RECT 523.150 4.000 524.610 4.280 ;
        RECT 525.450 4.000 526.910 4.280 ;
        RECT 527.750 4.000 529.210 4.280 ;
        RECT 530.050 4.000 531.510 4.280 ;
        RECT 532.350 4.000 533.810 4.280 ;
        RECT 534.650 4.000 536.110 4.280 ;
        RECT 536.950 4.000 538.410 4.280 ;
        RECT 539.250 4.000 540.250 4.280 ;
        RECT 541.090 4.000 542.550 4.280 ;
        RECT 543.390 4.000 544.850 4.280 ;
        RECT 545.690 4.000 547.150 4.280 ;
        RECT 547.990 4.000 549.450 4.280 ;
        RECT 550.290 4.000 551.750 4.280 ;
        RECT 552.590 4.000 554.050 4.280 ;
        RECT 554.890 4.000 556.350 4.280 ;
        RECT 557.190 4.000 558.650 4.280 ;
        RECT 559.490 4.000 560.490 4.280 ;
        RECT 561.330 4.000 562.790 4.280 ;
        RECT 563.630 4.000 565.090 4.280 ;
        RECT 565.930 4.000 567.390 4.280 ;
        RECT 568.230 4.000 569.690 4.280 ;
        RECT 570.530 4.000 571.990 4.280 ;
        RECT 572.830 4.000 574.290 4.280 ;
        RECT 575.130 4.000 576.590 4.280 ;
        RECT 577.430 4.000 578.430 4.280 ;
        RECT 579.270 4.000 580.730 4.280 ;
        RECT 581.570 4.000 583.030 4.280 ;
        RECT 583.870 4.000 585.330 4.280 ;
        RECT 586.170 4.000 587.630 4.280 ;
        RECT 588.470 4.000 589.930 4.280 ;
        RECT 590.770 4.000 592.230 4.280 ;
        RECT 593.070 4.000 594.530 4.280 ;
        RECT 595.370 4.000 596.370 4.280 ;
        RECT 597.210 4.000 598.670 4.280 ;
        RECT 599.510 4.000 600.970 4.280 ;
        RECT 601.810 4.000 603.270 4.280 ;
        RECT 604.110 4.000 605.570 4.280 ;
        RECT 606.410 4.000 607.870 4.280 ;
        RECT 608.710 4.000 610.170 4.280 ;
        RECT 611.010 4.000 612.470 4.280 ;
        RECT 613.310 4.000 614.770 4.280 ;
        RECT 615.610 4.000 616.610 4.280 ;
        RECT 617.450 4.000 618.910 4.280 ;
        RECT 619.750 4.000 621.210 4.280 ;
        RECT 622.050 4.000 623.510 4.280 ;
        RECT 624.350 4.000 625.810 4.280 ;
        RECT 626.650 4.000 628.110 4.280 ;
        RECT 628.950 4.000 630.410 4.280 ;
        RECT 631.250 4.000 632.710 4.280 ;
        RECT 633.550 4.000 634.550 4.280 ;
        RECT 635.390 4.000 636.850 4.280 ;
        RECT 637.690 4.000 639.150 4.280 ;
        RECT 639.990 4.000 641.450 4.280 ;
        RECT 642.290 4.000 643.750 4.280 ;
        RECT 644.590 4.000 646.050 4.280 ;
        RECT 646.890 4.000 648.350 4.280 ;
        RECT 649.190 4.000 650.650 4.280 ;
        RECT 651.490 4.000 652.490 4.280 ;
        RECT 653.330 4.000 654.790 4.280 ;
        RECT 655.630 4.000 657.090 4.280 ;
        RECT 657.930 4.000 659.390 4.280 ;
        RECT 660.230 4.000 661.690 4.280 ;
        RECT 662.530 4.000 663.990 4.280 ;
        RECT 664.830 4.000 666.290 4.280 ;
        RECT 667.130 4.000 668.590 4.280 ;
        RECT 669.430 4.000 670.430 4.280 ;
        RECT 671.270 4.000 672.730 4.280 ;
        RECT 673.570 4.000 675.030 4.280 ;
        RECT 675.870 4.000 677.330 4.280 ;
        RECT 678.170 4.000 679.630 4.280 ;
        RECT 680.470 4.000 681.930 4.280 ;
        RECT 682.770 4.000 684.230 4.280 ;
        RECT 685.070 4.000 686.530 4.280 ;
        RECT 687.370 4.000 688.830 4.280 ;
        RECT 689.670 4.000 690.670 4.280 ;
        RECT 691.510 4.000 692.970 4.280 ;
        RECT 693.810 4.000 695.270 4.280 ;
        RECT 696.110 4.000 697.570 4.280 ;
        RECT 698.410 4.000 699.870 4.280 ;
        RECT 700.710 4.000 702.170 4.280 ;
        RECT 703.010 4.000 704.470 4.280 ;
        RECT 705.310 4.000 706.770 4.280 ;
        RECT 707.610 4.000 708.610 4.280 ;
        RECT 709.450 4.000 710.910 4.280 ;
        RECT 711.750 4.000 713.210 4.280 ;
        RECT 714.050 4.000 715.510 4.280 ;
        RECT 716.350 4.000 717.810 4.280 ;
        RECT 718.650 4.000 720.110 4.280 ;
        RECT 720.950 4.000 722.410 4.280 ;
        RECT 723.250 4.000 724.710 4.280 ;
        RECT 725.550 4.000 726.550 4.280 ;
        RECT 727.390 4.000 728.850 4.280 ;
        RECT 729.690 4.000 731.150 4.280 ;
        RECT 731.990 4.000 733.450 4.280 ;
        RECT 734.290 4.000 735.750 4.280 ;
        RECT 736.590 4.000 738.050 4.280 ;
        RECT 738.890 4.000 740.350 4.280 ;
        RECT 741.190 4.000 742.650 4.280 ;
        RECT 743.490 4.000 744.950 4.280 ;
        RECT 745.790 4.000 746.790 4.280 ;
        RECT 747.630 4.000 749.090 4.280 ;
        RECT 749.930 4.000 751.390 4.280 ;
        RECT 752.230 4.000 753.690 4.280 ;
        RECT 754.530 4.000 755.990 4.280 ;
        RECT 756.830 4.000 758.290 4.280 ;
        RECT 759.130 4.000 760.590 4.280 ;
        RECT 761.430 4.000 762.890 4.280 ;
        RECT 763.730 4.000 764.730 4.280 ;
        RECT 765.570 4.000 767.030 4.280 ;
        RECT 767.870 4.000 769.330 4.280 ;
        RECT 770.170 4.000 771.630 4.280 ;
        RECT 772.470 4.000 773.930 4.280 ;
        RECT 774.770 4.000 776.230 4.280 ;
        RECT 777.070 4.000 778.530 4.280 ;
        RECT 779.370 4.000 780.830 4.280 ;
        RECT 781.670 4.000 782.670 4.280 ;
        RECT 783.510 4.000 784.970 4.280 ;
        RECT 785.810 4.000 787.270 4.280 ;
        RECT 788.110 4.000 789.570 4.280 ;
        RECT 790.410 4.000 791.870 4.280 ;
        RECT 792.710 4.000 794.170 4.280 ;
        RECT 795.010 4.000 796.470 4.280 ;
        RECT 797.310 4.000 798.770 4.280 ;
        RECT 799.610 4.000 801.070 4.280 ;
        RECT 801.910 4.000 802.910 4.280 ;
        RECT 803.750 4.000 805.210 4.280 ;
        RECT 806.050 4.000 807.510 4.280 ;
        RECT 808.350 4.000 809.810 4.280 ;
        RECT 810.650 4.000 812.110 4.280 ;
        RECT 812.950 4.000 814.410 4.280 ;
        RECT 815.250 4.000 816.710 4.280 ;
        RECT 817.550 4.000 819.010 4.280 ;
        RECT 819.850 4.000 820.850 4.280 ;
        RECT 821.690 4.000 823.150 4.280 ;
        RECT 823.990 4.000 825.450 4.280 ;
        RECT 826.290 4.000 827.750 4.280 ;
        RECT 828.590 4.000 830.050 4.280 ;
        RECT 830.890 4.000 832.350 4.280 ;
        RECT 833.190 4.000 834.650 4.280 ;
        RECT 835.490 4.000 836.950 4.280 ;
        RECT 837.790 4.000 838.790 4.280 ;
        RECT 839.630 4.000 841.090 4.280 ;
        RECT 841.930 4.000 843.390 4.280 ;
        RECT 844.230 4.000 845.690 4.280 ;
        RECT 846.530 4.000 847.990 4.280 ;
        RECT 848.830 4.000 850.290 4.280 ;
        RECT 851.130 4.000 852.590 4.280 ;
        RECT 853.430 4.000 854.890 4.280 ;
        RECT 855.730 4.000 857.190 4.280 ;
        RECT 858.030 4.000 859.030 4.280 ;
        RECT 859.870 4.000 861.330 4.280 ;
        RECT 862.170 4.000 863.630 4.280 ;
        RECT 864.470 4.000 865.930 4.280 ;
        RECT 866.770 4.000 868.230 4.280 ;
        RECT 869.070 4.000 870.530 4.280 ;
        RECT 871.370 4.000 872.830 4.280 ;
        RECT 873.670 4.000 875.130 4.280 ;
        RECT 875.970 4.000 876.970 4.280 ;
        RECT 877.810 4.000 879.270 4.280 ;
        RECT 880.110 4.000 881.570 4.280 ;
        RECT 882.410 4.000 883.870 4.280 ;
        RECT 884.710 4.000 886.170 4.280 ;
        RECT 887.010 4.000 888.470 4.280 ;
        RECT 889.310 4.000 890.770 4.280 ;
        RECT 891.610 4.000 893.070 4.280 ;
        RECT 893.910 4.000 894.910 4.280 ;
        RECT 895.750 4.000 897.210 4.280 ;
        RECT 898.050 4.000 899.510 4.280 ;
        RECT 900.350 4.000 901.810 4.280 ;
        RECT 902.650 4.000 904.110 4.280 ;
        RECT 904.950 4.000 906.410 4.280 ;
        RECT 907.250 4.000 908.710 4.280 ;
        RECT 909.550 4.000 911.010 4.280 ;
        RECT 911.850 4.000 912.850 4.280 ;
        RECT 913.690 4.000 915.150 4.280 ;
        RECT 915.990 4.000 917.450 4.280 ;
        RECT 918.290 4.000 919.750 4.280 ;
        RECT 920.590 4.000 922.050 4.280 ;
        RECT 922.890 4.000 924.350 4.280 ;
        RECT 925.190 4.000 926.650 4.280 ;
        RECT 927.490 4.000 928.950 4.280 ;
        RECT 929.790 4.000 931.250 4.280 ;
        RECT 932.090 4.000 933.090 4.280 ;
        RECT 933.930 4.000 935.390 4.280 ;
        RECT 936.230 4.000 937.690 4.280 ;
        RECT 938.530 4.000 939.990 4.280 ;
        RECT 940.830 4.000 942.290 4.280 ;
        RECT 943.130 4.000 944.590 4.280 ;
        RECT 945.430 4.000 946.890 4.280 ;
        RECT 947.730 4.000 949.190 4.280 ;
        RECT 950.030 4.000 951.030 4.280 ;
        RECT 951.870 4.000 953.330 4.280 ;
        RECT 954.170 4.000 955.630 4.280 ;
        RECT 956.470 4.000 957.930 4.280 ;
        RECT 958.770 4.000 960.230 4.280 ;
        RECT 961.070 4.000 962.530 4.280 ;
        RECT 963.370 4.000 964.830 4.280 ;
        RECT 965.670 4.000 967.130 4.280 ;
        RECT 967.970 4.000 968.970 4.280 ;
        RECT 969.810 4.000 971.270 4.280 ;
        RECT 972.110 4.000 973.570 4.280 ;
        RECT 974.410 4.000 975.870 4.280 ;
        RECT 976.710 4.000 978.170 4.280 ;
        RECT 979.010 4.000 980.470 4.280 ;
        RECT 981.310 4.000 982.770 4.280 ;
        RECT 983.610 4.000 985.070 4.280 ;
        RECT 985.910 4.000 987.370 4.280 ;
        RECT 988.210 4.000 989.210 4.280 ;
        RECT 990.050 4.000 991.510 4.280 ;
        RECT 992.350 4.000 993.810 4.280 ;
        RECT 994.650 4.000 996.110 4.280 ;
        RECT 996.950 4.000 998.410 4.280 ;
        RECT 999.250 4.000 1000.710 4.280 ;
        RECT 1001.550 4.000 1003.010 4.280 ;
        RECT 1003.850 4.000 1005.310 4.280 ;
        RECT 1006.150 4.000 1007.150 4.280 ;
        RECT 1007.990 4.000 1009.450 4.280 ;
        RECT 1010.290 4.000 1011.750 4.280 ;
        RECT 1012.590 4.000 1014.050 4.280 ;
        RECT 1014.890 4.000 1016.350 4.280 ;
        RECT 1017.190 4.000 1018.650 4.280 ;
        RECT 1019.490 4.000 1020.950 4.280 ;
        RECT 1021.790 4.000 1023.250 4.280 ;
        RECT 1024.090 4.000 1025.090 4.280 ;
        RECT 1025.930 4.000 1027.390 4.280 ;
        RECT 1028.230 4.000 1029.690 4.280 ;
        RECT 1030.530 4.000 1031.990 4.280 ;
        RECT 1032.830 4.000 1034.290 4.280 ;
        RECT 1035.130 4.000 1036.590 4.280 ;
        RECT 1037.430 4.000 1038.890 4.280 ;
        RECT 1039.730 4.000 1041.190 4.280 ;
        RECT 1042.030 4.000 1043.490 4.280 ;
        RECT 1044.330 4.000 1045.330 4.280 ;
        RECT 1046.170 4.000 1047.630 4.280 ;
        RECT 1048.470 4.000 1049.930 4.280 ;
        RECT 1050.770 4.000 1052.230 4.280 ;
        RECT 1053.070 4.000 1054.530 4.280 ;
        RECT 1055.370 4.000 1056.830 4.280 ;
        RECT 1057.670 4.000 1059.130 4.280 ;
        RECT 1059.970 4.000 1061.430 4.280 ;
        RECT 1062.270 4.000 1063.270 4.280 ;
        RECT 1064.110 4.000 1065.570 4.280 ;
        RECT 1066.410 4.000 1067.870 4.280 ;
        RECT 1068.710 4.000 1070.170 4.280 ;
        RECT 1071.010 4.000 1072.470 4.280 ;
        RECT 1073.310 4.000 1074.770 4.280 ;
        RECT 1075.610 4.000 1077.070 4.280 ;
        RECT 1077.910 4.000 1079.370 4.280 ;
        RECT 1080.210 4.000 1081.210 4.280 ;
        RECT 1082.050 4.000 1083.510 4.280 ;
        RECT 1084.350 4.000 1085.810 4.280 ;
        RECT 1086.650 4.000 1088.110 4.280 ;
        RECT 1088.950 4.000 1090.410 4.280 ;
        RECT 1091.250 4.000 1092.710 4.280 ;
        RECT 1093.550 4.000 1095.010 4.280 ;
        RECT 1095.850 4.000 1097.310 4.280 ;
      LAYER met3 ;
        RECT 0.005 4.255 1079.035 1088.165 ;
      LAYER met4 ;
        RECT 45.315 10.640 96.460 1088.240 ;
        RECT 98.860 10.640 1068.685 1088.240 ;
  END
END user_proj_example
END LIBRARY

