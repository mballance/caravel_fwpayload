magic
tech sky130A
magscale 1 2
timestamp 1608083996
<< obsli1 >>
rect 908 2159 238636 237745
<< obsm1 >>
rect 908 1096 239542 237776
<< metal2 >>
rect 834 239200 890 240000
rect 2858 239200 2914 240000
rect 4974 239200 5030 240000
rect 7090 239200 7146 240000
rect 9206 239200 9262 240000
rect 11322 239200 11378 240000
rect 13438 239200 13494 240000
rect 15554 239200 15610 240000
rect 17670 239200 17726 240000
rect 19694 239200 19750 240000
rect 21810 239200 21866 240000
rect 23926 239200 23982 240000
rect 26042 239200 26098 240000
rect 28158 239200 28214 240000
rect 30274 239200 30330 240000
rect 32390 239200 32446 240000
rect 34506 239200 34562 240000
rect 36622 239200 36678 240000
rect 38646 239200 38702 240000
rect 40762 239200 40818 240000
rect 42878 239200 42934 240000
rect 44994 239200 45050 240000
rect 47110 239200 47166 240000
rect 49226 239200 49282 240000
rect 51342 239200 51398 240000
rect 53458 239200 53514 240000
rect 55574 239200 55630 240000
rect 57598 239200 57654 240000
rect 59714 239200 59770 240000
rect 61830 239200 61886 240000
rect 63946 239200 64002 240000
rect 66062 239200 66118 240000
rect 68178 239200 68234 240000
rect 70294 239200 70350 240000
rect 72410 239200 72466 240000
rect 74526 239200 74582 240000
rect 76550 239200 76606 240000
rect 78666 239200 78722 240000
rect 80782 239200 80838 240000
rect 82898 239200 82954 240000
rect 85014 239200 85070 240000
rect 87130 239200 87186 240000
rect 89246 239200 89302 240000
rect 91362 239200 91418 240000
rect 93386 239200 93442 240000
rect 95502 239200 95558 240000
rect 97618 239200 97674 240000
rect 99734 239200 99790 240000
rect 101850 239200 101906 240000
rect 103966 239200 104022 240000
rect 106082 239200 106138 240000
rect 108198 239200 108254 240000
rect 110314 239200 110370 240000
rect 112338 239200 112394 240000
rect 114454 239200 114510 240000
rect 116570 239200 116626 240000
rect 118686 239200 118742 240000
rect 120802 239200 120858 240000
rect 122918 239200 122974 240000
rect 125034 239200 125090 240000
rect 127150 239200 127206 240000
rect 129266 239200 129322 240000
rect 131290 239200 131346 240000
rect 133406 239200 133462 240000
rect 135522 239200 135578 240000
rect 137638 239200 137694 240000
rect 139754 239200 139810 240000
rect 141870 239200 141926 240000
rect 143986 239200 144042 240000
rect 146102 239200 146158 240000
rect 148218 239200 148274 240000
rect 150242 239200 150298 240000
rect 152358 239200 152414 240000
rect 154474 239200 154530 240000
rect 156590 239200 156646 240000
rect 158706 239200 158762 240000
rect 160822 239200 160878 240000
rect 162938 239200 162994 240000
rect 165054 239200 165110 240000
rect 167078 239200 167134 240000
rect 169194 239200 169250 240000
rect 171310 239200 171366 240000
rect 173426 239200 173482 240000
rect 175542 239200 175598 240000
rect 177658 239200 177714 240000
rect 179774 239200 179830 240000
rect 181890 239200 181946 240000
rect 184006 239200 184062 240000
rect 186030 239200 186086 240000
rect 188146 239200 188202 240000
rect 190262 239200 190318 240000
rect 192378 239200 192434 240000
rect 194494 239200 194550 240000
rect 196610 239200 196666 240000
rect 198726 239200 198782 240000
rect 200842 239200 200898 240000
rect 202958 239200 203014 240000
rect 204982 239200 205038 240000
rect 207098 239200 207154 240000
rect 209214 239200 209270 240000
rect 211330 239200 211386 240000
rect 213446 239200 213502 240000
rect 215562 239200 215618 240000
rect 217678 239200 217734 240000
rect 219794 239200 219850 240000
rect 221910 239200 221966 240000
rect 223934 239200 223990 240000
rect 226050 239200 226106 240000
rect 228166 239200 228222 240000
rect 230282 239200 230338 240000
rect 232398 239200 232454 240000
rect 234514 239200 234570 240000
rect 236630 239200 236686 240000
rect 238746 239200 238802 240000
rect 6 0 62 800
rect 466 0 522 800
rect 926 0 982 800
rect 1386 0 1442 800
rect 1938 0 1994 800
rect 2398 0 2454 800
rect 2858 0 2914 800
rect 3410 0 3466 800
rect 3870 0 3926 800
rect 4330 0 4386 800
rect 4882 0 4938 800
rect 5342 0 5398 800
rect 5802 0 5858 800
rect 6354 0 6410 800
rect 6814 0 6870 800
rect 7274 0 7330 800
rect 7826 0 7882 800
rect 8286 0 8342 800
rect 8746 0 8802 800
rect 9298 0 9354 800
rect 9758 0 9814 800
rect 10218 0 10274 800
rect 10770 0 10826 800
rect 11230 0 11286 800
rect 11690 0 11746 800
rect 12242 0 12298 800
rect 12702 0 12758 800
rect 13162 0 13218 800
rect 13714 0 13770 800
rect 14174 0 14230 800
rect 14634 0 14690 800
rect 15186 0 15242 800
rect 15646 0 15702 800
rect 16106 0 16162 800
rect 16658 0 16714 800
rect 17118 0 17174 800
rect 17578 0 17634 800
rect 18130 0 18186 800
rect 18590 0 18646 800
rect 19050 0 19106 800
rect 19510 0 19566 800
rect 20062 0 20118 800
rect 20522 0 20578 800
rect 20982 0 21038 800
rect 21534 0 21590 800
rect 21994 0 22050 800
rect 22454 0 22510 800
rect 23006 0 23062 800
rect 23466 0 23522 800
rect 23926 0 23982 800
rect 24478 0 24534 800
rect 24938 0 24994 800
rect 25398 0 25454 800
rect 25950 0 26006 800
rect 26410 0 26466 800
rect 26870 0 26926 800
rect 27422 0 27478 800
rect 27882 0 27938 800
rect 28342 0 28398 800
rect 28894 0 28950 800
rect 29354 0 29410 800
rect 29814 0 29870 800
rect 30366 0 30422 800
rect 30826 0 30882 800
rect 31286 0 31342 800
rect 31838 0 31894 800
rect 32298 0 32354 800
rect 32758 0 32814 800
rect 33310 0 33366 800
rect 33770 0 33826 800
rect 34230 0 34286 800
rect 34782 0 34838 800
rect 35242 0 35298 800
rect 35702 0 35758 800
rect 36254 0 36310 800
rect 36714 0 36770 800
rect 37174 0 37230 800
rect 37634 0 37690 800
rect 38186 0 38242 800
rect 38646 0 38702 800
rect 39106 0 39162 800
rect 39658 0 39714 800
rect 40118 0 40174 800
rect 40578 0 40634 800
rect 41130 0 41186 800
rect 41590 0 41646 800
rect 42050 0 42106 800
rect 42602 0 42658 800
rect 43062 0 43118 800
rect 43522 0 43578 800
rect 44074 0 44130 800
rect 44534 0 44590 800
rect 44994 0 45050 800
rect 45546 0 45602 800
rect 46006 0 46062 800
rect 46466 0 46522 800
rect 47018 0 47074 800
rect 47478 0 47534 800
rect 47938 0 47994 800
rect 48490 0 48546 800
rect 48950 0 49006 800
rect 49410 0 49466 800
rect 49962 0 50018 800
rect 50422 0 50478 800
rect 50882 0 50938 800
rect 51434 0 51490 800
rect 51894 0 51950 800
rect 52354 0 52410 800
rect 52906 0 52962 800
rect 53366 0 53422 800
rect 53826 0 53882 800
rect 54378 0 54434 800
rect 54838 0 54894 800
rect 55298 0 55354 800
rect 55758 0 55814 800
rect 56310 0 56366 800
rect 56770 0 56826 800
rect 57230 0 57286 800
rect 57782 0 57838 800
rect 58242 0 58298 800
rect 58702 0 58758 800
rect 59254 0 59310 800
rect 59714 0 59770 800
rect 60174 0 60230 800
rect 60726 0 60782 800
rect 61186 0 61242 800
rect 61646 0 61702 800
rect 62198 0 62254 800
rect 62658 0 62714 800
rect 63118 0 63174 800
rect 63670 0 63726 800
rect 64130 0 64186 800
rect 64590 0 64646 800
rect 65142 0 65198 800
rect 65602 0 65658 800
rect 66062 0 66118 800
rect 66614 0 66670 800
rect 67074 0 67130 800
rect 67534 0 67590 800
rect 68086 0 68142 800
rect 68546 0 68602 800
rect 69006 0 69062 800
rect 69558 0 69614 800
rect 70018 0 70074 800
rect 70478 0 70534 800
rect 71030 0 71086 800
rect 71490 0 71546 800
rect 71950 0 72006 800
rect 72502 0 72558 800
rect 72962 0 73018 800
rect 73422 0 73478 800
rect 73882 0 73938 800
rect 74434 0 74490 800
rect 74894 0 74950 800
rect 75354 0 75410 800
rect 75906 0 75962 800
rect 76366 0 76422 800
rect 76826 0 76882 800
rect 77378 0 77434 800
rect 77838 0 77894 800
rect 78298 0 78354 800
rect 78850 0 78906 800
rect 79310 0 79366 800
rect 79770 0 79826 800
rect 80322 0 80378 800
rect 80782 0 80838 800
rect 81242 0 81298 800
rect 81794 0 81850 800
rect 82254 0 82310 800
rect 82714 0 82770 800
rect 83266 0 83322 800
rect 83726 0 83782 800
rect 84186 0 84242 800
rect 84738 0 84794 800
rect 85198 0 85254 800
rect 85658 0 85714 800
rect 86210 0 86266 800
rect 86670 0 86726 800
rect 87130 0 87186 800
rect 87682 0 87738 800
rect 88142 0 88198 800
rect 88602 0 88658 800
rect 89154 0 89210 800
rect 89614 0 89670 800
rect 90074 0 90130 800
rect 90626 0 90682 800
rect 91086 0 91142 800
rect 91546 0 91602 800
rect 92098 0 92154 800
rect 92558 0 92614 800
rect 93018 0 93074 800
rect 93478 0 93534 800
rect 94030 0 94086 800
rect 94490 0 94546 800
rect 94950 0 95006 800
rect 95502 0 95558 800
rect 95962 0 96018 800
rect 96422 0 96478 800
rect 96974 0 97030 800
rect 97434 0 97490 800
rect 97894 0 97950 800
rect 98446 0 98502 800
rect 98906 0 98962 800
rect 99366 0 99422 800
rect 99918 0 99974 800
rect 100378 0 100434 800
rect 100838 0 100894 800
rect 101390 0 101446 800
rect 101850 0 101906 800
rect 102310 0 102366 800
rect 102862 0 102918 800
rect 103322 0 103378 800
rect 103782 0 103838 800
rect 104334 0 104390 800
rect 104794 0 104850 800
rect 105254 0 105310 800
rect 105806 0 105862 800
rect 106266 0 106322 800
rect 106726 0 106782 800
rect 107278 0 107334 800
rect 107738 0 107794 800
rect 108198 0 108254 800
rect 108750 0 108806 800
rect 109210 0 109266 800
rect 109670 0 109726 800
rect 110222 0 110278 800
rect 110682 0 110738 800
rect 111142 0 111198 800
rect 111602 0 111658 800
rect 112154 0 112210 800
rect 112614 0 112670 800
rect 113074 0 113130 800
rect 113626 0 113682 800
rect 114086 0 114142 800
rect 114546 0 114602 800
rect 115098 0 115154 800
rect 115558 0 115614 800
rect 116018 0 116074 800
rect 116570 0 116626 800
rect 117030 0 117086 800
rect 117490 0 117546 800
rect 118042 0 118098 800
rect 118502 0 118558 800
rect 118962 0 119018 800
rect 119514 0 119570 800
rect 119974 0 120030 800
rect 120434 0 120490 800
rect 120986 0 121042 800
rect 121446 0 121502 800
rect 121906 0 121962 800
rect 122458 0 122514 800
rect 122918 0 122974 800
rect 123378 0 123434 800
rect 123930 0 123986 800
rect 124390 0 124446 800
rect 124850 0 124906 800
rect 125402 0 125458 800
rect 125862 0 125918 800
rect 126322 0 126378 800
rect 126874 0 126930 800
rect 127334 0 127390 800
rect 127794 0 127850 800
rect 128346 0 128402 800
rect 128806 0 128862 800
rect 129266 0 129322 800
rect 129726 0 129782 800
rect 130278 0 130334 800
rect 130738 0 130794 800
rect 131198 0 131254 800
rect 131750 0 131806 800
rect 132210 0 132266 800
rect 132670 0 132726 800
rect 133222 0 133278 800
rect 133682 0 133738 800
rect 134142 0 134198 800
rect 134694 0 134750 800
rect 135154 0 135210 800
rect 135614 0 135670 800
rect 136166 0 136222 800
rect 136626 0 136682 800
rect 137086 0 137142 800
rect 137638 0 137694 800
rect 138098 0 138154 800
rect 138558 0 138614 800
rect 139110 0 139166 800
rect 139570 0 139626 800
rect 140030 0 140086 800
rect 140582 0 140638 800
rect 141042 0 141098 800
rect 141502 0 141558 800
rect 142054 0 142110 800
rect 142514 0 142570 800
rect 142974 0 143030 800
rect 143526 0 143582 800
rect 143986 0 144042 800
rect 144446 0 144502 800
rect 144998 0 145054 800
rect 145458 0 145514 800
rect 145918 0 145974 800
rect 146470 0 146526 800
rect 146930 0 146986 800
rect 147390 0 147446 800
rect 147850 0 147906 800
rect 148402 0 148458 800
rect 148862 0 148918 800
rect 149322 0 149378 800
rect 149874 0 149930 800
rect 150334 0 150390 800
rect 150794 0 150850 800
rect 151346 0 151402 800
rect 151806 0 151862 800
rect 152266 0 152322 800
rect 152818 0 152874 800
rect 153278 0 153334 800
rect 153738 0 153794 800
rect 154290 0 154346 800
rect 154750 0 154806 800
rect 155210 0 155266 800
rect 155762 0 155818 800
rect 156222 0 156278 800
rect 156682 0 156738 800
rect 157234 0 157290 800
rect 157694 0 157750 800
rect 158154 0 158210 800
rect 158706 0 158762 800
rect 159166 0 159222 800
rect 159626 0 159682 800
rect 160178 0 160234 800
rect 160638 0 160694 800
rect 161098 0 161154 800
rect 161650 0 161706 800
rect 162110 0 162166 800
rect 162570 0 162626 800
rect 163122 0 163178 800
rect 163582 0 163638 800
rect 164042 0 164098 800
rect 164594 0 164650 800
rect 165054 0 165110 800
rect 165514 0 165570 800
rect 166066 0 166122 800
rect 166526 0 166582 800
rect 166986 0 167042 800
rect 167446 0 167502 800
rect 167998 0 168054 800
rect 168458 0 168514 800
rect 168918 0 168974 800
rect 169470 0 169526 800
rect 169930 0 169986 800
rect 170390 0 170446 800
rect 170942 0 170998 800
rect 171402 0 171458 800
rect 171862 0 171918 800
rect 172414 0 172470 800
rect 172874 0 172930 800
rect 173334 0 173390 800
rect 173886 0 173942 800
rect 174346 0 174402 800
rect 174806 0 174862 800
rect 175358 0 175414 800
rect 175818 0 175874 800
rect 176278 0 176334 800
rect 176830 0 176886 800
rect 177290 0 177346 800
rect 177750 0 177806 800
rect 178302 0 178358 800
rect 178762 0 178818 800
rect 179222 0 179278 800
rect 179774 0 179830 800
rect 180234 0 180290 800
rect 180694 0 180750 800
rect 181246 0 181302 800
rect 181706 0 181762 800
rect 182166 0 182222 800
rect 182718 0 182774 800
rect 183178 0 183234 800
rect 183638 0 183694 800
rect 184190 0 184246 800
rect 184650 0 184706 800
rect 185110 0 185166 800
rect 185570 0 185626 800
rect 186122 0 186178 800
rect 186582 0 186638 800
rect 187042 0 187098 800
rect 187594 0 187650 800
rect 188054 0 188110 800
rect 188514 0 188570 800
rect 189066 0 189122 800
rect 189526 0 189582 800
rect 189986 0 190042 800
rect 190538 0 190594 800
rect 190998 0 191054 800
rect 191458 0 191514 800
rect 192010 0 192066 800
rect 192470 0 192526 800
rect 192930 0 192986 800
rect 193482 0 193538 800
rect 193942 0 193998 800
rect 194402 0 194458 800
rect 194954 0 195010 800
rect 195414 0 195470 800
rect 195874 0 195930 800
rect 196426 0 196482 800
rect 196886 0 196942 800
rect 197346 0 197402 800
rect 197898 0 197954 800
rect 198358 0 198414 800
rect 198818 0 198874 800
rect 199370 0 199426 800
rect 199830 0 199886 800
rect 200290 0 200346 800
rect 200842 0 200898 800
rect 201302 0 201358 800
rect 201762 0 201818 800
rect 202314 0 202370 800
rect 202774 0 202830 800
rect 203234 0 203290 800
rect 203694 0 203750 800
rect 204246 0 204302 800
rect 204706 0 204762 800
rect 205166 0 205222 800
rect 205718 0 205774 800
rect 206178 0 206234 800
rect 206638 0 206694 800
rect 207190 0 207246 800
rect 207650 0 207706 800
rect 208110 0 208166 800
rect 208662 0 208718 800
rect 209122 0 209178 800
rect 209582 0 209638 800
rect 210134 0 210190 800
rect 210594 0 210650 800
rect 211054 0 211110 800
rect 211606 0 211662 800
rect 212066 0 212122 800
rect 212526 0 212582 800
rect 213078 0 213134 800
rect 213538 0 213594 800
rect 213998 0 214054 800
rect 214550 0 214606 800
rect 215010 0 215066 800
rect 215470 0 215526 800
rect 216022 0 216078 800
rect 216482 0 216538 800
rect 216942 0 216998 800
rect 217494 0 217550 800
rect 217954 0 218010 800
rect 218414 0 218470 800
rect 218966 0 219022 800
rect 219426 0 219482 800
rect 219886 0 219942 800
rect 220438 0 220494 800
rect 220898 0 220954 800
rect 221358 0 221414 800
rect 221818 0 221874 800
rect 222370 0 222426 800
rect 222830 0 222886 800
rect 223290 0 223346 800
rect 223842 0 223898 800
rect 224302 0 224358 800
rect 224762 0 224818 800
rect 225314 0 225370 800
rect 225774 0 225830 800
rect 226234 0 226290 800
rect 226786 0 226842 800
rect 227246 0 227302 800
rect 227706 0 227762 800
rect 228258 0 228314 800
rect 228718 0 228774 800
rect 229178 0 229234 800
rect 229730 0 229786 800
rect 230190 0 230246 800
rect 230650 0 230706 800
rect 231202 0 231258 800
rect 231662 0 231718 800
rect 232122 0 232178 800
rect 232674 0 232730 800
rect 233134 0 233190 800
rect 233594 0 233650 800
rect 234146 0 234202 800
rect 234606 0 234662 800
rect 235066 0 235122 800
rect 235618 0 235674 800
rect 236078 0 236134 800
rect 236538 0 236594 800
rect 237090 0 237146 800
rect 237550 0 237606 800
rect 238010 0 238066 800
rect 238562 0 238618 800
rect 239022 0 239078 800
rect 239482 0 239538 800
<< obsm2 >>
rect 6 239144 778 239200
rect 946 239144 2802 239200
rect 2970 239144 4918 239200
rect 5086 239144 7034 239200
rect 7202 239144 9150 239200
rect 9318 239144 11266 239200
rect 11434 239144 13382 239200
rect 13550 239144 15498 239200
rect 15666 239144 17614 239200
rect 17782 239144 19638 239200
rect 19806 239144 21754 239200
rect 21922 239144 23870 239200
rect 24038 239144 25986 239200
rect 26154 239144 28102 239200
rect 28270 239144 30218 239200
rect 30386 239144 32334 239200
rect 32502 239144 34450 239200
rect 34618 239144 36566 239200
rect 36734 239144 38590 239200
rect 38758 239144 40706 239200
rect 40874 239144 42822 239200
rect 42990 239144 44938 239200
rect 45106 239144 47054 239200
rect 47222 239144 49170 239200
rect 49338 239144 51286 239200
rect 51454 239144 53402 239200
rect 53570 239144 55518 239200
rect 55686 239144 57542 239200
rect 57710 239144 59658 239200
rect 59826 239144 61774 239200
rect 61942 239144 63890 239200
rect 64058 239144 66006 239200
rect 66174 239144 68122 239200
rect 68290 239144 70238 239200
rect 70406 239144 72354 239200
rect 72522 239144 74470 239200
rect 74638 239144 76494 239200
rect 76662 239144 78610 239200
rect 78778 239144 80726 239200
rect 80894 239144 82842 239200
rect 83010 239144 84958 239200
rect 85126 239144 87074 239200
rect 87242 239144 89190 239200
rect 89358 239144 91306 239200
rect 91474 239144 93330 239200
rect 93498 239144 95446 239200
rect 95614 239144 97562 239200
rect 97730 239144 99678 239200
rect 99846 239144 101794 239200
rect 101962 239144 103910 239200
rect 104078 239144 106026 239200
rect 106194 239144 108142 239200
rect 108310 239144 110258 239200
rect 110426 239144 112282 239200
rect 112450 239144 114398 239200
rect 114566 239144 116514 239200
rect 116682 239144 118630 239200
rect 118798 239144 120746 239200
rect 120914 239144 122862 239200
rect 123030 239144 124978 239200
rect 125146 239144 127094 239200
rect 127262 239144 129210 239200
rect 129378 239144 131234 239200
rect 131402 239144 133350 239200
rect 133518 239144 135466 239200
rect 135634 239144 137582 239200
rect 137750 239144 139698 239200
rect 139866 239144 141814 239200
rect 141982 239144 143930 239200
rect 144098 239144 146046 239200
rect 146214 239144 148162 239200
rect 148330 239144 150186 239200
rect 150354 239144 152302 239200
rect 152470 239144 154418 239200
rect 154586 239144 156534 239200
rect 156702 239144 158650 239200
rect 158818 239144 160766 239200
rect 160934 239144 162882 239200
rect 163050 239144 164998 239200
rect 165166 239144 167022 239200
rect 167190 239144 169138 239200
rect 169306 239144 171254 239200
rect 171422 239144 173370 239200
rect 173538 239144 175486 239200
rect 175654 239144 177602 239200
rect 177770 239144 179718 239200
rect 179886 239144 181834 239200
rect 182002 239144 183950 239200
rect 184118 239144 185974 239200
rect 186142 239144 188090 239200
rect 188258 239144 190206 239200
rect 190374 239144 192322 239200
rect 192490 239144 194438 239200
rect 194606 239144 196554 239200
rect 196722 239144 198670 239200
rect 198838 239144 200786 239200
rect 200954 239144 202902 239200
rect 203070 239144 204926 239200
rect 205094 239144 207042 239200
rect 207210 239144 209158 239200
rect 209326 239144 211274 239200
rect 211442 239144 213390 239200
rect 213558 239144 215506 239200
rect 215674 239144 217622 239200
rect 217790 239144 219738 239200
rect 219906 239144 221854 239200
rect 222022 239144 223878 239200
rect 224046 239144 225994 239200
rect 226162 239144 228110 239200
rect 228278 239144 230226 239200
rect 230394 239144 232342 239200
rect 232510 239144 234458 239200
rect 234626 239144 236574 239200
rect 236742 239144 238690 239200
rect 238858 239144 239536 239200
rect 6 856 239536 239144
rect 118 800 410 856
rect 578 800 870 856
rect 1038 800 1330 856
rect 1498 800 1882 856
rect 2050 800 2342 856
rect 2510 800 2802 856
rect 2970 800 3354 856
rect 3522 800 3814 856
rect 3982 800 4274 856
rect 4442 800 4826 856
rect 4994 800 5286 856
rect 5454 800 5746 856
rect 5914 800 6298 856
rect 6466 800 6758 856
rect 6926 800 7218 856
rect 7386 800 7770 856
rect 7938 800 8230 856
rect 8398 800 8690 856
rect 8858 800 9242 856
rect 9410 800 9702 856
rect 9870 800 10162 856
rect 10330 800 10714 856
rect 10882 800 11174 856
rect 11342 800 11634 856
rect 11802 800 12186 856
rect 12354 800 12646 856
rect 12814 800 13106 856
rect 13274 800 13658 856
rect 13826 800 14118 856
rect 14286 800 14578 856
rect 14746 800 15130 856
rect 15298 800 15590 856
rect 15758 800 16050 856
rect 16218 800 16602 856
rect 16770 800 17062 856
rect 17230 800 17522 856
rect 17690 800 18074 856
rect 18242 800 18534 856
rect 18702 800 18994 856
rect 19162 800 19454 856
rect 19622 800 20006 856
rect 20174 800 20466 856
rect 20634 800 20926 856
rect 21094 800 21478 856
rect 21646 800 21938 856
rect 22106 800 22398 856
rect 22566 800 22950 856
rect 23118 800 23410 856
rect 23578 800 23870 856
rect 24038 800 24422 856
rect 24590 800 24882 856
rect 25050 800 25342 856
rect 25510 800 25894 856
rect 26062 800 26354 856
rect 26522 800 26814 856
rect 26982 800 27366 856
rect 27534 800 27826 856
rect 27994 800 28286 856
rect 28454 800 28838 856
rect 29006 800 29298 856
rect 29466 800 29758 856
rect 29926 800 30310 856
rect 30478 800 30770 856
rect 30938 800 31230 856
rect 31398 800 31782 856
rect 31950 800 32242 856
rect 32410 800 32702 856
rect 32870 800 33254 856
rect 33422 800 33714 856
rect 33882 800 34174 856
rect 34342 800 34726 856
rect 34894 800 35186 856
rect 35354 800 35646 856
rect 35814 800 36198 856
rect 36366 800 36658 856
rect 36826 800 37118 856
rect 37286 800 37578 856
rect 37746 800 38130 856
rect 38298 800 38590 856
rect 38758 800 39050 856
rect 39218 800 39602 856
rect 39770 800 40062 856
rect 40230 800 40522 856
rect 40690 800 41074 856
rect 41242 800 41534 856
rect 41702 800 41994 856
rect 42162 800 42546 856
rect 42714 800 43006 856
rect 43174 800 43466 856
rect 43634 800 44018 856
rect 44186 800 44478 856
rect 44646 800 44938 856
rect 45106 800 45490 856
rect 45658 800 45950 856
rect 46118 800 46410 856
rect 46578 800 46962 856
rect 47130 800 47422 856
rect 47590 800 47882 856
rect 48050 800 48434 856
rect 48602 800 48894 856
rect 49062 800 49354 856
rect 49522 800 49906 856
rect 50074 800 50366 856
rect 50534 800 50826 856
rect 50994 800 51378 856
rect 51546 800 51838 856
rect 52006 800 52298 856
rect 52466 800 52850 856
rect 53018 800 53310 856
rect 53478 800 53770 856
rect 53938 800 54322 856
rect 54490 800 54782 856
rect 54950 800 55242 856
rect 55410 800 55702 856
rect 55870 800 56254 856
rect 56422 800 56714 856
rect 56882 800 57174 856
rect 57342 800 57726 856
rect 57894 800 58186 856
rect 58354 800 58646 856
rect 58814 800 59198 856
rect 59366 800 59658 856
rect 59826 800 60118 856
rect 60286 800 60670 856
rect 60838 800 61130 856
rect 61298 800 61590 856
rect 61758 800 62142 856
rect 62310 800 62602 856
rect 62770 800 63062 856
rect 63230 800 63614 856
rect 63782 800 64074 856
rect 64242 800 64534 856
rect 64702 800 65086 856
rect 65254 800 65546 856
rect 65714 800 66006 856
rect 66174 800 66558 856
rect 66726 800 67018 856
rect 67186 800 67478 856
rect 67646 800 68030 856
rect 68198 800 68490 856
rect 68658 800 68950 856
rect 69118 800 69502 856
rect 69670 800 69962 856
rect 70130 800 70422 856
rect 70590 800 70974 856
rect 71142 800 71434 856
rect 71602 800 71894 856
rect 72062 800 72446 856
rect 72614 800 72906 856
rect 73074 800 73366 856
rect 73534 800 73826 856
rect 73994 800 74378 856
rect 74546 800 74838 856
rect 75006 800 75298 856
rect 75466 800 75850 856
rect 76018 800 76310 856
rect 76478 800 76770 856
rect 76938 800 77322 856
rect 77490 800 77782 856
rect 77950 800 78242 856
rect 78410 800 78794 856
rect 78962 800 79254 856
rect 79422 800 79714 856
rect 79882 800 80266 856
rect 80434 800 80726 856
rect 80894 800 81186 856
rect 81354 800 81738 856
rect 81906 800 82198 856
rect 82366 800 82658 856
rect 82826 800 83210 856
rect 83378 800 83670 856
rect 83838 800 84130 856
rect 84298 800 84682 856
rect 84850 800 85142 856
rect 85310 800 85602 856
rect 85770 800 86154 856
rect 86322 800 86614 856
rect 86782 800 87074 856
rect 87242 800 87626 856
rect 87794 800 88086 856
rect 88254 800 88546 856
rect 88714 800 89098 856
rect 89266 800 89558 856
rect 89726 800 90018 856
rect 90186 800 90570 856
rect 90738 800 91030 856
rect 91198 800 91490 856
rect 91658 800 92042 856
rect 92210 800 92502 856
rect 92670 800 92962 856
rect 93130 800 93422 856
rect 93590 800 93974 856
rect 94142 800 94434 856
rect 94602 800 94894 856
rect 95062 800 95446 856
rect 95614 800 95906 856
rect 96074 800 96366 856
rect 96534 800 96918 856
rect 97086 800 97378 856
rect 97546 800 97838 856
rect 98006 800 98390 856
rect 98558 800 98850 856
rect 99018 800 99310 856
rect 99478 800 99862 856
rect 100030 800 100322 856
rect 100490 800 100782 856
rect 100950 800 101334 856
rect 101502 800 101794 856
rect 101962 800 102254 856
rect 102422 800 102806 856
rect 102974 800 103266 856
rect 103434 800 103726 856
rect 103894 800 104278 856
rect 104446 800 104738 856
rect 104906 800 105198 856
rect 105366 800 105750 856
rect 105918 800 106210 856
rect 106378 800 106670 856
rect 106838 800 107222 856
rect 107390 800 107682 856
rect 107850 800 108142 856
rect 108310 800 108694 856
rect 108862 800 109154 856
rect 109322 800 109614 856
rect 109782 800 110166 856
rect 110334 800 110626 856
rect 110794 800 111086 856
rect 111254 800 111546 856
rect 111714 800 112098 856
rect 112266 800 112558 856
rect 112726 800 113018 856
rect 113186 800 113570 856
rect 113738 800 114030 856
rect 114198 800 114490 856
rect 114658 800 115042 856
rect 115210 800 115502 856
rect 115670 800 115962 856
rect 116130 800 116514 856
rect 116682 800 116974 856
rect 117142 800 117434 856
rect 117602 800 117986 856
rect 118154 800 118446 856
rect 118614 800 118906 856
rect 119074 800 119458 856
rect 119626 800 119918 856
rect 120086 800 120378 856
rect 120546 800 120930 856
rect 121098 800 121390 856
rect 121558 800 121850 856
rect 122018 800 122402 856
rect 122570 800 122862 856
rect 123030 800 123322 856
rect 123490 800 123874 856
rect 124042 800 124334 856
rect 124502 800 124794 856
rect 124962 800 125346 856
rect 125514 800 125806 856
rect 125974 800 126266 856
rect 126434 800 126818 856
rect 126986 800 127278 856
rect 127446 800 127738 856
rect 127906 800 128290 856
rect 128458 800 128750 856
rect 128918 800 129210 856
rect 129378 800 129670 856
rect 129838 800 130222 856
rect 130390 800 130682 856
rect 130850 800 131142 856
rect 131310 800 131694 856
rect 131862 800 132154 856
rect 132322 800 132614 856
rect 132782 800 133166 856
rect 133334 800 133626 856
rect 133794 800 134086 856
rect 134254 800 134638 856
rect 134806 800 135098 856
rect 135266 800 135558 856
rect 135726 800 136110 856
rect 136278 800 136570 856
rect 136738 800 137030 856
rect 137198 800 137582 856
rect 137750 800 138042 856
rect 138210 800 138502 856
rect 138670 800 139054 856
rect 139222 800 139514 856
rect 139682 800 139974 856
rect 140142 800 140526 856
rect 140694 800 140986 856
rect 141154 800 141446 856
rect 141614 800 141998 856
rect 142166 800 142458 856
rect 142626 800 142918 856
rect 143086 800 143470 856
rect 143638 800 143930 856
rect 144098 800 144390 856
rect 144558 800 144942 856
rect 145110 800 145402 856
rect 145570 800 145862 856
rect 146030 800 146414 856
rect 146582 800 146874 856
rect 147042 800 147334 856
rect 147502 800 147794 856
rect 147962 800 148346 856
rect 148514 800 148806 856
rect 148974 800 149266 856
rect 149434 800 149818 856
rect 149986 800 150278 856
rect 150446 800 150738 856
rect 150906 800 151290 856
rect 151458 800 151750 856
rect 151918 800 152210 856
rect 152378 800 152762 856
rect 152930 800 153222 856
rect 153390 800 153682 856
rect 153850 800 154234 856
rect 154402 800 154694 856
rect 154862 800 155154 856
rect 155322 800 155706 856
rect 155874 800 156166 856
rect 156334 800 156626 856
rect 156794 800 157178 856
rect 157346 800 157638 856
rect 157806 800 158098 856
rect 158266 800 158650 856
rect 158818 800 159110 856
rect 159278 800 159570 856
rect 159738 800 160122 856
rect 160290 800 160582 856
rect 160750 800 161042 856
rect 161210 800 161594 856
rect 161762 800 162054 856
rect 162222 800 162514 856
rect 162682 800 163066 856
rect 163234 800 163526 856
rect 163694 800 163986 856
rect 164154 800 164538 856
rect 164706 800 164998 856
rect 165166 800 165458 856
rect 165626 800 166010 856
rect 166178 800 166470 856
rect 166638 800 166930 856
rect 167098 800 167390 856
rect 167558 800 167942 856
rect 168110 800 168402 856
rect 168570 800 168862 856
rect 169030 800 169414 856
rect 169582 800 169874 856
rect 170042 800 170334 856
rect 170502 800 170886 856
rect 171054 800 171346 856
rect 171514 800 171806 856
rect 171974 800 172358 856
rect 172526 800 172818 856
rect 172986 800 173278 856
rect 173446 800 173830 856
rect 173998 800 174290 856
rect 174458 800 174750 856
rect 174918 800 175302 856
rect 175470 800 175762 856
rect 175930 800 176222 856
rect 176390 800 176774 856
rect 176942 800 177234 856
rect 177402 800 177694 856
rect 177862 800 178246 856
rect 178414 800 178706 856
rect 178874 800 179166 856
rect 179334 800 179718 856
rect 179886 800 180178 856
rect 180346 800 180638 856
rect 180806 800 181190 856
rect 181358 800 181650 856
rect 181818 800 182110 856
rect 182278 800 182662 856
rect 182830 800 183122 856
rect 183290 800 183582 856
rect 183750 800 184134 856
rect 184302 800 184594 856
rect 184762 800 185054 856
rect 185222 800 185514 856
rect 185682 800 186066 856
rect 186234 800 186526 856
rect 186694 800 186986 856
rect 187154 800 187538 856
rect 187706 800 187998 856
rect 188166 800 188458 856
rect 188626 800 189010 856
rect 189178 800 189470 856
rect 189638 800 189930 856
rect 190098 800 190482 856
rect 190650 800 190942 856
rect 191110 800 191402 856
rect 191570 800 191954 856
rect 192122 800 192414 856
rect 192582 800 192874 856
rect 193042 800 193426 856
rect 193594 800 193886 856
rect 194054 800 194346 856
rect 194514 800 194898 856
rect 195066 800 195358 856
rect 195526 800 195818 856
rect 195986 800 196370 856
rect 196538 800 196830 856
rect 196998 800 197290 856
rect 197458 800 197842 856
rect 198010 800 198302 856
rect 198470 800 198762 856
rect 198930 800 199314 856
rect 199482 800 199774 856
rect 199942 800 200234 856
rect 200402 800 200786 856
rect 200954 800 201246 856
rect 201414 800 201706 856
rect 201874 800 202258 856
rect 202426 800 202718 856
rect 202886 800 203178 856
rect 203346 800 203638 856
rect 203806 800 204190 856
rect 204358 800 204650 856
rect 204818 800 205110 856
rect 205278 800 205662 856
rect 205830 800 206122 856
rect 206290 800 206582 856
rect 206750 800 207134 856
rect 207302 800 207594 856
rect 207762 800 208054 856
rect 208222 800 208606 856
rect 208774 800 209066 856
rect 209234 800 209526 856
rect 209694 800 210078 856
rect 210246 800 210538 856
rect 210706 800 210998 856
rect 211166 800 211550 856
rect 211718 800 212010 856
rect 212178 800 212470 856
rect 212638 800 213022 856
rect 213190 800 213482 856
rect 213650 800 213942 856
rect 214110 800 214494 856
rect 214662 800 214954 856
rect 215122 800 215414 856
rect 215582 800 215966 856
rect 216134 800 216426 856
rect 216594 800 216886 856
rect 217054 800 217438 856
rect 217606 800 217898 856
rect 218066 800 218358 856
rect 218526 800 218910 856
rect 219078 800 219370 856
rect 219538 800 219830 856
rect 219998 800 220382 856
rect 220550 800 220842 856
rect 221010 800 221302 856
rect 221470 800 221762 856
rect 221930 800 222314 856
rect 222482 800 222774 856
rect 222942 800 223234 856
rect 223402 800 223786 856
rect 223954 800 224246 856
rect 224414 800 224706 856
rect 224874 800 225258 856
rect 225426 800 225718 856
rect 225886 800 226178 856
rect 226346 800 226730 856
rect 226898 800 227190 856
rect 227358 800 227650 856
rect 227818 800 228202 856
rect 228370 800 228662 856
rect 228830 800 229122 856
rect 229290 800 229674 856
rect 229842 800 230134 856
rect 230302 800 230594 856
rect 230762 800 231146 856
rect 231314 800 231606 856
rect 231774 800 232066 856
rect 232234 800 232618 856
rect 232786 800 233078 856
rect 233246 800 233538 856
rect 233706 800 234090 856
rect 234258 800 234550 856
rect 234718 800 235010 856
rect 235178 800 235562 856
rect 235730 800 236022 856
rect 236190 800 236482 856
rect 236650 800 237034 856
rect 237202 800 237494 856
rect 237662 800 237954 856
rect 238122 800 238506 856
rect 238674 800 238966 856
rect 239134 800 239426 856
<< obsm3 >>
rect 1 851 235587 237761
<< metal4 >>
rect 4012 2128 4332 237776
rect 19372 2128 19692 237776
<< obsm4 >>
rect 19183 2128 19292 237776
rect 19772 2128 234732 237776
<< labels >>
rlabel metal2 s 834 239200 890 240000 6 io_in[0]
port 1 nsew default input
rlabel metal2 s 63946 239200 64002 240000 6 io_in[10]
port 2 nsew default input
rlabel metal2 s 70294 239200 70350 240000 6 io_in[11]
port 3 nsew default input
rlabel metal2 s 76550 239200 76606 240000 6 io_in[12]
port 4 nsew default input
rlabel metal2 s 82898 239200 82954 240000 6 io_in[13]
port 5 nsew default input
rlabel metal2 s 89246 239200 89302 240000 6 io_in[14]
port 6 nsew default input
rlabel metal2 s 95502 239200 95558 240000 6 io_in[15]
port 7 nsew default input
rlabel metal2 s 101850 239200 101906 240000 6 io_in[16]
port 8 nsew default input
rlabel metal2 s 108198 239200 108254 240000 6 io_in[17]
port 9 nsew default input
rlabel metal2 s 114454 239200 114510 240000 6 io_in[18]
port 10 nsew default input
rlabel metal2 s 120802 239200 120858 240000 6 io_in[19]
port 11 nsew default input
rlabel metal2 s 7090 239200 7146 240000 6 io_in[1]
port 12 nsew default input
rlabel metal2 s 127150 239200 127206 240000 6 io_in[20]
port 13 nsew default input
rlabel metal2 s 133406 239200 133462 240000 6 io_in[21]
port 14 nsew default input
rlabel metal2 s 139754 239200 139810 240000 6 io_in[22]
port 15 nsew default input
rlabel metal2 s 146102 239200 146158 240000 6 io_in[23]
port 16 nsew default input
rlabel metal2 s 152358 239200 152414 240000 6 io_in[24]
port 17 nsew default input
rlabel metal2 s 158706 239200 158762 240000 6 io_in[25]
port 18 nsew default input
rlabel metal2 s 165054 239200 165110 240000 6 io_in[26]
port 19 nsew default input
rlabel metal2 s 171310 239200 171366 240000 6 io_in[27]
port 20 nsew default input
rlabel metal2 s 177658 239200 177714 240000 6 io_in[28]
port 21 nsew default input
rlabel metal2 s 184006 239200 184062 240000 6 io_in[29]
port 22 nsew default input
rlabel metal2 s 13438 239200 13494 240000 6 io_in[2]
port 23 nsew default input
rlabel metal2 s 190262 239200 190318 240000 6 io_in[30]
port 24 nsew default input
rlabel metal2 s 196610 239200 196666 240000 6 io_in[31]
port 25 nsew default input
rlabel metal2 s 202958 239200 203014 240000 6 io_in[32]
port 26 nsew default input
rlabel metal2 s 209214 239200 209270 240000 6 io_in[33]
port 27 nsew default input
rlabel metal2 s 215562 239200 215618 240000 6 io_in[34]
port 28 nsew default input
rlabel metal2 s 221910 239200 221966 240000 6 io_in[35]
port 29 nsew default input
rlabel metal2 s 228166 239200 228222 240000 6 io_in[36]
port 30 nsew default input
rlabel metal2 s 234514 239200 234570 240000 6 io_in[37]
port 31 nsew default input
rlabel metal2 s 19694 239200 19750 240000 6 io_in[3]
port 32 nsew default input
rlabel metal2 s 26042 239200 26098 240000 6 io_in[4]
port 33 nsew default input
rlabel metal2 s 32390 239200 32446 240000 6 io_in[5]
port 34 nsew default input
rlabel metal2 s 38646 239200 38702 240000 6 io_in[6]
port 35 nsew default input
rlabel metal2 s 44994 239200 45050 240000 6 io_in[7]
port 36 nsew default input
rlabel metal2 s 51342 239200 51398 240000 6 io_in[8]
port 37 nsew default input
rlabel metal2 s 57598 239200 57654 240000 6 io_in[9]
port 38 nsew default input
rlabel metal2 s 2858 239200 2914 240000 6 io_oeb[0]
port 39 nsew default output
rlabel metal2 s 66062 239200 66118 240000 6 io_oeb[10]
port 40 nsew default output
rlabel metal2 s 72410 239200 72466 240000 6 io_oeb[11]
port 41 nsew default output
rlabel metal2 s 78666 239200 78722 240000 6 io_oeb[12]
port 42 nsew default output
rlabel metal2 s 85014 239200 85070 240000 6 io_oeb[13]
port 43 nsew default output
rlabel metal2 s 91362 239200 91418 240000 6 io_oeb[14]
port 44 nsew default output
rlabel metal2 s 97618 239200 97674 240000 6 io_oeb[15]
port 45 nsew default output
rlabel metal2 s 103966 239200 104022 240000 6 io_oeb[16]
port 46 nsew default output
rlabel metal2 s 110314 239200 110370 240000 6 io_oeb[17]
port 47 nsew default output
rlabel metal2 s 116570 239200 116626 240000 6 io_oeb[18]
port 48 nsew default output
rlabel metal2 s 122918 239200 122974 240000 6 io_oeb[19]
port 49 nsew default output
rlabel metal2 s 9206 239200 9262 240000 6 io_oeb[1]
port 50 nsew default output
rlabel metal2 s 129266 239200 129322 240000 6 io_oeb[20]
port 51 nsew default output
rlabel metal2 s 135522 239200 135578 240000 6 io_oeb[21]
port 52 nsew default output
rlabel metal2 s 141870 239200 141926 240000 6 io_oeb[22]
port 53 nsew default output
rlabel metal2 s 148218 239200 148274 240000 6 io_oeb[23]
port 54 nsew default output
rlabel metal2 s 154474 239200 154530 240000 6 io_oeb[24]
port 55 nsew default output
rlabel metal2 s 160822 239200 160878 240000 6 io_oeb[25]
port 56 nsew default output
rlabel metal2 s 167078 239200 167134 240000 6 io_oeb[26]
port 57 nsew default output
rlabel metal2 s 173426 239200 173482 240000 6 io_oeb[27]
port 58 nsew default output
rlabel metal2 s 179774 239200 179830 240000 6 io_oeb[28]
port 59 nsew default output
rlabel metal2 s 186030 239200 186086 240000 6 io_oeb[29]
port 60 nsew default output
rlabel metal2 s 15554 239200 15610 240000 6 io_oeb[2]
port 61 nsew default output
rlabel metal2 s 192378 239200 192434 240000 6 io_oeb[30]
port 62 nsew default output
rlabel metal2 s 198726 239200 198782 240000 6 io_oeb[31]
port 63 nsew default output
rlabel metal2 s 204982 239200 205038 240000 6 io_oeb[32]
port 64 nsew default output
rlabel metal2 s 211330 239200 211386 240000 6 io_oeb[33]
port 65 nsew default output
rlabel metal2 s 217678 239200 217734 240000 6 io_oeb[34]
port 66 nsew default output
rlabel metal2 s 223934 239200 223990 240000 6 io_oeb[35]
port 67 nsew default output
rlabel metal2 s 230282 239200 230338 240000 6 io_oeb[36]
port 68 nsew default output
rlabel metal2 s 236630 239200 236686 240000 6 io_oeb[37]
port 69 nsew default output
rlabel metal2 s 21810 239200 21866 240000 6 io_oeb[3]
port 70 nsew default output
rlabel metal2 s 28158 239200 28214 240000 6 io_oeb[4]
port 71 nsew default output
rlabel metal2 s 34506 239200 34562 240000 6 io_oeb[5]
port 72 nsew default output
rlabel metal2 s 40762 239200 40818 240000 6 io_oeb[6]
port 73 nsew default output
rlabel metal2 s 47110 239200 47166 240000 6 io_oeb[7]
port 74 nsew default output
rlabel metal2 s 53458 239200 53514 240000 6 io_oeb[8]
port 75 nsew default output
rlabel metal2 s 59714 239200 59770 240000 6 io_oeb[9]
port 76 nsew default output
rlabel metal2 s 4974 239200 5030 240000 6 io_out[0]
port 77 nsew default output
rlabel metal2 s 68178 239200 68234 240000 6 io_out[10]
port 78 nsew default output
rlabel metal2 s 74526 239200 74582 240000 6 io_out[11]
port 79 nsew default output
rlabel metal2 s 80782 239200 80838 240000 6 io_out[12]
port 80 nsew default output
rlabel metal2 s 87130 239200 87186 240000 6 io_out[13]
port 81 nsew default output
rlabel metal2 s 93386 239200 93442 240000 6 io_out[14]
port 82 nsew default output
rlabel metal2 s 99734 239200 99790 240000 6 io_out[15]
port 83 nsew default output
rlabel metal2 s 106082 239200 106138 240000 6 io_out[16]
port 84 nsew default output
rlabel metal2 s 112338 239200 112394 240000 6 io_out[17]
port 85 nsew default output
rlabel metal2 s 118686 239200 118742 240000 6 io_out[18]
port 86 nsew default output
rlabel metal2 s 125034 239200 125090 240000 6 io_out[19]
port 87 nsew default output
rlabel metal2 s 11322 239200 11378 240000 6 io_out[1]
port 88 nsew default output
rlabel metal2 s 131290 239200 131346 240000 6 io_out[20]
port 89 nsew default output
rlabel metal2 s 137638 239200 137694 240000 6 io_out[21]
port 90 nsew default output
rlabel metal2 s 143986 239200 144042 240000 6 io_out[22]
port 91 nsew default output
rlabel metal2 s 150242 239200 150298 240000 6 io_out[23]
port 92 nsew default output
rlabel metal2 s 156590 239200 156646 240000 6 io_out[24]
port 93 nsew default output
rlabel metal2 s 162938 239200 162994 240000 6 io_out[25]
port 94 nsew default output
rlabel metal2 s 169194 239200 169250 240000 6 io_out[26]
port 95 nsew default output
rlabel metal2 s 175542 239200 175598 240000 6 io_out[27]
port 96 nsew default output
rlabel metal2 s 181890 239200 181946 240000 6 io_out[28]
port 97 nsew default output
rlabel metal2 s 188146 239200 188202 240000 6 io_out[29]
port 98 nsew default output
rlabel metal2 s 17670 239200 17726 240000 6 io_out[2]
port 99 nsew default output
rlabel metal2 s 194494 239200 194550 240000 6 io_out[30]
port 100 nsew default output
rlabel metal2 s 200842 239200 200898 240000 6 io_out[31]
port 101 nsew default output
rlabel metal2 s 207098 239200 207154 240000 6 io_out[32]
port 102 nsew default output
rlabel metal2 s 213446 239200 213502 240000 6 io_out[33]
port 103 nsew default output
rlabel metal2 s 219794 239200 219850 240000 6 io_out[34]
port 104 nsew default output
rlabel metal2 s 226050 239200 226106 240000 6 io_out[35]
port 105 nsew default output
rlabel metal2 s 232398 239200 232454 240000 6 io_out[36]
port 106 nsew default output
rlabel metal2 s 238746 239200 238802 240000 6 io_out[37]
port 107 nsew default output
rlabel metal2 s 23926 239200 23982 240000 6 io_out[3]
port 108 nsew default output
rlabel metal2 s 30274 239200 30330 240000 6 io_out[4]
port 109 nsew default output
rlabel metal2 s 36622 239200 36678 240000 6 io_out[5]
port 110 nsew default output
rlabel metal2 s 42878 239200 42934 240000 6 io_out[6]
port 111 nsew default output
rlabel metal2 s 49226 239200 49282 240000 6 io_out[7]
port 112 nsew default output
rlabel metal2 s 55574 239200 55630 240000 6 io_out[8]
port 113 nsew default output
rlabel metal2 s 61830 239200 61886 240000 6 io_out[9]
port 114 nsew default output
rlabel metal2 s 51894 0 51950 800 6 la_data_in[0]
port 115 nsew default input
rlabel metal2 s 198818 0 198874 800 6 la_data_in[100]
port 116 nsew default input
rlabel metal2 s 200290 0 200346 800 6 la_data_in[101]
port 117 nsew default input
rlabel metal2 s 201762 0 201818 800 6 la_data_in[102]
port 118 nsew default input
rlabel metal2 s 203234 0 203290 800 6 la_data_in[103]
port 119 nsew default input
rlabel metal2 s 204706 0 204762 800 6 la_data_in[104]
port 120 nsew default input
rlabel metal2 s 206178 0 206234 800 6 la_data_in[105]
port 121 nsew default input
rlabel metal2 s 207650 0 207706 800 6 la_data_in[106]
port 122 nsew default input
rlabel metal2 s 209122 0 209178 800 6 la_data_in[107]
port 123 nsew default input
rlabel metal2 s 210594 0 210650 800 6 la_data_in[108]
port 124 nsew default input
rlabel metal2 s 212066 0 212122 800 6 la_data_in[109]
port 125 nsew default input
rlabel metal2 s 66614 0 66670 800 6 la_data_in[10]
port 126 nsew default input
rlabel metal2 s 213538 0 213594 800 6 la_data_in[110]
port 127 nsew default input
rlabel metal2 s 215010 0 215066 800 6 la_data_in[111]
port 128 nsew default input
rlabel metal2 s 216482 0 216538 800 6 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 217954 0 218010 800 6 la_data_in[113]
port 130 nsew default input
rlabel metal2 s 219426 0 219482 800 6 la_data_in[114]
port 131 nsew default input
rlabel metal2 s 220898 0 220954 800 6 la_data_in[115]
port 132 nsew default input
rlabel metal2 s 222370 0 222426 800 6 la_data_in[116]
port 133 nsew default input
rlabel metal2 s 223842 0 223898 800 6 la_data_in[117]
port 134 nsew default input
rlabel metal2 s 225314 0 225370 800 6 la_data_in[118]
port 135 nsew default input
rlabel metal2 s 226786 0 226842 800 6 la_data_in[119]
port 136 nsew default input
rlabel metal2 s 68086 0 68142 800 6 la_data_in[11]
port 137 nsew default input
rlabel metal2 s 228258 0 228314 800 6 la_data_in[120]
port 138 nsew default input
rlabel metal2 s 229730 0 229786 800 6 la_data_in[121]
port 139 nsew default input
rlabel metal2 s 231202 0 231258 800 6 la_data_in[122]
port 140 nsew default input
rlabel metal2 s 232674 0 232730 800 6 la_data_in[123]
port 141 nsew default input
rlabel metal2 s 234146 0 234202 800 6 la_data_in[124]
port 142 nsew default input
rlabel metal2 s 235618 0 235674 800 6 la_data_in[125]
port 143 nsew default input
rlabel metal2 s 237090 0 237146 800 6 la_data_in[126]
port 144 nsew default input
rlabel metal2 s 238562 0 238618 800 6 la_data_in[127]
port 145 nsew default input
rlabel metal2 s 69558 0 69614 800 6 la_data_in[12]
port 146 nsew default input
rlabel metal2 s 71030 0 71086 800 6 la_data_in[13]
port 147 nsew default input
rlabel metal2 s 72502 0 72558 800 6 la_data_in[14]
port 148 nsew default input
rlabel metal2 s 73882 0 73938 800 6 la_data_in[15]
port 149 nsew default input
rlabel metal2 s 75354 0 75410 800 6 la_data_in[16]
port 150 nsew default input
rlabel metal2 s 76826 0 76882 800 6 la_data_in[17]
port 151 nsew default input
rlabel metal2 s 78298 0 78354 800 6 la_data_in[18]
port 152 nsew default input
rlabel metal2 s 79770 0 79826 800 6 la_data_in[19]
port 153 nsew default input
rlabel metal2 s 53366 0 53422 800 6 la_data_in[1]
port 154 nsew default input
rlabel metal2 s 81242 0 81298 800 6 la_data_in[20]
port 155 nsew default input
rlabel metal2 s 82714 0 82770 800 6 la_data_in[21]
port 156 nsew default input
rlabel metal2 s 84186 0 84242 800 6 la_data_in[22]
port 157 nsew default input
rlabel metal2 s 85658 0 85714 800 6 la_data_in[23]
port 158 nsew default input
rlabel metal2 s 87130 0 87186 800 6 la_data_in[24]
port 159 nsew default input
rlabel metal2 s 88602 0 88658 800 6 la_data_in[25]
port 160 nsew default input
rlabel metal2 s 90074 0 90130 800 6 la_data_in[26]
port 161 nsew default input
rlabel metal2 s 91546 0 91602 800 6 la_data_in[27]
port 162 nsew default input
rlabel metal2 s 93018 0 93074 800 6 la_data_in[28]
port 163 nsew default input
rlabel metal2 s 94490 0 94546 800 6 la_data_in[29]
port 164 nsew default input
rlabel metal2 s 54838 0 54894 800 6 la_data_in[2]
port 165 nsew default input
rlabel metal2 s 95962 0 96018 800 6 la_data_in[30]
port 166 nsew default input
rlabel metal2 s 97434 0 97490 800 6 la_data_in[31]
port 167 nsew default input
rlabel metal2 s 98906 0 98962 800 6 la_data_in[32]
port 168 nsew default input
rlabel metal2 s 100378 0 100434 800 6 la_data_in[33]
port 169 nsew default input
rlabel metal2 s 101850 0 101906 800 6 la_data_in[34]
port 170 nsew default input
rlabel metal2 s 103322 0 103378 800 6 la_data_in[35]
port 171 nsew default input
rlabel metal2 s 104794 0 104850 800 6 la_data_in[36]
port 172 nsew default input
rlabel metal2 s 106266 0 106322 800 6 la_data_in[37]
port 173 nsew default input
rlabel metal2 s 107738 0 107794 800 6 la_data_in[38]
port 174 nsew default input
rlabel metal2 s 109210 0 109266 800 6 la_data_in[39]
port 175 nsew default input
rlabel metal2 s 56310 0 56366 800 6 la_data_in[3]
port 176 nsew default input
rlabel metal2 s 110682 0 110738 800 6 la_data_in[40]
port 177 nsew default input
rlabel metal2 s 112154 0 112210 800 6 la_data_in[41]
port 178 nsew default input
rlabel metal2 s 113626 0 113682 800 6 la_data_in[42]
port 179 nsew default input
rlabel metal2 s 115098 0 115154 800 6 la_data_in[43]
port 180 nsew default input
rlabel metal2 s 116570 0 116626 800 6 la_data_in[44]
port 181 nsew default input
rlabel metal2 s 118042 0 118098 800 6 la_data_in[45]
port 182 nsew default input
rlabel metal2 s 119514 0 119570 800 6 la_data_in[46]
port 183 nsew default input
rlabel metal2 s 120986 0 121042 800 6 la_data_in[47]
port 184 nsew default input
rlabel metal2 s 122458 0 122514 800 6 la_data_in[48]
port 185 nsew default input
rlabel metal2 s 123930 0 123986 800 6 la_data_in[49]
port 186 nsew default input
rlabel metal2 s 57782 0 57838 800 6 la_data_in[4]
port 187 nsew default input
rlabel metal2 s 125402 0 125458 800 6 la_data_in[50]
port 188 nsew default input
rlabel metal2 s 126874 0 126930 800 6 la_data_in[51]
port 189 nsew default input
rlabel metal2 s 128346 0 128402 800 6 la_data_in[52]
port 190 nsew default input
rlabel metal2 s 129726 0 129782 800 6 la_data_in[53]
port 191 nsew default input
rlabel metal2 s 131198 0 131254 800 6 la_data_in[54]
port 192 nsew default input
rlabel metal2 s 132670 0 132726 800 6 la_data_in[55]
port 193 nsew default input
rlabel metal2 s 134142 0 134198 800 6 la_data_in[56]
port 194 nsew default input
rlabel metal2 s 135614 0 135670 800 6 la_data_in[57]
port 195 nsew default input
rlabel metal2 s 137086 0 137142 800 6 la_data_in[58]
port 196 nsew default input
rlabel metal2 s 138558 0 138614 800 6 la_data_in[59]
port 197 nsew default input
rlabel metal2 s 59254 0 59310 800 6 la_data_in[5]
port 198 nsew default input
rlabel metal2 s 140030 0 140086 800 6 la_data_in[60]
port 199 nsew default input
rlabel metal2 s 141502 0 141558 800 6 la_data_in[61]
port 200 nsew default input
rlabel metal2 s 142974 0 143030 800 6 la_data_in[62]
port 201 nsew default input
rlabel metal2 s 144446 0 144502 800 6 la_data_in[63]
port 202 nsew default input
rlabel metal2 s 145918 0 145974 800 6 la_data_in[64]
port 203 nsew default input
rlabel metal2 s 147390 0 147446 800 6 la_data_in[65]
port 204 nsew default input
rlabel metal2 s 148862 0 148918 800 6 la_data_in[66]
port 205 nsew default input
rlabel metal2 s 150334 0 150390 800 6 la_data_in[67]
port 206 nsew default input
rlabel metal2 s 151806 0 151862 800 6 la_data_in[68]
port 207 nsew default input
rlabel metal2 s 153278 0 153334 800 6 la_data_in[69]
port 208 nsew default input
rlabel metal2 s 60726 0 60782 800 6 la_data_in[6]
port 209 nsew default input
rlabel metal2 s 154750 0 154806 800 6 la_data_in[70]
port 210 nsew default input
rlabel metal2 s 156222 0 156278 800 6 la_data_in[71]
port 211 nsew default input
rlabel metal2 s 157694 0 157750 800 6 la_data_in[72]
port 212 nsew default input
rlabel metal2 s 159166 0 159222 800 6 la_data_in[73]
port 213 nsew default input
rlabel metal2 s 160638 0 160694 800 6 la_data_in[74]
port 214 nsew default input
rlabel metal2 s 162110 0 162166 800 6 la_data_in[75]
port 215 nsew default input
rlabel metal2 s 163582 0 163638 800 6 la_data_in[76]
port 216 nsew default input
rlabel metal2 s 165054 0 165110 800 6 la_data_in[77]
port 217 nsew default input
rlabel metal2 s 166526 0 166582 800 6 la_data_in[78]
port 218 nsew default input
rlabel metal2 s 167998 0 168054 800 6 la_data_in[79]
port 219 nsew default input
rlabel metal2 s 62198 0 62254 800 6 la_data_in[7]
port 220 nsew default input
rlabel metal2 s 169470 0 169526 800 6 la_data_in[80]
port 221 nsew default input
rlabel metal2 s 170942 0 170998 800 6 la_data_in[81]
port 222 nsew default input
rlabel metal2 s 172414 0 172470 800 6 la_data_in[82]
port 223 nsew default input
rlabel metal2 s 173886 0 173942 800 6 la_data_in[83]
port 224 nsew default input
rlabel metal2 s 175358 0 175414 800 6 la_data_in[84]
port 225 nsew default input
rlabel metal2 s 176830 0 176886 800 6 la_data_in[85]
port 226 nsew default input
rlabel metal2 s 178302 0 178358 800 6 la_data_in[86]
port 227 nsew default input
rlabel metal2 s 179774 0 179830 800 6 la_data_in[87]
port 228 nsew default input
rlabel metal2 s 181246 0 181302 800 6 la_data_in[88]
port 229 nsew default input
rlabel metal2 s 182718 0 182774 800 6 la_data_in[89]
port 230 nsew default input
rlabel metal2 s 63670 0 63726 800 6 la_data_in[8]
port 231 nsew default input
rlabel metal2 s 184190 0 184246 800 6 la_data_in[90]
port 232 nsew default input
rlabel metal2 s 185570 0 185626 800 6 la_data_in[91]
port 233 nsew default input
rlabel metal2 s 187042 0 187098 800 6 la_data_in[92]
port 234 nsew default input
rlabel metal2 s 188514 0 188570 800 6 la_data_in[93]
port 235 nsew default input
rlabel metal2 s 189986 0 190042 800 6 la_data_in[94]
port 236 nsew default input
rlabel metal2 s 191458 0 191514 800 6 la_data_in[95]
port 237 nsew default input
rlabel metal2 s 192930 0 192986 800 6 la_data_in[96]
port 238 nsew default input
rlabel metal2 s 194402 0 194458 800 6 la_data_in[97]
port 239 nsew default input
rlabel metal2 s 195874 0 195930 800 6 la_data_in[98]
port 240 nsew default input
rlabel metal2 s 197346 0 197402 800 6 la_data_in[99]
port 241 nsew default input
rlabel metal2 s 65142 0 65198 800 6 la_data_in[9]
port 242 nsew default input
rlabel metal2 s 52354 0 52410 800 6 la_data_out[0]
port 243 nsew default output
rlabel metal2 s 199370 0 199426 800 6 la_data_out[100]
port 244 nsew default output
rlabel metal2 s 200842 0 200898 800 6 la_data_out[101]
port 245 nsew default output
rlabel metal2 s 202314 0 202370 800 6 la_data_out[102]
port 246 nsew default output
rlabel metal2 s 203694 0 203750 800 6 la_data_out[103]
port 247 nsew default output
rlabel metal2 s 205166 0 205222 800 6 la_data_out[104]
port 248 nsew default output
rlabel metal2 s 206638 0 206694 800 6 la_data_out[105]
port 249 nsew default output
rlabel metal2 s 208110 0 208166 800 6 la_data_out[106]
port 250 nsew default output
rlabel metal2 s 209582 0 209638 800 6 la_data_out[107]
port 251 nsew default output
rlabel metal2 s 211054 0 211110 800 6 la_data_out[108]
port 252 nsew default output
rlabel metal2 s 212526 0 212582 800 6 la_data_out[109]
port 253 nsew default output
rlabel metal2 s 67074 0 67130 800 6 la_data_out[10]
port 254 nsew default output
rlabel metal2 s 213998 0 214054 800 6 la_data_out[110]
port 255 nsew default output
rlabel metal2 s 215470 0 215526 800 6 la_data_out[111]
port 256 nsew default output
rlabel metal2 s 216942 0 216998 800 6 la_data_out[112]
port 257 nsew default output
rlabel metal2 s 218414 0 218470 800 6 la_data_out[113]
port 258 nsew default output
rlabel metal2 s 219886 0 219942 800 6 la_data_out[114]
port 259 nsew default output
rlabel metal2 s 221358 0 221414 800 6 la_data_out[115]
port 260 nsew default output
rlabel metal2 s 222830 0 222886 800 6 la_data_out[116]
port 261 nsew default output
rlabel metal2 s 224302 0 224358 800 6 la_data_out[117]
port 262 nsew default output
rlabel metal2 s 225774 0 225830 800 6 la_data_out[118]
port 263 nsew default output
rlabel metal2 s 227246 0 227302 800 6 la_data_out[119]
port 264 nsew default output
rlabel metal2 s 68546 0 68602 800 6 la_data_out[11]
port 265 nsew default output
rlabel metal2 s 228718 0 228774 800 6 la_data_out[120]
port 266 nsew default output
rlabel metal2 s 230190 0 230246 800 6 la_data_out[121]
port 267 nsew default output
rlabel metal2 s 231662 0 231718 800 6 la_data_out[122]
port 268 nsew default output
rlabel metal2 s 233134 0 233190 800 6 la_data_out[123]
port 269 nsew default output
rlabel metal2 s 234606 0 234662 800 6 la_data_out[124]
port 270 nsew default output
rlabel metal2 s 236078 0 236134 800 6 la_data_out[125]
port 271 nsew default output
rlabel metal2 s 237550 0 237606 800 6 la_data_out[126]
port 272 nsew default output
rlabel metal2 s 239022 0 239078 800 6 la_data_out[127]
port 273 nsew default output
rlabel metal2 s 70018 0 70074 800 6 la_data_out[12]
port 274 nsew default output
rlabel metal2 s 71490 0 71546 800 6 la_data_out[13]
port 275 nsew default output
rlabel metal2 s 72962 0 73018 800 6 la_data_out[14]
port 276 nsew default output
rlabel metal2 s 74434 0 74490 800 6 la_data_out[15]
port 277 nsew default output
rlabel metal2 s 75906 0 75962 800 6 la_data_out[16]
port 278 nsew default output
rlabel metal2 s 77378 0 77434 800 6 la_data_out[17]
port 279 nsew default output
rlabel metal2 s 78850 0 78906 800 6 la_data_out[18]
port 280 nsew default output
rlabel metal2 s 80322 0 80378 800 6 la_data_out[19]
port 281 nsew default output
rlabel metal2 s 53826 0 53882 800 6 la_data_out[1]
port 282 nsew default output
rlabel metal2 s 81794 0 81850 800 6 la_data_out[20]
port 283 nsew default output
rlabel metal2 s 83266 0 83322 800 6 la_data_out[21]
port 284 nsew default output
rlabel metal2 s 84738 0 84794 800 6 la_data_out[22]
port 285 nsew default output
rlabel metal2 s 86210 0 86266 800 6 la_data_out[23]
port 286 nsew default output
rlabel metal2 s 87682 0 87738 800 6 la_data_out[24]
port 287 nsew default output
rlabel metal2 s 89154 0 89210 800 6 la_data_out[25]
port 288 nsew default output
rlabel metal2 s 90626 0 90682 800 6 la_data_out[26]
port 289 nsew default output
rlabel metal2 s 92098 0 92154 800 6 la_data_out[27]
port 290 nsew default output
rlabel metal2 s 93478 0 93534 800 6 la_data_out[28]
port 291 nsew default output
rlabel metal2 s 94950 0 95006 800 6 la_data_out[29]
port 292 nsew default output
rlabel metal2 s 55298 0 55354 800 6 la_data_out[2]
port 293 nsew default output
rlabel metal2 s 96422 0 96478 800 6 la_data_out[30]
port 294 nsew default output
rlabel metal2 s 97894 0 97950 800 6 la_data_out[31]
port 295 nsew default output
rlabel metal2 s 99366 0 99422 800 6 la_data_out[32]
port 296 nsew default output
rlabel metal2 s 100838 0 100894 800 6 la_data_out[33]
port 297 nsew default output
rlabel metal2 s 102310 0 102366 800 6 la_data_out[34]
port 298 nsew default output
rlabel metal2 s 103782 0 103838 800 6 la_data_out[35]
port 299 nsew default output
rlabel metal2 s 105254 0 105310 800 6 la_data_out[36]
port 300 nsew default output
rlabel metal2 s 106726 0 106782 800 6 la_data_out[37]
port 301 nsew default output
rlabel metal2 s 108198 0 108254 800 6 la_data_out[38]
port 302 nsew default output
rlabel metal2 s 109670 0 109726 800 6 la_data_out[39]
port 303 nsew default output
rlabel metal2 s 56770 0 56826 800 6 la_data_out[3]
port 304 nsew default output
rlabel metal2 s 111142 0 111198 800 6 la_data_out[40]
port 305 nsew default output
rlabel metal2 s 112614 0 112670 800 6 la_data_out[41]
port 306 nsew default output
rlabel metal2 s 114086 0 114142 800 6 la_data_out[42]
port 307 nsew default output
rlabel metal2 s 115558 0 115614 800 6 la_data_out[43]
port 308 nsew default output
rlabel metal2 s 117030 0 117086 800 6 la_data_out[44]
port 309 nsew default output
rlabel metal2 s 118502 0 118558 800 6 la_data_out[45]
port 310 nsew default output
rlabel metal2 s 119974 0 120030 800 6 la_data_out[46]
port 311 nsew default output
rlabel metal2 s 121446 0 121502 800 6 la_data_out[47]
port 312 nsew default output
rlabel metal2 s 122918 0 122974 800 6 la_data_out[48]
port 313 nsew default output
rlabel metal2 s 124390 0 124446 800 6 la_data_out[49]
port 314 nsew default output
rlabel metal2 s 58242 0 58298 800 6 la_data_out[4]
port 315 nsew default output
rlabel metal2 s 125862 0 125918 800 6 la_data_out[50]
port 316 nsew default output
rlabel metal2 s 127334 0 127390 800 6 la_data_out[51]
port 317 nsew default output
rlabel metal2 s 128806 0 128862 800 6 la_data_out[52]
port 318 nsew default output
rlabel metal2 s 130278 0 130334 800 6 la_data_out[53]
port 319 nsew default output
rlabel metal2 s 131750 0 131806 800 6 la_data_out[54]
port 320 nsew default output
rlabel metal2 s 133222 0 133278 800 6 la_data_out[55]
port 321 nsew default output
rlabel metal2 s 134694 0 134750 800 6 la_data_out[56]
port 322 nsew default output
rlabel metal2 s 136166 0 136222 800 6 la_data_out[57]
port 323 nsew default output
rlabel metal2 s 137638 0 137694 800 6 la_data_out[58]
port 324 nsew default output
rlabel metal2 s 139110 0 139166 800 6 la_data_out[59]
port 325 nsew default output
rlabel metal2 s 59714 0 59770 800 6 la_data_out[5]
port 326 nsew default output
rlabel metal2 s 140582 0 140638 800 6 la_data_out[60]
port 327 nsew default output
rlabel metal2 s 142054 0 142110 800 6 la_data_out[61]
port 328 nsew default output
rlabel metal2 s 143526 0 143582 800 6 la_data_out[62]
port 329 nsew default output
rlabel metal2 s 144998 0 145054 800 6 la_data_out[63]
port 330 nsew default output
rlabel metal2 s 146470 0 146526 800 6 la_data_out[64]
port 331 nsew default output
rlabel metal2 s 147850 0 147906 800 6 la_data_out[65]
port 332 nsew default output
rlabel metal2 s 149322 0 149378 800 6 la_data_out[66]
port 333 nsew default output
rlabel metal2 s 150794 0 150850 800 6 la_data_out[67]
port 334 nsew default output
rlabel metal2 s 152266 0 152322 800 6 la_data_out[68]
port 335 nsew default output
rlabel metal2 s 153738 0 153794 800 6 la_data_out[69]
port 336 nsew default output
rlabel metal2 s 61186 0 61242 800 6 la_data_out[6]
port 337 nsew default output
rlabel metal2 s 155210 0 155266 800 6 la_data_out[70]
port 338 nsew default output
rlabel metal2 s 156682 0 156738 800 6 la_data_out[71]
port 339 nsew default output
rlabel metal2 s 158154 0 158210 800 6 la_data_out[72]
port 340 nsew default output
rlabel metal2 s 159626 0 159682 800 6 la_data_out[73]
port 341 nsew default output
rlabel metal2 s 161098 0 161154 800 6 la_data_out[74]
port 342 nsew default output
rlabel metal2 s 162570 0 162626 800 6 la_data_out[75]
port 343 nsew default output
rlabel metal2 s 164042 0 164098 800 6 la_data_out[76]
port 344 nsew default output
rlabel metal2 s 165514 0 165570 800 6 la_data_out[77]
port 345 nsew default output
rlabel metal2 s 166986 0 167042 800 6 la_data_out[78]
port 346 nsew default output
rlabel metal2 s 168458 0 168514 800 6 la_data_out[79]
port 347 nsew default output
rlabel metal2 s 62658 0 62714 800 6 la_data_out[7]
port 348 nsew default output
rlabel metal2 s 169930 0 169986 800 6 la_data_out[80]
port 349 nsew default output
rlabel metal2 s 171402 0 171458 800 6 la_data_out[81]
port 350 nsew default output
rlabel metal2 s 172874 0 172930 800 6 la_data_out[82]
port 351 nsew default output
rlabel metal2 s 174346 0 174402 800 6 la_data_out[83]
port 352 nsew default output
rlabel metal2 s 175818 0 175874 800 6 la_data_out[84]
port 353 nsew default output
rlabel metal2 s 177290 0 177346 800 6 la_data_out[85]
port 354 nsew default output
rlabel metal2 s 178762 0 178818 800 6 la_data_out[86]
port 355 nsew default output
rlabel metal2 s 180234 0 180290 800 6 la_data_out[87]
port 356 nsew default output
rlabel metal2 s 181706 0 181762 800 6 la_data_out[88]
port 357 nsew default output
rlabel metal2 s 183178 0 183234 800 6 la_data_out[89]
port 358 nsew default output
rlabel metal2 s 64130 0 64186 800 6 la_data_out[8]
port 359 nsew default output
rlabel metal2 s 184650 0 184706 800 6 la_data_out[90]
port 360 nsew default output
rlabel metal2 s 186122 0 186178 800 6 la_data_out[91]
port 361 nsew default output
rlabel metal2 s 187594 0 187650 800 6 la_data_out[92]
port 362 nsew default output
rlabel metal2 s 189066 0 189122 800 6 la_data_out[93]
port 363 nsew default output
rlabel metal2 s 190538 0 190594 800 6 la_data_out[94]
port 364 nsew default output
rlabel metal2 s 192010 0 192066 800 6 la_data_out[95]
port 365 nsew default output
rlabel metal2 s 193482 0 193538 800 6 la_data_out[96]
port 366 nsew default output
rlabel metal2 s 194954 0 195010 800 6 la_data_out[97]
port 367 nsew default output
rlabel metal2 s 196426 0 196482 800 6 la_data_out[98]
port 368 nsew default output
rlabel metal2 s 197898 0 197954 800 6 la_data_out[99]
port 369 nsew default output
rlabel metal2 s 65602 0 65658 800 6 la_data_out[9]
port 370 nsew default output
rlabel metal2 s 52906 0 52962 800 6 la_oen[0]
port 371 nsew default input
rlabel metal2 s 199830 0 199886 800 6 la_oen[100]
port 372 nsew default input
rlabel metal2 s 201302 0 201358 800 6 la_oen[101]
port 373 nsew default input
rlabel metal2 s 202774 0 202830 800 6 la_oen[102]
port 374 nsew default input
rlabel metal2 s 204246 0 204302 800 6 la_oen[103]
port 375 nsew default input
rlabel metal2 s 205718 0 205774 800 6 la_oen[104]
port 376 nsew default input
rlabel metal2 s 207190 0 207246 800 6 la_oen[105]
port 377 nsew default input
rlabel metal2 s 208662 0 208718 800 6 la_oen[106]
port 378 nsew default input
rlabel metal2 s 210134 0 210190 800 6 la_oen[107]
port 379 nsew default input
rlabel metal2 s 211606 0 211662 800 6 la_oen[108]
port 380 nsew default input
rlabel metal2 s 213078 0 213134 800 6 la_oen[109]
port 381 nsew default input
rlabel metal2 s 67534 0 67590 800 6 la_oen[10]
port 382 nsew default input
rlabel metal2 s 214550 0 214606 800 6 la_oen[110]
port 383 nsew default input
rlabel metal2 s 216022 0 216078 800 6 la_oen[111]
port 384 nsew default input
rlabel metal2 s 217494 0 217550 800 6 la_oen[112]
port 385 nsew default input
rlabel metal2 s 218966 0 219022 800 6 la_oen[113]
port 386 nsew default input
rlabel metal2 s 220438 0 220494 800 6 la_oen[114]
port 387 nsew default input
rlabel metal2 s 221818 0 221874 800 6 la_oen[115]
port 388 nsew default input
rlabel metal2 s 223290 0 223346 800 6 la_oen[116]
port 389 nsew default input
rlabel metal2 s 224762 0 224818 800 6 la_oen[117]
port 390 nsew default input
rlabel metal2 s 226234 0 226290 800 6 la_oen[118]
port 391 nsew default input
rlabel metal2 s 227706 0 227762 800 6 la_oen[119]
port 392 nsew default input
rlabel metal2 s 69006 0 69062 800 6 la_oen[11]
port 393 nsew default input
rlabel metal2 s 229178 0 229234 800 6 la_oen[120]
port 394 nsew default input
rlabel metal2 s 230650 0 230706 800 6 la_oen[121]
port 395 nsew default input
rlabel metal2 s 232122 0 232178 800 6 la_oen[122]
port 396 nsew default input
rlabel metal2 s 233594 0 233650 800 6 la_oen[123]
port 397 nsew default input
rlabel metal2 s 235066 0 235122 800 6 la_oen[124]
port 398 nsew default input
rlabel metal2 s 236538 0 236594 800 6 la_oen[125]
port 399 nsew default input
rlabel metal2 s 238010 0 238066 800 6 la_oen[126]
port 400 nsew default input
rlabel metal2 s 239482 0 239538 800 6 la_oen[127]
port 401 nsew default input
rlabel metal2 s 70478 0 70534 800 6 la_oen[12]
port 402 nsew default input
rlabel metal2 s 71950 0 72006 800 6 la_oen[13]
port 403 nsew default input
rlabel metal2 s 73422 0 73478 800 6 la_oen[14]
port 404 nsew default input
rlabel metal2 s 74894 0 74950 800 6 la_oen[15]
port 405 nsew default input
rlabel metal2 s 76366 0 76422 800 6 la_oen[16]
port 406 nsew default input
rlabel metal2 s 77838 0 77894 800 6 la_oen[17]
port 407 nsew default input
rlabel metal2 s 79310 0 79366 800 6 la_oen[18]
port 408 nsew default input
rlabel metal2 s 80782 0 80838 800 6 la_oen[19]
port 409 nsew default input
rlabel metal2 s 54378 0 54434 800 6 la_oen[1]
port 410 nsew default input
rlabel metal2 s 82254 0 82310 800 6 la_oen[20]
port 411 nsew default input
rlabel metal2 s 83726 0 83782 800 6 la_oen[21]
port 412 nsew default input
rlabel metal2 s 85198 0 85254 800 6 la_oen[22]
port 413 nsew default input
rlabel metal2 s 86670 0 86726 800 6 la_oen[23]
port 414 nsew default input
rlabel metal2 s 88142 0 88198 800 6 la_oen[24]
port 415 nsew default input
rlabel metal2 s 89614 0 89670 800 6 la_oen[25]
port 416 nsew default input
rlabel metal2 s 91086 0 91142 800 6 la_oen[26]
port 417 nsew default input
rlabel metal2 s 92558 0 92614 800 6 la_oen[27]
port 418 nsew default input
rlabel metal2 s 94030 0 94086 800 6 la_oen[28]
port 419 nsew default input
rlabel metal2 s 95502 0 95558 800 6 la_oen[29]
port 420 nsew default input
rlabel metal2 s 55758 0 55814 800 6 la_oen[2]
port 421 nsew default input
rlabel metal2 s 96974 0 97030 800 6 la_oen[30]
port 422 nsew default input
rlabel metal2 s 98446 0 98502 800 6 la_oen[31]
port 423 nsew default input
rlabel metal2 s 99918 0 99974 800 6 la_oen[32]
port 424 nsew default input
rlabel metal2 s 101390 0 101446 800 6 la_oen[33]
port 425 nsew default input
rlabel metal2 s 102862 0 102918 800 6 la_oen[34]
port 426 nsew default input
rlabel metal2 s 104334 0 104390 800 6 la_oen[35]
port 427 nsew default input
rlabel metal2 s 105806 0 105862 800 6 la_oen[36]
port 428 nsew default input
rlabel metal2 s 107278 0 107334 800 6 la_oen[37]
port 429 nsew default input
rlabel metal2 s 108750 0 108806 800 6 la_oen[38]
port 430 nsew default input
rlabel metal2 s 110222 0 110278 800 6 la_oen[39]
port 431 nsew default input
rlabel metal2 s 57230 0 57286 800 6 la_oen[3]
port 432 nsew default input
rlabel metal2 s 111602 0 111658 800 6 la_oen[40]
port 433 nsew default input
rlabel metal2 s 113074 0 113130 800 6 la_oen[41]
port 434 nsew default input
rlabel metal2 s 114546 0 114602 800 6 la_oen[42]
port 435 nsew default input
rlabel metal2 s 116018 0 116074 800 6 la_oen[43]
port 436 nsew default input
rlabel metal2 s 117490 0 117546 800 6 la_oen[44]
port 437 nsew default input
rlabel metal2 s 118962 0 119018 800 6 la_oen[45]
port 438 nsew default input
rlabel metal2 s 120434 0 120490 800 6 la_oen[46]
port 439 nsew default input
rlabel metal2 s 121906 0 121962 800 6 la_oen[47]
port 440 nsew default input
rlabel metal2 s 123378 0 123434 800 6 la_oen[48]
port 441 nsew default input
rlabel metal2 s 124850 0 124906 800 6 la_oen[49]
port 442 nsew default input
rlabel metal2 s 58702 0 58758 800 6 la_oen[4]
port 443 nsew default input
rlabel metal2 s 126322 0 126378 800 6 la_oen[50]
port 444 nsew default input
rlabel metal2 s 127794 0 127850 800 6 la_oen[51]
port 445 nsew default input
rlabel metal2 s 129266 0 129322 800 6 la_oen[52]
port 446 nsew default input
rlabel metal2 s 130738 0 130794 800 6 la_oen[53]
port 447 nsew default input
rlabel metal2 s 132210 0 132266 800 6 la_oen[54]
port 448 nsew default input
rlabel metal2 s 133682 0 133738 800 6 la_oen[55]
port 449 nsew default input
rlabel metal2 s 135154 0 135210 800 6 la_oen[56]
port 450 nsew default input
rlabel metal2 s 136626 0 136682 800 6 la_oen[57]
port 451 nsew default input
rlabel metal2 s 138098 0 138154 800 6 la_oen[58]
port 452 nsew default input
rlabel metal2 s 139570 0 139626 800 6 la_oen[59]
port 453 nsew default input
rlabel metal2 s 60174 0 60230 800 6 la_oen[5]
port 454 nsew default input
rlabel metal2 s 141042 0 141098 800 6 la_oen[60]
port 455 nsew default input
rlabel metal2 s 142514 0 142570 800 6 la_oen[61]
port 456 nsew default input
rlabel metal2 s 143986 0 144042 800 6 la_oen[62]
port 457 nsew default input
rlabel metal2 s 145458 0 145514 800 6 la_oen[63]
port 458 nsew default input
rlabel metal2 s 146930 0 146986 800 6 la_oen[64]
port 459 nsew default input
rlabel metal2 s 148402 0 148458 800 6 la_oen[65]
port 460 nsew default input
rlabel metal2 s 149874 0 149930 800 6 la_oen[66]
port 461 nsew default input
rlabel metal2 s 151346 0 151402 800 6 la_oen[67]
port 462 nsew default input
rlabel metal2 s 152818 0 152874 800 6 la_oen[68]
port 463 nsew default input
rlabel metal2 s 154290 0 154346 800 6 la_oen[69]
port 464 nsew default input
rlabel metal2 s 61646 0 61702 800 6 la_oen[6]
port 465 nsew default input
rlabel metal2 s 155762 0 155818 800 6 la_oen[70]
port 466 nsew default input
rlabel metal2 s 157234 0 157290 800 6 la_oen[71]
port 467 nsew default input
rlabel metal2 s 158706 0 158762 800 6 la_oen[72]
port 468 nsew default input
rlabel metal2 s 160178 0 160234 800 6 la_oen[73]
port 469 nsew default input
rlabel metal2 s 161650 0 161706 800 6 la_oen[74]
port 470 nsew default input
rlabel metal2 s 163122 0 163178 800 6 la_oen[75]
port 471 nsew default input
rlabel metal2 s 164594 0 164650 800 6 la_oen[76]
port 472 nsew default input
rlabel metal2 s 166066 0 166122 800 6 la_oen[77]
port 473 nsew default input
rlabel metal2 s 167446 0 167502 800 6 la_oen[78]
port 474 nsew default input
rlabel metal2 s 168918 0 168974 800 6 la_oen[79]
port 475 nsew default input
rlabel metal2 s 63118 0 63174 800 6 la_oen[7]
port 476 nsew default input
rlabel metal2 s 170390 0 170446 800 6 la_oen[80]
port 477 nsew default input
rlabel metal2 s 171862 0 171918 800 6 la_oen[81]
port 478 nsew default input
rlabel metal2 s 173334 0 173390 800 6 la_oen[82]
port 479 nsew default input
rlabel metal2 s 174806 0 174862 800 6 la_oen[83]
port 480 nsew default input
rlabel metal2 s 176278 0 176334 800 6 la_oen[84]
port 481 nsew default input
rlabel metal2 s 177750 0 177806 800 6 la_oen[85]
port 482 nsew default input
rlabel metal2 s 179222 0 179278 800 6 la_oen[86]
port 483 nsew default input
rlabel metal2 s 180694 0 180750 800 6 la_oen[87]
port 484 nsew default input
rlabel metal2 s 182166 0 182222 800 6 la_oen[88]
port 485 nsew default input
rlabel metal2 s 183638 0 183694 800 6 la_oen[89]
port 486 nsew default input
rlabel metal2 s 64590 0 64646 800 6 la_oen[8]
port 487 nsew default input
rlabel metal2 s 185110 0 185166 800 6 la_oen[90]
port 488 nsew default input
rlabel metal2 s 186582 0 186638 800 6 la_oen[91]
port 489 nsew default input
rlabel metal2 s 188054 0 188110 800 6 la_oen[92]
port 490 nsew default input
rlabel metal2 s 189526 0 189582 800 6 la_oen[93]
port 491 nsew default input
rlabel metal2 s 190998 0 191054 800 6 la_oen[94]
port 492 nsew default input
rlabel metal2 s 192470 0 192526 800 6 la_oen[95]
port 493 nsew default input
rlabel metal2 s 193942 0 193998 800 6 la_oen[96]
port 494 nsew default input
rlabel metal2 s 195414 0 195470 800 6 la_oen[97]
port 495 nsew default input
rlabel metal2 s 196886 0 196942 800 6 la_oen[98]
port 496 nsew default input
rlabel metal2 s 198358 0 198414 800 6 la_oen[99]
port 497 nsew default input
rlabel metal2 s 66062 0 66118 800 6 la_oen[9]
port 498 nsew default input
rlabel metal2 s 6 0 62 800 6 wb_clk_i
port 499 nsew default input
rlabel metal2 s 466 0 522 800 6 wb_rst_i
port 500 nsew default input
rlabel metal2 s 926 0 982 800 6 wbs_ack_o
port 501 nsew default output
rlabel metal2 s 2858 0 2914 800 6 wbs_adr_i[0]
port 502 nsew default input
rlabel metal2 s 19510 0 19566 800 6 wbs_adr_i[10]
port 503 nsew default input
rlabel metal2 s 20982 0 21038 800 6 wbs_adr_i[11]
port 504 nsew default input
rlabel metal2 s 22454 0 22510 800 6 wbs_adr_i[12]
port 505 nsew default input
rlabel metal2 s 23926 0 23982 800 6 wbs_adr_i[13]
port 506 nsew default input
rlabel metal2 s 25398 0 25454 800 6 wbs_adr_i[14]
port 507 nsew default input
rlabel metal2 s 26870 0 26926 800 6 wbs_adr_i[15]
port 508 nsew default input
rlabel metal2 s 28342 0 28398 800 6 wbs_adr_i[16]
port 509 nsew default input
rlabel metal2 s 29814 0 29870 800 6 wbs_adr_i[17]
port 510 nsew default input
rlabel metal2 s 31286 0 31342 800 6 wbs_adr_i[18]
port 511 nsew default input
rlabel metal2 s 32758 0 32814 800 6 wbs_adr_i[19]
port 512 nsew default input
rlabel metal2 s 4882 0 4938 800 6 wbs_adr_i[1]
port 513 nsew default input
rlabel metal2 s 34230 0 34286 800 6 wbs_adr_i[20]
port 514 nsew default input
rlabel metal2 s 35702 0 35758 800 6 wbs_adr_i[21]
port 515 nsew default input
rlabel metal2 s 37174 0 37230 800 6 wbs_adr_i[22]
port 516 nsew default input
rlabel metal2 s 38646 0 38702 800 6 wbs_adr_i[23]
port 517 nsew default input
rlabel metal2 s 40118 0 40174 800 6 wbs_adr_i[24]
port 518 nsew default input
rlabel metal2 s 41590 0 41646 800 6 wbs_adr_i[25]
port 519 nsew default input
rlabel metal2 s 43062 0 43118 800 6 wbs_adr_i[26]
port 520 nsew default input
rlabel metal2 s 44534 0 44590 800 6 wbs_adr_i[27]
port 521 nsew default input
rlabel metal2 s 46006 0 46062 800 6 wbs_adr_i[28]
port 522 nsew default input
rlabel metal2 s 47478 0 47534 800 6 wbs_adr_i[29]
port 523 nsew default input
rlabel metal2 s 6814 0 6870 800 6 wbs_adr_i[2]
port 524 nsew default input
rlabel metal2 s 48950 0 49006 800 6 wbs_adr_i[30]
port 525 nsew default input
rlabel metal2 s 50422 0 50478 800 6 wbs_adr_i[31]
port 526 nsew default input
rlabel metal2 s 8746 0 8802 800 6 wbs_adr_i[3]
port 527 nsew default input
rlabel metal2 s 10770 0 10826 800 6 wbs_adr_i[4]
port 528 nsew default input
rlabel metal2 s 12242 0 12298 800 6 wbs_adr_i[5]
port 529 nsew default input
rlabel metal2 s 13714 0 13770 800 6 wbs_adr_i[6]
port 530 nsew default input
rlabel metal2 s 15186 0 15242 800 6 wbs_adr_i[7]
port 531 nsew default input
rlabel metal2 s 16658 0 16714 800 6 wbs_adr_i[8]
port 532 nsew default input
rlabel metal2 s 18130 0 18186 800 6 wbs_adr_i[9]
port 533 nsew default input
rlabel metal2 s 1386 0 1442 800 6 wbs_cyc_i
port 534 nsew default input
rlabel metal2 s 3410 0 3466 800 6 wbs_dat_i[0]
port 535 nsew default input
rlabel metal2 s 20062 0 20118 800 6 wbs_dat_i[10]
port 536 nsew default input
rlabel metal2 s 21534 0 21590 800 6 wbs_dat_i[11]
port 537 nsew default input
rlabel metal2 s 23006 0 23062 800 6 wbs_dat_i[12]
port 538 nsew default input
rlabel metal2 s 24478 0 24534 800 6 wbs_dat_i[13]
port 539 nsew default input
rlabel metal2 s 25950 0 26006 800 6 wbs_dat_i[14]
port 540 nsew default input
rlabel metal2 s 27422 0 27478 800 6 wbs_dat_i[15]
port 541 nsew default input
rlabel metal2 s 28894 0 28950 800 6 wbs_dat_i[16]
port 542 nsew default input
rlabel metal2 s 30366 0 30422 800 6 wbs_dat_i[17]
port 543 nsew default input
rlabel metal2 s 31838 0 31894 800 6 wbs_dat_i[18]
port 544 nsew default input
rlabel metal2 s 33310 0 33366 800 6 wbs_dat_i[19]
port 545 nsew default input
rlabel metal2 s 5342 0 5398 800 6 wbs_dat_i[1]
port 546 nsew default input
rlabel metal2 s 34782 0 34838 800 6 wbs_dat_i[20]
port 547 nsew default input
rlabel metal2 s 36254 0 36310 800 6 wbs_dat_i[21]
port 548 nsew default input
rlabel metal2 s 37634 0 37690 800 6 wbs_dat_i[22]
port 549 nsew default input
rlabel metal2 s 39106 0 39162 800 6 wbs_dat_i[23]
port 550 nsew default input
rlabel metal2 s 40578 0 40634 800 6 wbs_dat_i[24]
port 551 nsew default input
rlabel metal2 s 42050 0 42106 800 6 wbs_dat_i[25]
port 552 nsew default input
rlabel metal2 s 43522 0 43578 800 6 wbs_dat_i[26]
port 553 nsew default input
rlabel metal2 s 44994 0 45050 800 6 wbs_dat_i[27]
port 554 nsew default input
rlabel metal2 s 46466 0 46522 800 6 wbs_dat_i[28]
port 555 nsew default input
rlabel metal2 s 47938 0 47994 800 6 wbs_dat_i[29]
port 556 nsew default input
rlabel metal2 s 7274 0 7330 800 6 wbs_dat_i[2]
port 557 nsew default input
rlabel metal2 s 49410 0 49466 800 6 wbs_dat_i[30]
port 558 nsew default input
rlabel metal2 s 50882 0 50938 800 6 wbs_dat_i[31]
port 559 nsew default input
rlabel metal2 s 9298 0 9354 800 6 wbs_dat_i[3]
port 560 nsew default input
rlabel metal2 s 11230 0 11286 800 6 wbs_dat_i[4]
port 561 nsew default input
rlabel metal2 s 12702 0 12758 800 6 wbs_dat_i[5]
port 562 nsew default input
rlabel metal2 s 14174 0 14230 800 6 wbs_dat_i[6]
port 563 nsew default input
rlabel metal2 s 15646 0 15702 800 6 wbs_dat_i[7]
port 564 nsew default input
rlabel metal2 s 17118 0 17174 800 6 wbs_dat_i[8]
port 565 nsew default input
rlabel metal2 s 18590 0 18646 800 6 wbs_dat_i[9]
port 566 nsew default input
rlabel metal2 s 3870 0 3926 800 6 wbs_dat_o[0]
port 567 nsew default output
rlabel metal2 s 20522 0 20578 800 6 wbs_dat_o[10]
port 568 nsew default output
rlabel metal2 s 21994 0 22050 800 6 wbs_dat_o[11]
port 569 nsew default output
rlabel metal2 s 23466 0 23522 800 6 wbs_dat_o[12]
port 570 nsew default output
rlabel metal2 s 24938 0 24994 800 6 wbs_dat_o[13]
port 571 nsew default output
rlabel metal2 s 26410 0 26466 800 6 wbs_dat_o[14]
port 572 nsew default output
rlabel metal2 s 27882 0 27938 800 6 wbs_dat_o[15]
port 573 nsew default output
rlabel metal2 s 29354 0 29410 800 6 wbs_dat_o[16]
port 574 nsew default output
rlabel metal2 s 30826 0 30882 800 6 wbs_dat_o[17]
port 575 nsew default output
rlabel metal2 s 32298 0 32354 800 6 wbs_dat_o[18]
port 576 nsew default output
rlabel metal2 s 33770 0 33826 800 6 wbs_dat_o[19]
port 577 nsew default output
rlabel metal2 s 5802 0 5858 800 6 wbs_dat_o[1]
port 578 nsew default output
rlabel metal2 s 35242 0 35298 800 6 wbs_dat_o[20]
port 579 nsew default output
rlabel metal2 s 36714 0 36770 800 6 wbs_dat_o[21]
port 580 nsew default output
rlabel metal2 s 38186 0 38242 800 6 wbs_dat_o[22]
port 581 nsew default output
rlabel metal2 s 39658 0 39714 800 6 wbs_dat_o[23]
port 582 nsew default output
rlabel metal2 s 41130 0 41186 800 6 wbs_dat_o[24]
port 583 nsew default output
rlabel metal2 s 42602 0 42658 800 6 wbs_dat_o[25]
port 584 nsew default output
rlabel metal2 s 44074 0 44130 800 6 wbs_dat_o[26]
port 585 nsew default output
rlabel metal2 s 45546 0 45602 800 6 wbs_dat_o[27]
port 586 nsew default output
rlabel metal2 s 47018 0 47074 800 6 wbs_dat_o[28]
port 587 nsew default output
rlabel metal2 s 48490 0 48546 800 6 wbs_dat_o[29]
port 588 nsew default output
rlabel metal2 s 7826 0 7882 800 6 wbs_dat_o[2]
port 589 nsew default output
rlabel metal2 s 49962 0 50018 800 6 wbs_dat_o[30]
port 590 nsew default output
rlabel metal2 s 51434 0 51490 800 6 wbs_dat_o[31]
port 591 nsew default output
rlabel metal2 s 9758 0 9814 800 6 wbs_dat_o[3]
port 592 nsew default output
rlabel metal2 s 11690 0 11746 800 6 wbs_dat_o[4]
port 593 nsew default output
rlabel metal2 s 13162 0 13218 800 6 wbs_dat_o[5]
port 594 nsew default output
rlabel metal2 s 14634 0 14690 800 6 wbs_dat_o[6]
port 595 nsew default output
rlabel metal2 s 16106 0 16162 800 6 wbs_dat_o[7]
port 596 nsew default output
rlabel metal2 s 17578 0 17634 800 6 wbs_dat_o[8]
port 597 nsew default output
rlabel metal2 s 19050 0 19106 800 6 wbs_dat_o[9]
port 598 nsew default output
rlabel metal2 s 4330 0 4386 800 6 wbs_sel_i[0]
port 599 nsew default input
rlabel metal2 s 6354 0 6410 800 6 wbs_sel_i[1]
port 600 nsew default input
rlabel metal2 s 8286 0 8342 800 6 wbs_sel_i[2]
port 601 nsew default input
rlabel metal2 s 10218 0 10274 800 6 wbs_sel_i[3]
port 602 nsew default input
rlabel metal2 s 1938 0 1994 800 6 wbs_stb_i
port 603 nsew default input
rlabel metal2 s 2398 0 2454 800 6 wbs_we_i
port 604 nsew default input
rlabel metal4 s 4012 2128 4332 237776 6 VPWR
port 605 nsew power input
rlabel metal4 s 19372 2128 19692 237776 6 VGND
port 606 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 1 0 239542 240000
string LEFview TRUE
<< end >>
