magic
tech sky130A
magscale 1 2
timestamp 1608158347
<< locali >>
rect 364533 676243 364567 685797
rect 429577 666587 429611 684437
rect 494069 666587 494103 676141
rect 559297 666587 559331 684437
rect 364533 608651 364567 618205
rect 429393 601715 429427 608549
rect 559113 601715 559147 608549
rect 364625 589339 364659 598893
rect 429577 589339 429611 598893
rect 559297 589339 559331 598893
rect 289737 579479 289771 579581
rect 289921 579479 289955 579513
rect 454049 579479 454083 579581
rect 289863 579445 289955 579479
rect 318809 579343 318843 579445
rect 252109 578595 252143 579309
rect 254225 578663 254259 579309
rect 294613 579003 294647 579309
rect 299305 579003 299339 579309
rect 312001 579275 312035 579309
rect 311851 579241 312035 579275
rect 328377 579275 328411 579445
rect 338129 579343 338163 579445
rect 331321 579275 331355 579309
rect 331171 579241 331355 579275
rect 347697 579275 347731 579445
rect 357449 579343 357483 579445
rect 350641 579275 350675 579309
rect 350491 579241 350675 579275
rect 367017 579275 367051 579445
rect 376769 579343 376803 579445
rect 369961 579275 369995 579309
rect 369811 579241 369995 579275
rect 386337 579275 386371 579445
rect 396089 579343 396123 579445
rect 389281 579275 389315 579309
rect 389131 579241 389315 579275
rect 405657 579275 405691 579445
rect 408509 579275 408543 579445
rect 415317 579343 415351 579445
rect 299155 578833 299397 578867
rect 299247 578765 299305 578799
rect 299155 578629 299305 578663
rect 299063 578561 299213 578595
rect 415685 578527 415719 579377
rect 298971 578493 299121 578527
rect 428381 578459 428415 579377
rect 441077 578391 441111 579309
rect 444297 579275 444331 579445
rect 444389 579275 444423 579445
rect 453589 578323 453623 579377
rect 455797 578255 455831 579377
rect 463617 579343 463651 579581
rect 464445 577915 464479 579309
rect 260481 337399 260515 337569
rect 86969 336991 87003 337093
rect 103437 336991 103471 337229
rect 113189 336787 113223 337229
rect 122757 336787 122791 337229
rect 284401 335223 284435 338045
rect 379471 338045 379529 338079
rect 302249 337195 302283 337773
rect 316693 337331 316727 338045
rect 250177 328491 250211 334441
rect 302525 328491 302559 334713
rect 321845 329171 321879 337229
rect 335829 336787 335863 337501
rect 335921 337467 335955 337841
rect 336013 337671 336047 337841
rect 344293 337637 344661 337671
rect 344293 337535 344327 337637
rect 335921 337433 336105 337467
rect 341717 336719 341751 337161
rect 342821 337127 342855 337501
rect 345673 336787 345707 337569
rect 348985 337467 349019 337705
rect 347789 337331 347823 337433
rect 360117 337331 360151 337705
rect 364349 337399 364383 337705
rect 364475 337501 364717 337535
rect 364993 337127 365027 337637
rect 365729 337603 365763 337841
rect 412557 337807 412591 337977
rect 451197 337807 451231 337977
rect 460581 337943 460615 338113
rect 412465 337671 412499 337773
rect 413971 337637 414305 337671
rect 369869 337195 369903 337365
rect 374653 337195 374687 337433
rect 412649 337331 412683 337569
rect 431877 337195 431911 337501
rect 345857 336991 345891 337093
rect 345615 336753 345707 336787
rect 432245 336991 432279 337705
rect 451105 337671 451139 337773
rect 443469 337399 443503 337637
rect 451289 337535 451323 337773
rect 345765 336787 345799 336957
rect 454693 336787 454727 337909
rect 461593 337603 461627 337977
rect 456993 337331 457027 337569
rect 460397 337263 460431 337569
rect 457177 336787 457211 337229
rect 461593 336855 461627 337297
rect 466285 336719 466319 337977
rect 466377 337807 466411 338113
rect 466469 336923 466503 337297
rect 469229 337263 469263 337909
rect 259837 318835 259871 328389
rect 330217 327199 330251 336685
rect 331413 327131 331447 336073
rect 341717 328491 341751 335529
rect 374469 327131 374503 336685
rect 375849 327131 375883 336685
rect 337209 320875 337243 321589
rect 341441 318835 341475 321589
rect 230857 309179 230891 318733
rect 236285 309247 236319 318733
rect 239229 309179 239263 318733
rect 244473 309179 244507 311797
rect 236285 299591 236319 309077
rect 259653 299591 259687 309077
rect 236285 289867 236319 299421
rect 262597 298231 262631 315945
rect 284677 314211 284711 318733
rect 357449 317475 357483 327029
rect 360393 317475 360427 327029
rect 389557 318835 389591 328389
rect 470609 318835 470643 328389
rect 273453 311899 273487 313429
rect 299765 299523 299799 317373
rect 310897 307887 310931 311933
rect 325893 307819 325927 317373
rect 337209 311763 337243 317373
rect 310713 298163 310747 307717
rect 239229 289867 239263 292553
rect 251465 289867 251499 294661
rect 236285 280279 236319 289697
rect 244473 280211 244507 289765
rect 266737 288439 266771 298061
rect 267749 288439 267783 298061
rect 270785 285651 270819 292485
rect 285965 288439 285999 298061
rect 294245 287079 294279 289833
rect 310897 282795 310931 293029
rect 323317 288439 323351 299421
rect 324697 289867 324731 299421
rect 327181 298163 327215 307717
rect 337209 298163 337243 307717
rect 341165 299523 341199 309077
rect 357817 299523 357851 309077
rect 358737 299523 358771 309077
rect 375849 307819 375883 317373
rect 327181 283611 327215 289765
rect 236285 270555 236319 280109
rect 239137 270555 239171 280109
rect 251465 270555 251499 280109
rect 259561 273071 259595 280109
rect 323501 278783 323535 283577
rect 236285 260967 236319 270385
rect 236285 251243 236319 260797
rect 239137 251243 239171 260797
rect 250085 259471 250119 269025
rect 310897 263483 310931 278681
rect 330125 269127 330159 273853
rect 331413 270555 331447 280109
rect 337209 276063 337243 285617
rect 341165 280211 341199 282897
rect 357449 280211 357483 289765
rect 358737 288439 358771 298061
rect 372721 289867 372755 299421
rect 374377 289867 374411 307717
rect 389281 299523 389315 309009
rect 470609 299523 470643 309077
rect 375849 289867 375883 299421
rect 389373 280211 389407 289765
rect 470609 280211 470643 289765
rect 338865 270555 338899 280109
rect 372721 270555 372755 280109
rect 377137 270555 377171 280109
rect 389373 260899 389407 270453
rect 470609 260899 470643 270453
rect 250177 251107 250211 259301
rect 251465 251243 251499 260797
rect 259561 253759 259595 260797
rect 262597 259471 262631 260865
rect 259561 244171 259595 251141
rect 270693 251107 270727 260797
rect 306757 248387 306791 258009
rect 310897 251311 310931 256037
rect 272165 241587 272199 244409
rect 266737 230503 266771 234821
rect 267749 231795 267783 240057
rect 272165 234515 272199 240057
rect 285965 234515 285999 244953
rect 310713 241519 310747 251141
rect 337117 247163 337151 253997
rect 338865 251243 338899 260797
rect 341073 253759 341107 260797
rect 357541 249815 357575 259369
rect 372721 251243 372755 260797
rect 377137 251243 377171 260797
rect 463709 251243 463743 260797
rect 337117 244239 337151 246993
rect 470609 241519 470643 251141
rect 290381 230435 290415 238697
rect 295625 229143 295659 238697
rect 299489 231863 299523 241417
rect 306941 230503 306975 238765
rect 331413 231863 331447 241417
rect 389281 234651 389315 241417
rect 270693 220847 270727 224961
rect 310805 222207 310839 231761
rect 290197 212483 290231 219385
rect 291669 212483 291703 219385
rect 299489 212551 299523 222105
rect 337117 220847 337151 231625
rect 341073 222207 341107 224961
rect 270693 202895 270727 205649
rect 302617 202895 302651 207757
rect 310805 202895 310839 212449
rect 250085 186303 250119 200073
rect 267749 183583 267783 186337
rect 270693 183583 270727 186337
rect 232329 172567 232363 182121
rect 259653 173995 259687 179537
rect 232237 164203 232271 172465
rect 265265 161483 265299 179333
rect 284769 171139 284803 180761
rect 288725 179435 288759 188989
rect 299857 180863 299891 190417
rect 302525 180863 302559 190417
rect 306849 180863 306883 190417
rect 339785 183583 339819 188377
rect 367017 183583 367051 193137
rect 267841 162775 267875 171037
rect 294429 161483 294463 171037
rect 337117 164203 337151 172465
rect 341257 169779 341291 179333
rect 358737 173859 358771 181985
rect 366925 173927 366959 174029
rect 259653 145027 259687 154173
rect 267841 151827 267875 161381
rect 250269 133943 250303 143497
rect 264989 142171 265023 151725
rect 291485 149107 291519 160021
rect 294429 150467 294463 160021
rect 306849 151827 306883 161381
rect 270693 139995 270727 144857
rect 294245 140811 294279 150297
rect 310805 147611 310839 153153
rect 337209 152371 337243 154513
rect 284677 126939 284711 132413
rect 235089 113203 235123 122757
rect 239137 118031 239171 122757
rect 251465 115991 251499 125545
rect 270693 120683 270727 125545
rect 272165 120683 272199 125545
rect 288817 121499 288851 122825
rect 230857 95251 230891 104805
rect 232329 87023 232363 100045
rect 251465 96679 251499 106233
rect 265173 96611 265207 104805
rect 266645 96679 266679 106233
rect 267841 106199 267875 114461
rect 290013 113203 290047 122757
rect 291485 121499 291519 139349
rect 296821 132515 296855 142069
rect 301145 132515 301179 142069
rect 302525 124219 302559 133841
rect 306757 124219 306791 133841
rect 310805 128299 310839 138669
rect 325985 132515 326019 143497
rect 330125 138703 330159 143497
rect 339785 142171 339819 151725
rect 341257 143395 341291 160021
rect 358737 154547 358771 162809
rect 372813 159307 372847 164169
rect 367017 144959 367051 154513
rect 375849 143599 375883 153153
rect 358737 135235 358771 143497
rect 360301 137955 360335 143497
rect 372721 135303 372755 138125
rect 327181 129727 327215 135201
rect 295809 111843 295843 121397
rect 296913 113203 296947 122689
rect 301145 114427 301179 122757
rect 306665 113203 306699 122757
rect 310805 116059 310839 125477
rect 337117 124219 337151 133841
rect 310805 108987 310839 115889
rect 325893 104907 325927 117997
rect 330125 113203 330159 122757
rect 337209 118031 337243 122757
rect 358737 114563 358771 124117
rect 367017 116059 367051 125545
rect 372721 115991 372755 125545
rect 375849 124219 375883 133841
rect 389465 122859 389499 133841
rect 236285 87023 236319 96577
rect 247141 89675 247175 96577
rect 267841 95251 267875 104805
rect 272257 96543 272291 104805
rect 273545 95251 273579 104805
rect 327181 103547 327215 113101
rect 367017 106335 367051 115889
rect 374377 104975 374411 114461
rect 375849 104975 375883 114461
rect 377045 106335 377079 115889
rect 285965 93891 285999 103445
rect 295533 92531 295567 101949
rect 232329 75939 232363 85493
rect 236285 75939 236319 85493
rect 247233 77299 247267 80189
rect 251465 77299 251499 86921
rect 284769 85595 284803 90185
rect 301145 86887 301179 93789
rect 291577 84235 291611 85561
rect 306757 84235 306791 93789
rect 317797 89675 317831 96577
rect 330217 86955 330251 98685
rect 337209 93891 337243 103445
rect 244473 66283 244507 70465
rect 250085 66283 250119 75837
rect 265265 73219 265299 82773
rect 270785 74579 270819 84133
rect 230765 48331 230799 61421
rect 232329 56627 232363 66181
rect 266737 64923 266771 74477
rect 272165 66283 272199 75837
rect 284769 75803 284803 84133
rect 273545 67643 273579 70465
rect 285965 66283 285999 78489
rect 301237 73219 301271 82773
rect 302617 73219 302651 82773
rect 323409 75939 323443 77265
rect 324605 75939 324639 85493
rect 232237 38743 232271 53057
rect 236285 48399 236319 61421
rect 250085 51051 250119 56525
rect 262689 55267 262723 60333
rect 265265 53839 265299 63461
rect 270693 52411 270727 66181
rect 230765 37315 230799 38709
rect 236285 37315 236319 46869
rect 247141 34527 247175 46869
rect 250085 37315 250119 46869
rect 251373 37315 251407 46869
rect 270877 42891 270911 52377
rect 265265 35955 265299 41429
rect 236377 19363 236411 28917
rect 251465 26299 251499 35853
rect 266645 34459 266679 41361
rect 273545 38675 273579 48229
rect 285965 46971 285999 56525
rect 294245 55267 294279 64821
rect 295533 48331 295567 57001
rect 296821 56219 296855 66181
rect 301053 55199 301087 69649
rect 337209 66283 337243 84065
rect 339785 77299 339819 95149
rect 341073 77299 341107 103445
rect 357633 95251 357667 104805
rect 358737 95251 358771 104805
rect 374377 99331 374411 104805
rect 367017 87023 367051 96577
rect 375849 95251 375883 104805
rect 377137 99331 377171 106233
rect 389373 87907 389407 99161
rect 341073 70295 341107 77129
rect 357541 75939 357575 85493
rect 360209 77299 360243 86921
rect 372721 66283 372755 75837
rect 389373 67643 389407 77197
rect 310805 60707 310839 66181
rect 300995 55165 301087 55199
rect 302525 46971 302559 59517
rect 323317 48331 323351 66181
rect 324697 56627 324731 66181
rect 329941 56627 329975 66181
rect 339693 46971 339727 56525
rect 341349 50915 341383 57885
rect 367017 48331 367051 57885
rect 389189 48331 389223 57885
rect 470609 48331 470643 57885
rect 358737 46971 358771 48297
rect 284769 29019 284803 44693
rect 296821 43979 296855 46801
rect 288725 27659 288759 37213
rect 230673 11135 230707 12461
rect 244381 8347 244415 24769
rect 265173 18003 265207 27557
rect 285965 18003 285999 27557
rect 288817 16643 288851 26197
rect 273453 10931 273487 16541
rect 295533 12291 295567 27557
rect 299857 18003 299891 37349
rect 303813 32419 303847 42041
rect 323317 37315 323351 46869
rect 324697 37315 324731 46869
rect 327365 38539 327399 46869
rect 330125 37315 330159 46869
rect 338497 27659 338531 45509
rect 341441 38607 341475 41429
rect 377137 38743 377171 41293
rect 367017 29087 367051 38573
rect 372721 29019 372755 31841
rect 301145 18003 301179 27489
rect 310897 16643 310931 26197
rect 327273 9639 327307 17901
rect 330125 9707 330159 27557
rect 337117 19363 337151 24293
rect 358553 9707 358587 27557
rect 367017 19363 367051 28917
rect 375849 19363 375883 28917
rect 377137 22083 377171 28917
rect 366925 12359 366959 19261
rect 389373 8347 389407 17901
rect 227545 6987 227579 7633
rect 268393 5015 268427 5253
rect 220277 4267 220311 4777
rect 249073 4267 249107 4981
rect 278053 5015 278087 5253
rect 287713 5015 287747 5457
rect 297097 5015 297131 5457
rect 258733 4267 258767 4981
rect 307033 4199 307067 4981
rect 319545 4947 319579 5525
rect 320683 4845 320833 4879
rect 320097 4539 320131 4709
rect 320925 4539 320959 4913
rect 324145 4607 324179 5049
rect 325157 4811 325191 4981
rect 326353 4675 326387 4913
rect 327181 4811 327215 5049
rect 326629 4607 326663 4777
rect 326295 4573 326663 4607
rect 45477 3179 45511 3349
rect 82921 2975 82955 3145
rect 93869 2839 93903 2941
rect 263885 1275 263919 4029
rect 278053 3859 278087 4097
rect 282929 3791 282963 4029
rect 287621 3995 287655 4165
rect 287713 3791 287747 3961
rect 318717 3961 319027 3995
rect 273269 3043 273303 3213
rect 282837 3043 282871 3349
rect 287621 3111 287655 3689
rect 318717 3655 318751 3961
rect 318993 3927 319027 3961
rect 318901 3587 318935 3893
rect 331413 3723 331447 3825
rect 332367 3757 332517 3791
rect 338221 3723 338255 3825
rect 322949 2907 322983 3621
rect 326353 3043 326387 3689
rect 349169 3383 349203 4097
rect 322799 2873 322983 2907
rect 335553 2839 335587 3077
rect 336197 2975 336231 3281
rect 345581 3281 345857 3315
rect 345581 2839 345615 3281
rect 350181 3247 350215 4437
rect 350549 4403 350583 4505
rect 351285 4131 351319 4369
rect 339911 2805 340003 2839
rect 354321 3247 354355 4097
rect 345673 2839 345707 3213
rect 354413 2975 354447 3213
rect 359565 2975 359599 3961
rect 360853 3927 360887 4097
rect 360761 2907 360795 3893
rect 361899 3757 361991 3791
rect 361957 3451 361991 3757
rect 362049 3315 362083 3689
rect 363705 3043 363739 3145
rect 369777 2907 369811 3961
rect 376769 3519 376803 4369
rect 445585 3927 445619 4097
rect 445493 3791 445527 3893
rect 376861 3315 376895 3689
rect 413109 3587 413143 3689
rect 420561 3587 420595 3757
rect 376803 3281 376895 3315
rect 422309 2839 422343 3689
rect 425253 3451 425287 3621
rect 431233 3043 431267 3621
rect 431877 2839 431911 3689
rect 433901 3247 433935 3349
rect 441629 3247 441663 3689
rect 446321 3247 446355 4029
rect 446413 3655 446447 3893
rect 446505 3383 446539 3825
rect 446413 2839 446447 3349
rect 446689 3315 446723 3757
rect 451933 2975 451967 3621
rect 451231 2873 451381 2907
rect 451841 2839 451875 2941
rect 339969 2771 340003 2805
rect 454693 2771 454727 4913
rect 461225 4879 461259 5117
rect 466101 4947 466135 5253
rect 471345 4811 471379 5049
rect 471437 4811 471471 5525
rect 456809 2907 456843 3689
rect 460121 3519 460155 3689
rect 460213 3587 460247 3825
rect 466101 3825 466377 3859
rect 460213 3553 460949 3587
rect 461593 3043 461627 3621
rect 461777 3587 461811 3689
rect 463157 3587 463191 3689
rect 466101 3587 466135 3825
rect 463157 3553 463525 3587
rect 466227 3485 466319 3519
rect 466285 2907 466319 3485
rect 466285 2873 466377 2907
rect 471529 595 471563 5593
rect 518173 3043 518207 3213
<< viali >>
rect 364533 685797 364567 685831
rect 364533 676209 364567 676243
rect 429577 684437 429611 684471
rect 559297 684437 559331 684471
rect 429577 666553 429611 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 559297 666553 559331 666587
rect 364533 618205 364567 618239
rect 364533 608617 364567 608651
rect 429393 608549 429427 608583
rect 429393 601681 429427 601715
rect 559113 608549 559147 608583
rect 559113 601681 559147 601715
rect 364625 598893 364659 598927
rect 364625 589305 364659 589339
rect 429577 598893 429611 598927
rect 429577 589305 429611 589339
rect 559297 598893 559331 598927
rect 559297 589305 559331 589339
rect 289737 579581 289771 579615
rect 454049 579581 454083 579615
rect 289921 579513 289955 579547
rect 289737 579445 289771 579479
rect 289829 579445 289863 579479
rect 318809 579445 318843 579479
rect 252109 579309 252143 579343
rect 254225 579309 254259 579343
rect 294613 579309 294647 579343
rect 294613 578969 294647 579003
rect 299305 579309 299339 579343
rect 312001 579309 312035 579343
rect 318809 579309 318843 579343
rect 328377 579445 328411 579479
rect 311817 579241 311851 579275
rect 338129 579445 338163 579479
rect 331321 579309 331355 579343
rect 338129 579309 338163 579343
rect 347697 579445 347731 579479
rect 328377 579241 328411 579275
rect 331137 579241 331171 579275
rect 357449 579445 357483 579479
rect 350641 579309 350675 579343
rect 357449 579309 357483 579343
rect 367017 579445 367051 579479
rect 347697 579241 347731 579275
rect 350457 579241 350491 579275
rect 376769 579445 376803 579479
rect 369961 579309 369995 579343
rect 376769 579309 376803 579343
rect 386337 579445 386371 579479
rect 367017 579241 367051 579275
rect 369777 579241 369811 579275
rect 396089 579445 396123 579479
rect 389281 579309 389315 579343
rect 396089 579309 396123 579343
rect 405657 579445 405691 579479
rect 386337 579241 386371 579275
rect 389097 579241 389131 579275
rect 405657 579241 405691 579275
rect 408509 579445 408543 579479
rect 415317 579445 415351 579479
rect 444297 579445 444331 579479
rect 415317 579309 415351 579343
rect 415685 579377 415719 579411
rect 408509 579241 408543 579275
rect 299305 578969 299339 579003
rect 299121 578833 299155 578867
rect 299397 578833 299431 578867
rect 299213 578765 299247 578799
rect 299305 578765 299339 578799
rect 254225 578629 254259 578663
rect 299121 578629 299155 578663
rect 299305 578629 299339 578663
rect 252109 578561 252143 578595
rect 299029 578561 299063 578595
rect 299213 578561 299247 578595
rect 298937 578493 298971 578527
rect 299121 578493 299155 578527
rect 415685 578493 415719 578527
rect 428381 579377 428415 579411
rect 428381 578425 428415 578459
rect 441077 579309 441111 579343
rect 444297 579241 444331 579275
rect 444389 579445 444423 579479
rect 454049 579445 454083 579479
rect 463617 579581 463651 579615
rect 444389 579241 444423 579275
rect 453589 579377 453623 579411
rect 441077 578357 441111 578391
rect 453589 578289 453623 578323
rect 455797 579377 455831 579411
rect 463617 579309 463651 579343
rect 464445 579309 464479 579343
rect 455797 578221 455831 578255
rect 464445 577881 464479 577915
rect 460581 338113 460615 338147
rect 284401 338045 284435 338079
rect 260481 337569 260515 337603
rect 260481 337365 260515 337399
rect 103437 337229 103471 337263
rect 86969 337093 87003 337127
rect 86969 336957 87003 336991
rect 103437 336957 103471 336991
rect 113189 337229 113223 337263
rect 113189 336753 113223 336787
rect 122757 337229 122791 337263
rect 122757 336753 122791 336787
rect 316693 338045 316727 338079
rect 379437 338045 379471 338079
rect 379529 338045 379563 338079
rect 302249 337773 302283 337807
rect 412557 337977 412591 338011
rect 335921 337841 335955 337875
rect 316693 337297 316727 337331
rect 335829 337501 335863 337535
rect 302249 337161 302283 337195
rect 321845 337229 321879 337263
rect 284401 335189 284435 335223
rect 302525 334713 302559 334747
rect 250177 334441 250211 334475
rect 250177 328457 250211 328491
rect 336013 337841 336047 337875
rect 365729 337841 365763 337875
rect 348985 337705 349019 337739
rect 336013 337637 336047 337671
rect 344661 337637 344695 337671
rect 342821 337501 342855 337535
rect 344293 337501 344327 337535
rect 345673 337569 345707 337603
rect 336105 337433 336139 337467
rect 335829 336753 335863 336787
rect 341717 337161 341751 337195
rect 342821 337093 342855 337127
rect 347789 337433 347823 337467
rect 348985 337433 349019 337467
rect 360117 337705 360151 337739
rect 347789 337297 347823 337331
rect 364349 337705 364383 337739
rect 364993 337637 365027 337671
rect 364441 337501 364475 337535
rect 364717 337501 364751 337535
rect 364349 337365 364383 337399
rect 360117 337297 360151 337331
rect 451197 337977 451231 338011
rect 466377 338113 466411 338147
rect 454693 337909 454727 337943
rect 460581 337909 460615 337943
rect 461593 337977 461627 338011
rect 412465 337773 412499 337807
rect 412557 337773 412591 337807
rect 451105 337773 451139 337807
rect 451197 337773 451231 337807
rect 451289 337773 451323 337807
rect 432245 337705 432279 337739
rect 412465 337637 412499 337671
rect 413937 337637 413971 337671
rect 414305 337637 414339 337671
rect 365729 337569 365763 337603
rect 412649 337569 412683 337603
rect 374653 337433 374687 337467
rect 369869 337365 369903 337399
rect 369869 337161 369903 337195
rect 412649 337297 412683 337331
rect 431877 337501 431911 337535
rect 374653 337161 374687 337195
rect 431877 337161 431911 337195
rect 345857 337093 345891 337127
rect 364993 337093 365027 337127
rect 345581 336753 345615 336787
rect 345765 336957 345799 336991
rect 345857 336957 345891 336991
rect 443469 337637 443503 337671
rect 451105 337637 451139 337671
rect 451289 337501 451323 337535
rect 443469 337365 443503 337399
rect 432245 336957 432279 336991
rect 345765 336753 345799 336787
rect 456993 337569 457027 337603
rect 456993 337297 457027 337331
rect 460397 337569 460431 337603
rect 461593 337569 461627 337603
rect 466285 337977 466319 338011
rect 454693 336753 454727 336787
rect 457177 337229 457211 337263
rect 460397 337229 460431 337263
rect 461593 337297 461627 337331
rect 461593 336821 461627 336855
rect 457177 336753 457211 336787
rect 466377 337773 466411 337807
rect 469229 337909 469263 337943
rect 466469 337297 466503 337331
rect 469229 337229 469263 337263
rect 466469 336889 466503 336923
rect 321845 329137 321879 329171
rect 330217 336685 330251 336719
rect 341717 336685 341751 336719
rect 374469 336685 374503 336719
rect 302525 328457 302559 328491
rect 259837 328389 259871 328423
rect 330217 327165 330251 327199
rect 331413 336073 331447 336107
rect 341717 335529 341751 335563
rect 341717 328457 341751 328491
rect 331413 327097 331447 327131
rect 374469 327097 374503 327131
rect 375849 336685 375883 336719
rect 466285 336685 466319 336719
rect 375849 327097 375883 327131
rect 389557 328389 389591 328423
rect 357449 327029 357483 327063
rect 337209 321589 337243 321623
rect 337209 320841 337243 320875
rect 341441 321589 341475 321623
rect 259837 318801 259871 318835
rect 341441 318801 341475 318835
rect 230857 318733 230891 318767
rect 236285 318733 236319 318767
rect 236285 309213 236319 309247
rect 239229 318733 239263 318767
rect 230857 309145 230891 309179
rect 284677 318733 284711 318767
rect 262597 315945 262631 315979
rect 239229 309145 239263 309179
rect 244473 311797 244507 311831
rect 244473 309145 244507 309179
rect 236285 309077 236319 309111
rect 236285 299557 236319 299591
rect 259653 309077 259687 309111
rect 259653 299557 259687 299591
rect 236285 299421 236319 299455
rect 357449 317441 357483 317475
rect 360393 327029 360427 327063
rect 389557 318801 389591 318835
rect 470609 328389 470643 328423
rect 470609 318801 470643 318835
rect 360393 317441 360427 317475
rect 284677 314177 284711 314211
rect 299765 317373 299799 317407
rect 273453 313429 273487 313463
rect 273453 311865 273487 311899
rect 325893 317373 325927 317407
rect 310897 311933 310931 311967
rect 310897 307853 310931 307887
rect 337209 317373 337243 317407
rect 337209 311729 337243 311763
rect 375849 317373 375883 317407
rect 325893 307785 325927 307819
rect 341165 309077 341199 309111
rect 299765 299489 299799 299523
rect 310713 307717 310747 307751
rect 262597 298197 262631 298231
rect 327181 307717 327215 307751
rect 310713 298129 310747 298163
rect 323317 299421 323351 299455
rect 266737 298061 266771 298095
rect 251465 294661 251499 294695
rect 236285 289833 236319 289867
rect 239229 292553 239263 292587
rect 239229 289833 239263 289867
rect 251465 289833 251499 289867
rect 244473 289765 244507 289799
rect 236285 289697 236319 289731
rect 236285 280245 236319 280279
rect 266737 288405 266771 288439
rect 267749 298061 267783 298095
rect 285965 298061 285999 298095
rect 267749 288405 267783 288439
rect 270785 292485 270819 292519
rect 310897 293029 310931 293063
rect 285965 288405 285999 288439
rect 294245 289833 294279 289867
rect 294245 287045 294279 287079
rect 270785 285617 270819 285651
rect 324697 299421 324731 299455
rect 327181 298129 327215 298163
rect 337209 307717 337243 307751
rect 341165 299489 341199 299523
rect 357817 309077 357851 309111
rect 357817 299489 357851 299523
rect 358737 309077 358771 309111
rect 470609 309077 470643 309111
rect 375849 307785 375883 307819
rect 389281 309009 389315 309043
rect 358737 299489 358771 299523
rect 374377 307717 374411 307751
rect 337209 298129 337243 298163
rect 372721 299421 372755 299455
rect 324697 289833 324731 289867
rect 358737 298061 358771 298095
rect 323317 288405 323351 288439
rect 327181 289765 327215 289799
rect 357449 289765 357483 289799
rect 310897 282761 310931 282795
rect 323501 283577 323535 283611
rect 327181 283577 327215 283611
rect 337209 285617 337243 285651
rect 244473 280177 244507 280211
rect 236285 280109 236319 280143
rect 236285 270521 236319 270555
rect 239137 280109 239171 280143
rect 239137 270521 239171 270555
rect 251465 280109 251499 280143
rect 259561 280109 259595 280143
rect 323501 278749 323535 278783
rect 331413 280109 331447 280143
rect 259561 273037 259595 273071
rect 310897 278681 310931 278715
rect 251465 270521 251499 270555
rect 236285 270385 236319 270419
rect 236285 260933 236319 260967
rect 250085 269025 250119 269059
rect 236285 260797 236319 260831
rect 236285 251209 236319 251243
rect 239137 260797 239171 260831
rect 330125 273853 330159 273887
rect 341165 282897 341199 282931
rect 341165 280177 341199 280211
rect 372721 289833 372755 289867
rect 389281 299489 389315 299523
rect 470609 299489 470643 299523
rect 374377 289833 374411 289867
rect 375849 299421 375883 299455
rect 375849 289833 375883 289867
rect 358737 288405 358771 288439
rect 389373 289765 389407 289799
rect 357449 280177 357483 280211
rect 389373 280177 389407 280211
rect 470609 289765 470643 289799
rect 470609 280177 470643 280211
rect 337209 276029 337243 276063
rect 338865 280109 338899 280143
rect 331413 270521 331447 270555
rect 338865 270521 338899 270555
rect 372721 280109 372755 280143
rect 372721 270521 372755 270555
rect 377137 280109 377171 280143
rect 377137 270521 377171 270555
rect 330125 269093 330159 269127
rect 389373 270453 389407 270487
rect 310897 263449 310931 263483
rect 262597 260865 262631 260899
rect 389373 260865 389407 260899
rect 470609 270453 470643 270487
rect 470609 260865 470643 260899
rect 250085 259437 250119 259471
rect 251465 260797 251499 260831
rect 239137 251209 239171 251243
rect 250177 259301 250211 259335
rect 259561 260797 259595 260831
rect 262597 259437 262631 259471
rect 270693 260797 270727 260831
rect 259561 253725 259595 253759
rect 251465 251209 251499 251243
rect 250177 251073 250211 251107
rect 259561 251141 259595 251175
rect 338865 260797 338899 260831
rect 270693 251073 270727 251107
rect 306757 258009 306791 258043
rect 310897 256037 310931 256071
rect 310897 251277 310931 251311
rect 337117 253997 337151 254031
rect 306757 248353 306791 248387
rect 310713 251141 310747 251175
rect 285965 244953 285999 244987
rect 259561 244137 259595 244171
rect 272165 244409 272199 244443
rect 272165 241553 272199 241587
rect 267749 240057 267783 240091
rect 266737 234821 266771 234855
rect 272165 240057 272199 240091
rect 272165 234481 272199 234515
rect 341073 260797 341107 260831
rect 372721 260797 372755 260831
rect 341073 253725 341107 253759
rect 357541 259369 357575 259403
rect 338865 251209 338899 251243
rect 372721 251209 372755 251243
rect 377137 260797 377171 260831
rect 377137 251209 377171 251243
rect 463709 260797 463743 260831
rect 463709 251209 463743 251243
rect 357541 249781 357575 249815
rect 470609 251141 470643 251175
rect 337117 247129 337151 247163
rect 337117 246993 337151 247027
rect 337117 244205 337151 244239
rect 310713 241485 310747 241519
rect 470609 241485 470643 241519
rect 299489 241417 299523 241451
rect 285965 234481 285999 234515
rect 290381 238697 290415 238731
rect 267749 231761 267783 231795
rect 266737 230469 266771 230503
rect 290381 230401 290415 230435
rect 295625 238697 295659 238731
rect 331413 241417 331447 241451
rect 299489 231829 299523 231863
rect 306941 238765 306975 238799
rect 389281 241417 389315 241451
rect 389281 234617 389315 234651
rect 331413 231829 331447 231863
rect 306941 230469 306975 230503
rect 310805 231761 310839 231795
rect 295625 229109 295659 229143
rect 270693 224961 270727 224995
rect 310805 222173 310839 222207
rect 337117 231625 337151 231659
rect 270693 220813 270727 220847
rect 299489 222105 299523 222139
rect 290197 219385 290231 219419
rect 290197 212449 290231 212483
rect 291669 219385 291703 219419
rect 341073 224961 341107 224995
rect 341073 222173 341107 222207
rect 337117 220813 337151 220847
rect 299489 212517 299523 212551
rect 291669 212449 291703 212483
rect 310805 212449 310839 212483
rect 302617 207757 302651 207791
rect 270693 205649 270727 205683
rect 270693 202861 270727 202895
rect 302617 202861 302651 202895
rect 310805 202861 310839 202895
rect 250085 200073 250119 200107
rect 367017 193137 367051 193171
rect 299857 190417 299891 190451
rect 288725 188989 288759 189023
rect 250085 186269 250119 186303
rect 267749 186337 267783 186371
rect 267749 183549 267783 183583
rect 270693 186337 270727 186371
rect 270693 183549 270727 183583
rect 232329 182121 232363 182155
rect 284769 180761 284803 180795
rect 259653 179537 259687 179571
rect 259653 173961 259687 173995
rect 265265 179333 265299 179367
rect 232329 172533 232363 172567
rect 232237 172465 232271 172499
rect 232237 164169 232271 164203
rect 299857 180829 299891 180863
rect 302525 190417 302559 190451
rect 302525 180829 302559 180863
rect 306849 190417 306883 190451
rect 339785 188377 339819 188411
rect 339785 183549 339819 183583
rect 367017 183549 367051 183583
rect 306849 180829 306883 180863
rect 358737 181985 358771 182019
rect 288725 179401 288759 179435
rect 341257 179333 341291 179367
rect 284769 171105 284803 171139
rect 337117 172465 337151 172499
rect 267841 171037 267875 171071
rect 267841 162741 267875 162775
rect 294429 171037 294463 171071
rect 265265 161449 265299 161483
rect 366925 174029 366959 174063
rect 366925 173893 366959 173927
rect 358737 173825 358771 173859
rect 341257 169745 341291 169779
rect 337117 164169 337151 164203
rect 372813 164169 372847 164203
rect 294429 161449 294463 161483
rect 358737 162809 358771 162843
rect 267841 161381 267875 161415
rect 259653 154173 259687 154207
rect 306849 161381 306883 161415
rect 267841 151793 267875 151827
rect 291485 160021 291519 160055
rect 259653 144993 259687 145027
rect 264989 151725 265023 151759
rect 250269 143497 250303 143531
rect 294429 160021 294463 160055
rect 341257 160021 341291 160055
rect 337209 154513 337243 154547
rect 306849 151793 306883 151827
rect 310805 153153 310839 153187
rect 294429 150433 294463 150467
rect 291485 149073 291519 149107
rect 294245 150297 294279 150331
rect 264989 142137 265023 142171
rect 270693 144857 270727 144891
rect 337209 152337 337243 152371
rect 310805 147577 310839 147611
rect 339785 151725 339819 151759
rect 325985 143497 326019 143531
rect 294245 140777 294279 140811
rect 296821 142069 296855 142103
rect 270693 139961 270727 139995
rect 250269 133909 250303 133943
rect 291485 139349 291519 139383
rect 284677 132413 284711 132447
rect 284677 126905 284711 126939
rect 251465 125545 251499 125579
rect 235089 122757 235123 122791
rect 239137 122757 239171 122791
rect 239137 117997 239171 118031
rect 270693 125545 270727 125579
rect 270693 120649 270727 120683
rect 272165 125545 272199 125579
rect 288817 122825 288851 122859
rect 288817 121465 288851 121499
rect 290013 122757 290047 122791
rect 272165 120649 272199 120683
rect 251465 115957 251499 115991
rect 235089 113169 235123 113203
rect 267841 114461 267875 114495
rect 251465 106233 251499 106267
rect 230857 104805 230891 104839
rect 230857 95217 230891 95251
rect 232329 100045 232363 100079
rect 266645 106233 266679 106267
rect 251465 96645 251499 96679
rect 265173 104805 265207 104839
rect 296821 132481 296855 132515
rect 301145 142069 301179 142103
rect 310805 138669 310839 138703
rect 301145 132481 301179 132515
rect 302525 133841 302559 133875
rect 302525 124185 302559 124219
rect 306757 133841 306791 133875
rect 330125 143497 330159 143531
rect 372813 159273 372847 159307
rect 358737 154513 358771 154547
rect 367017 154513 367051 154547
rect 367017 144925 367051 144959
rect 375849 153153 375883 153187
rect 375849 143565 375883 143599
rect 341257 143361 341291 143395
rect 358737 143497 358771 143531
rect 339785 142137 339819 142171
rect 330125 138669 330159 138703
rect 360301 143497 360335 143531
rect 360301 137921 360335 137955
rect 372721 138125 372755 138159
rect 372721 135269 372755 135303
rect 325985 132481 326019 132515
rect 327181 135201 327215 135235
rect 358737 135201 358771 135235
rect 327181 129693 327215 129727
rect 337117 133841 337151 133875
rect 310805 128265 310839 128299
rect 306757 124185 306791 124219
rect 310805 125477 310839 125511
rect 301145 122757 301179 122791
rect 291485 121465 291519 121499
rect 296913 122689 296947 122723
rect 290013 113169 290047 113203
rect 295809 121397 295843 121431
rect 301145 114393 301179 114427
rect 306665 122757 306699 122791
rect 296913 113169 296947 113203
rect 375849 133841 375883 133875
rect 337117 124185 337151 124219
rect 367017 125545 367051 125579
rect 358737 124117 358771 124151
rect 330125 122757 330159 122791
rect 310805 116025 310839 116059
rect 325893 117997 325927 118031
rect 306665 113169 306699 113203
rect 310805 115889 310839 115923
rect 295809 111809 295843 111843
rect 310805 108953 310839 108987
rect 267841 106165 267875 106199
rect 337209 122757 337243 122791
rect 337209 117997 337243 118031
rect 367017 116025 367051 116059
rect 372721 125545 372755 125579
rect 375849 124185 375883 124219
rect 389465 133841 389499 133875
rect 389465 122825 389499 122859
rect 372721 115957 372755 115991
rect 358737 114529 358771 114563
rect 367017 115889 367051 115923
rect 330125 113169 330159 113203
rect 325893 104873 325927 104907
rect 327181 113101 327215 113135
rect 266645 96645 266679 96679
rect 267841 104805 267875 104839
rect 232329 86989 232363 87023
rect 236285 96577 236319 96611
rect 247141 96577 247175 96611
rect 265173 96577 265207 96611
rect 272257 104805 272291 104839
rect 272257 96509 272291 96543
rect 273545 104805 273579 104839
rect 267841 95217 267875 95251
rect 377045 115889 377079 115923
rect 367017 106301 367051 106335
rect 374377 114461 374411 114495
rect 374377 104941 374411 104975
rect 375849 114461 375883 114495
rect 377045 106301 377079 106335
rect 375849 104941 375883 104975
rect 377137 106233 377171 106267
rect 327181 103513 327215 103547
rect 357633 104805 357667 104839
rect 273545 95217 273579 95251
rect 285965 103445 285999 103479
rect 337209 103445 337243 103479
rect 285965 93857 285999 93891
rect 295533 101949 295567 101983
rect 330217 98685 330251 98719
rect 317797 96577 317831 96611
rect 295533 92497 295567 92531
rect 301145 93789 301179 93823
rect 247141 89641 247175 89675
rect 284769 90185 284803 90219
rect 236285 86989 236319 87023
rect 251465 86921 251499 86955
rect 232329 85493 232363 85527
rect 232329 75905 232363 75939
rect 236285 85493 236319 85527
rect 247233 80189 247267 80223
rect 247233 77265 247267 77299
rect 301145 86853 301179 86887
rect 306757 93789 306791 93823
rect 284769 85561 284803 85595
rect 291577 85561 291611 85595
rect 291577 84201 291611 84235
rect 317797 89641 317831 89675
rect 341073 103445 341107 103479
rect 337209 93857 337243 93891
rect 339785 95149 339819 95183
rect 330217 86921 330251 86955
rect 306757 84201 306791 84235
rect 324605 85493 324639 85527
rect 270785 84133 270819 84167
rect 251465 77265 251499 77299
rect 265265 82773 265299 82807
rect 236285 75905 236319 75939
rect 250085 75837 250119 75871
rect 244473 70465 244507 70499
rect 244473 66249 244507 66283
rect 284769 84133 284803 84167
rect 270785 74545 270819 74579
rect 272165 75837 272199 75871
rect 265265 73185 265299 73219
rect 266737 74477 266771 74511
rect 250085 66249 250119 66283
rect 232329 66181 232363 66215
rect 230765 61421 230799 61455
rect 301237 82773 301271 82807
rect 284769 75769 284803 75803
rect 285965 78489 285999 78523
rect 273545 70465 273579 70499
rect 273545 67609 273579 67643
rect 272165 66249 272199 66283
rect 301237 73185 301271 73219
rect 302617 82773 302651 82807
rect 323409 77265 323443 77299
rect 323409 75905 323443 75939
rect 324605 75905 324639 75939
rect 337209 84065 337243 84099
rect 302617 73185 302651 73219
rect 285965 66249 285999 66283
rect 301053 69649 301087 69683
rect 266737 64889 266771 64923
rect 270693 66181 270727 66215
rect 265265 63461 265299 63495
rect 232329 56593 232363 56627
rect 236285 61421 236319 61455
rect 230765 48297 230799 48331
rect 232237 53057 232271 53091
rect 262689 60333 262723 60367
rect 250085 56525 250119 56559
rect 262689 55233 262723 55267
rect 265265 53805 265299 53839
rect 296821 66181 296855 66215
rect 294245 64821 294279 64855
rect 285965 56525 285999 56559
rect 270693 52377 270727 52411
rect 270877 52377 270911 52411
rect 250085 51017 250119 51051
rect 236285 48365 236319 48399
rect 230765 38709 230799 38743
rect 232237 38709 232271 38743
rect 236285 46869 236319 46903
rect 230765 37281 230799 37315
rect 236285 37281 236319 37315
rect 247141 46869 247175 46903
rect 250085 46869 250119 46903
rect 250085 37281 250119 37315
rect 251373 46869 251407 46903
rect 270877 42857 270911 42891
rect 273545 48229 273579 48263
rect 251373 37281 251407 37315
rect 265265 41429 265299 41463
rect 265265 35921 265299 35955
rect 266645 41361 266679 41395
rect 247141 34493 247175 34527
rect 251465 35853 251499 35887
rect 236377 28917 236411 28951
rect 294245 55233 294279 55267
rect 295533 57001 295567 57035
rect 296821 56185 296855 56219
rect 339785 77265 339819 77299
rect 357633 95217 357667 95251
rect 358737 104805 358771 104839
rect 374377 104805 374411 104839
rect 374377 99297 374411 99331
rect 375849 104805 375883 104839
rect 358737 95217 358771 95251
rect 367017 96577 367051 96611
rect 377137 99297 377171 99331
rect 375849 95217 375883 95251
rect 389373 99161 389407 99195
rect 389373 87873 389407 87907
rect 367017 86989 367051 87023
rect 360209 86921 360243 86955
rect 341073 77265 341107 77299
rect 357541 85493 357575 85527
rect 341073 77129 341107 77163
rect 360209 77265 360243 77299
rect 357541 75905 357575 75939
rect 389373 77197 389407 77231
rect 341073 70261 341107 70295
rect 372721 75837 372755 75871
rect 337209 66249 337243 66283
rect 389373 67609 389407 67643
rect 372721 66249 372755 66283
rect 310805 66181 310839 66215
rect 310805 60673 310839 60707
rect 323317 66181 323351 66215
rect 300961 55165 300995 55199
rect 302525 59517 302559 59551
rect 295533 48297 295567 48331
rect 285965 46937 285999 46971
rect 324697 66181 324731 66215
rect 324697 56593 324731 56627
rect 329941 66181 329975 66215
rect 329941 56593 329975 56627
rect 341349 57885 341383 57919
rect 323317 48297 323351 48331
rect 339693 56525 339727 56559
rect 302525 46937 302559 46971
rect 341349 50881 341383 50915
rect 367017 57885 367051 57919
rect 339693 46937 339727 46971
rect 358737 48297 358771 48331
rect 367017 48297 367051 48331
rect 389189 57885 389223 57919
rect 389189 48297 389223 48331
rect 470609 57885 470643 57919
rect 470609 48297 470643 48331
rect 358737 46937 358771 46971
rect 323317 46869 323351 46903
rect 296821 46801 296855 46835
rect 273545 38641 273579 38675
rect 284769 44693 284803 44727
rect 266645 34425 266679 34459
rect 296821 43945 296855 43979
rect 303813 42041 303847 42075
rect 299857 37349 299891 37383
rect 284769 28985 284803 29019
rect 288725 37213 288759 37247
rect 288725 27625 288759 27659
rect 251465 26265 251499 26299
rect 265173 27557 265207 27591
rect 236377 19329 236411 19363
rect 244381 24769 244415 24803
rect 230673 12461 230707 12495
rect 230673 11101 230707 11135
rect 265173 17969 265207 18003
rect 285965 27557 285999 27591
rect 295533 27557 295567 27591
rect 285965 17969 285999 18003
rect 288817 26197 288851 26231
rect 288817 16609 288851 16643
rect 273453 16541 273487 16575
rect 323317 37281 323351 37315
rect 324697 46869 324731 46903
rect 327365 46869 327399 46903
rect 327365 38505 327399 38539
rect 330125 46869 330159 46903
rect 324697 37281 324731 37315
rect 330125 37281 330159 37315
rect 338497 45509 338531 45543
rect 303813 32385 303847 32419
rect 341441 41429 341475 41463
rect 377137 41293 377171 41327
rect 377137 38709 377171 38743
rect 341441 38573 341475 38607
rect 367017 38573 367051 38607
rect 367017 29053 367051 29087
rect 372721 31841 372755 31875
rect 372721 28985 372755 29019
rect 338497 27625 338531 27659
rect 367017 28917 367051 28951
rect 330125 27557 330159 27591
rect 299857 17969 299891 18003
rect 301145 27489 301179 27523
rect 301145 17969 301179 18003
rect 310897 26197 310931 26231
rect 310897 16609 310931 16643
rect 327273 17901 327307 17935
rect 295533 12257 295567 12291
rect 273453 10897 273487 10931
rect 358553 27557 358587 27591
rect 337117 24293 337151 24327
rect 337117 19329 337151 19363
rect 330125 9673 330159 9707
rect 367017 19329 367051 19363
rect 375849 28917 375883 28951
rect 377137 28917 377171 28951
rect 377137 22049 377171 22083
rect 375849 19329 375883 19363
rect 366925 19261 366959 19295
rect 366925 12325 366959 12359
rect 389373 17901 389407 17935
rect 358553 9673 358587 9707
rect 327273 9605 327307 9639
rect 244381 8313 244415 8347
rect 389373 8313 389407 8347
rect 227545 7633 227579 7667
rect 227545 6953 227579 6987
rect 471529 5593 471563 5627
rect 319545 5525 319579 5559
rect 287713 5457 287747 5491
rect 268393 5253 268427 5287
rect 249073 4981 249107 5015
rect 220277 4777 220311 4811
rect 220277 4233 220311 4267
rect 249073 4233 249107 4267
rect 258733 4981 258767 5015
rect 268393 4981 268427 5015
rect 278053 5253 278087 5287
rect 278053 4981 278087 5015
rect 287713 4981 287747 5015
rect 297097 5457 297131 5491
rect 297097 4981 297131 5015
rect 307033 4981 307067 5015
rect 258733 4233 258767 4267
rect 471437 5525 471471 5559
rect 466101 5253 466135 5287
rect 461225 5117 461259 5151
rect 324145 5049 324179 5083
rect 319545 4913 319579 4947
rect 320925 4913 320959 4947
rect 320649 4845 320683 4879
rect 320833 4845 320867 4879
rect 320097 4709 320131 4743
rect 320097 4505 320131 4539
rect 327181 5049 327215 5083
rect 325157 4981 325191 5015
rect 325157 4777 325191 4811
rect 326353 4913 326387 4947
rect 326353 4641 326387 4675
rect 326629 4777 326663 4811
rect 327181 4777 327215 4811
rect 454693 4913 454727 4947
rect 324145 4573 324179 4607
rect 326261 4573 326295 4607
rect 320925 4505 320959 4539
rect 350549 4505 350583 4539
rect 287621 4165 287655 4199
rect 307033 4165 307067 4199
rect 350181 4437 350215 4471
rect 278053 4097 278087 4131
rect 263885 4029 263919 4063
rect 45477 3349 45511 3383
rect 45477 3145 45511 3179
rect 82921 3145 82955 3179
rect 82921 2941 82955 2975
rect 93869 2941 93903 2975
rect 93869 2805 93903 2839
rect 278053 3825 278087 3859
rect 282929 4029 282963 4063
rect 349169 4097 349203 4131
rect 287621 3961 287655 3995
rect 287713 3961 287747 3995
rect 282929 3757 282963 3791
rect 287713 3757 287747 3791
rect 287621 3689 287655 3723
rect 282837 3349 282871 3383
rect 273269 3213 273303 3247
rect 273269 3009 273303 3043
rect 318717 3621 318751 3655
rect 318901 3893 318935 3927
rect 318993 3893 319027 3927
rect 331413 3825 331447 3859
rect 338221 3825 338255 3859
rect 332333 3757 332367 3791
rect 332517 3757 332551 3791
rect 326353 3689 326387 3723
rect 331413 3689 331447 3723
rect 338221 3689 338255 3723
rect 318901 3553 318935 3587
rect 322949 3621 322983 3655
rect 287621 3077 287655 3111
rect 282837 3009 282871 3043
rect 349169 3349 349203 3383
rect 336197 3281 336231 3315
rect 326353 3009 326387 3043
rect 335553 3077 335587 3111
rect 322765 2873 322799 2907
rect 336197 2941 336231 2975
rect 345857 3281 345891 3315
rect 350549 4369 350583 4403
rect 351285 4369 351319 4403
rect 376769 4369 376803 4403
rect 351285 4097 351319 4131
rect 354321 4097 354355 4131
rect 335553 2805 335587 2839
rect 339877 2805 339911 2839
rect 345581 2805 345615 2839
rect 345673 3213 345707 3247
rect 350181 3213 350215 3247
rect 360853 4097 360887 4131
rect 359565 3961 359599 3995
rect 354321 3213 354355 3247
rect 354413 3213 354447 3247
rect 354413 2941 354447 2975
rect 359565 2941 359599 2975
rect 360761 3893 360795 3927
rect 360853 3893 360887 3927
rect 369777 3961 369811 3995
rect 361865 3757 361899 3791
rect 361957 3417 361991 3451
rect 362049 3689 362083 3723
rect 362049 3281 362083 3315
rect 363705 3145 363739 3179
rect 363705 3009 363739 3043
rect 360761 2873 360795 2907
rect 445585 4097 445619 4131
rect 445493 3893 445527 3927
rect 445585 3893 445619 3927
rect 446321 4029 446355 4063
rect 420561 3757 420595 3791
rect 445493 3757 445527 3791
rect 376769 3485 376803 3519
rect 376861 3689 376895 3723
rect 413109 3689 413143 3723
rect 413109 3553 413143 3587
rect 420561 3553 420595 3587
rect 422309 3689 422343 3723
rect 376769 3281 376803 3315
rect 369777 2873 369811 2907
rect 345673 2805 345707 2839
rect 431877 3689 431911 3723
rect 425253 3621 425287 3655
rect 425253 3417 425287 3451
rect 431233 3621 431267 3655
rect 431233 3009 431267 3043
rect 422309 2805 422343 2839
rect 441629 3689 441663 3723
rect 433901 3349 433935 3383
rect 433901 3213 433935 3247
rect 441629 3213 441663 3247
rect 446413 3893 446447 3927
rect 446413 3621 446447 3655
rect 446505 3825 446539 3859
rect 446321 3213 446355 3247
rect 446413 3349 446447 3383
rect 446505 3349 446539 3383
rect 446689 3757 446723 3791
rect 431877 2805 431911 2839
rect 446689 3281 446723 3315
rect 451933 3621 451967 3655
rect 451841 2941 451875 2975
rect 451933 2941 451967 2975
rect 451197 2873 451231 2907
rect 451381 2873 451415 2907
rect 446413 2805 446447 2839
rect 451841 2805 451875 2839
rect 339969 2737 340003 2771
rect 466101 4913 466135 4947
rect 471345 5049 471379 5083
rect 461225 4845 461259 4879
rect 471345 4777 471379 4811
rect 471437 4777 471471 4811
rect 460213 3825 460247 3859
rect 456809 3689 456843 3723
rect 460121 3689 460155 3723
rect 466377 3825 466411 3859
rect 461777 3689 461811 3723
rect 461593 3621 461627 3655
rect 460949 3553 460983 3587
rect 460121 3485 460155 3519
rect 461777 3553 461811 3587
rect 463157 3689 463191 3723
rect 463525 3553 463559 3587
rect 466101 3553 466135 3587
rect 466193 3485 466227 3519
rect 461593 3009 461627 3043
rect 456809 2873 456843 2907
rect 466377 2873 466411 2907
rect 454693 2737 454727 2771
rect 263885 1241 263919 1275
rect 518173 3213 518207 3247
rect 518173 3009 518207 3043
rect 471529 561 471563 595
<< metal1 >>
rect 202782 700952 202788 701004
rect 202840 700992 202846 701004
rect 358814 700992 358820 701004
rect 202840 700964 358820 700992
rect 202840 700952 202846 700964
rect 358814 700952 358820 700964
rect 358872 700952 358878 701004
rect 170306 700884 170312 700936
rect 170364 700924 170370 700936
rect 362954 700924 362960 700936
rect 170364 700896 362960 700924
rect 170364 700884 170370 700896
rect 362954 700884 362960 700896
rect 363012 700884 363018 700936
rect 328362 700816 328368 700868
rect 328420 700856 328426 700868
rect 527174 700856 527180 700868
rect 328420 700828 527180 700856
rect 328420 700816 328426 700828
rect 527174 700816 527180 700828
rect 527232 700816 527238 700868
rect 329742 700748 329748 700800
rect 329800 700788 329806 700800
rect 543458 700788 543464 700800
rect 329800 700760 543464 700788
rect 329800 700748 329806 700760
rect 543458 700748 543464 700760
rect 543516 700748 543522 700800
rect 154114 700680 154120 700732
rect 154172 700720 154178 700732
rect 367094 700720 367100 700732
rect 154172 700692 367100 700720
rect 154172 700680 154178 700692
rect 367094 700680 367100 700692
rect 367152 700680 367158 700732
rect 137830 700612 137836 700664
rect 137888 700652 137894 700664
rect 364334 700652 364340 700664
rect 137888 700624 364340 700652
rect 137888 700612 137894 700624
rect 364334 700612 364340 700624
rect 364392 700612 364398 700664
rect 105446 700544 105452 700596
rect 105504 700584 105510 700596
rect 368474 700584 368480 700596
rect 105504 700556 368480 700584
rect 105504 700544 105510 700556
rect 368474 700544 368480 700556
rect 368532 700544 368538 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 373994 700516 374000 700528
rect 89220 700488 374000 700516
rect 89220 700476 89226 700488
rect 373994 700476 374000 700488
rect 374052 700476 374058 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 371234 700448 371240 700460
rect 73028 700420 371240 700448
rect 73028 700408 73034 700420
rect 371234 700408 371240 700420
rect 371292 700408 371298 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 375374 700380 375380 700392
rect 40552 700352 375380 700380
rect 40552 700340 40558 700352
rect 375374 700340 375380 700352
rect 375432 700340 375438 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 379514 700312 379520 700324
rect 24360 700284 379520 700312
rect 24360 700272 24366 700284
rect 379514 700272 379520 700284
rect 379572 700272 379578 700324
rect 218974 700204 218980 700256
rect 219032 700244 219038 700256
rect 360194 700244 360200 700256
rect 219032 700216 360200 700244
rect 219032 700204 219038 700216
rect 360194 700204 360200 700216
rect 360252 700204 360258 700256
rect 336642 700136 336648 700188
rect 336700 700176 336706 700188
rect 478506 700176 478512 700188
rect 336700 700148 478512 700176
rect 336700 700136 336706 700148
rect 478506 700136 478512 700148
rect 478564 700136 478570 700188
rect 335262 700068 335268 700120
rect 335320 700108 335326 700120
rect 462314 700108 462320 700120
rect 335320 700080 462320 700108
rect 335320 700068 335326 700080
rect 462314 700068 462320 700080
rect 462372 700068 462378 700120
rect 235166 700000 235172 700052
rect 235224 700040 235230 700052
rect 356054 700040 356060 700052
rect 235224 700012 356060 700040
rect 235224 700000 235230 700012
rect 356054 700000 356060 700012
rect 356112 700000 356118 700052
rect 267642 699932 267648 699984
rect 267700 699972 267706 699984
rect 351914 699972 351920 699984
rect 267700 699944 351920 699972
rect 267700 699932 267706 699944
rect 351914 699932 351920 699944
rect 351972 699932 351978 699984
rect 283834 699864 283840 699916
rect 283892 699904 283898 699916
rect 354674 699904 354680 699916
rect 283892 699876 354680 699904
rect 283892 699864 283898 699876
rect 354674 699864 354680 699876
rect 354732 699864 354738 699916
rect 343542 699796 343548 699848
rect 343600 699836 343606 699848
rect 413646 699836 413652 699848
rect 343600 699808 413652 699836
rect 343600 699796 343606 699808
rect 413646 699796 413652 699808
rect 413704 699796 413710 699848
rect 340782 699728 340788 699780
rect 340840 699768 340846 699780
rect 397454 699768 397460 699780
rect 340840 699740 397460 699768
rect 340840 699728 340846 699740
rect 397454 699728 397460 699740
rect 397512 699728 397518 699780
rect 300118 699660 300124 699712
rect 300176 699700 300182 699712
rect 300762 699700 300768 699712
rect 300176 699672 300768 699700
rect 300176 699660 300182 699672
rect 300762 699660 300768 699672
rect 300820 699660 300826 699712
rect 332502 699660 332508 699712
rect 332560 699700 332566 699712
rect 346394 699700 346400 699712
rect 332560 699672 346400 699700
rect 332560 699660 332566 699672
rect 346394 699660 346400 699672
rect 346452 699660 346458 699712
rect 347774 699660 347780 699712
rect 347832 699700 347838 699712
rect 348786 699700 348792 699712
rect 347832 699672 348792 699700
rect 347832 699660 347838 699672
rect 348786 699660 348792 699672
rect 348844 699660 348850 699712
rect 321462 696940 321468 696992
rect 321520 696980 321526 696992
rect 580166 696980 580172 696992
rect 321520 696952 580172 696980
rect 321520 696940 321526 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 429378 688576 429384 688628
rect 429436 688616 429442 688628
rect 429838 688616 429844 688628
rect 429436 688588 429844 688616
rect 429436 688576 429442 688588
rect 429838 688576 429844 688588
rect 429896 688576 429902 688628
rect 559098 688576 559104 688628
rect 559156 688616 559162 688628
rect 559650 688616 559656 688628
rect 559156 688588 559656 688616
rect 559156 688576 559162 688588
rect 559650 688576 559656 688588
rect 559708 688576 559714 688628
rect 364610 687760 364616 687812
rect 364668 687800 364674 687812
rect 365162 687800 365168 687812
rect 364668 687772 365168 687800
rect 364668 687760 364674 687772
rect 365162 687760 365168 687772
rect 365220 687760 365226 687812
rect 429212 685936 429976 685964
rect 324222 685856 324228 685908
rect 324280 685896 324286 685908
rect 429212 685896 429240 685936
rect 324280 685868 429240 685896
rect 429948 685896 429976 685936
rect 552584 685936 559788 685964
rect 552584 685896 552612 685936
rect 429948 685868 552612 685896
rect 559760 685896 559788 685936
rect 580166 685896 580172 685908
rect 559760 685868 580172 685896
rect 324280 685856 324286 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 364521 685831 364579 685837
rect 364521 685797 364533 685831
rect 364567 685828 364579 685831
rect 364610 685828 364616 685840
rect 364567 685800 364616 685828
rect 364567 685797 364579 685800
rect 364521 685791 364579 685797
rect 364610 685788 364616 685800
rect 364668 685788 364674 685840
rect 429286 684428 429292 684480
rect 429344 684468 429350 684480
rect 429565 684471 429623 684477
rect 429565 684468 429577 684471
rect 429344 684440 429577 684468
rect 429344 684428 429350 684440
rect 429565 684437 429577 684440
rect 429611 684437 429623 684471
rect 429565 684431 429623 684437
rect 559006 684428 559012 684480
rect 559064 684468 559070 684480
rect 559285 684471 559343 684477
rect 559285 684468 559297 684471
rect 559064 684440 559297 684468
rect 559064 684428 559070 684440
rect 559285 684437 559297 684440
rect 559331 684437 559343 684471
rect 559285 684431 559343 684437
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 382274 681748 382280 681760
rect 3568 681720 382280 681748
rect 3568 681708 3574 681720
rect 382274 681708 382280 681720
rect 382332 681708 382338 681760
rect 364518 676240 364524 676252
rect 364479 676212 364524 676240
rect 364518 676200 364524 676212
rect 364576 676200 364582 676252
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 320082 673480 320088 673532
rect 320140 673520 320146 673532
rect 580166 673520 580172 673532
rect 320140 673492 580172 673520
rect 320140 673480 320146 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 386414 667944 386420 667956
rect 3476 667916 386420 667944
rect 3476 667904 3482 667916
rect 386414 667904 386420 667916
rect 386472 667904 386478 667956
rect 429565 666587 429623 666593
rect 429565 666553 429577 666587
rect 429611 666584 429623 666587
rect 429654 666584 429660 666596
rect 429611 666556 429660 666584
rect 429611 666553 429623 666556
rect 429565 666547 429623 666553
rect 429654 666544 429660 666556
rect 429712 666544 429718 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 383654 652780 383660 652792
rect 3108 652752 383660 652780
rect 3108 652740 3114 652752
rect 383654 652740 383660 652752
rect 383712 652740 383718 652792
rect 315942 650020 315948 650072
rect 316000 650060 316006 650072
rect 580166 650060 580172 650072
rect 316000 650032 580172 650060
rect 316000 650020 316006 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 429378 647232 429384 647284
rect 429436 647272 429442 647284
rect 429470 647272 429476 647284
rect 429436 647244 429476 647272
rect 429436 647232 429442 647244
rect 429470 647232 429476 647244
rect 429528 647232 429534 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 429378 640364 429384 640416
rect 429436 640404 429442 640416
rect 429470 640404 429476 640416
rect 429436 640376 429476 640404
rect 429436 640364 429442 640376
rect 429470 640364 429476 640376
rect 429528 640364 429534 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 317322 638936 317328 638988
rect 317380 638976 317386 638988
rect 580166 638976 580172 638988
rect 317380 638948 580172 638976
rect 317380 638936 317386 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 429286 630640 429292 630692
rect 429344 630680 429350 630692
rect 429470 630680 429476 630692
rect 429344 630652 429476 630680
rect 429344 630640 429350 630652
rect 429470 630640 429476 630652
rect 429528 630640 429534 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 313182 626560 313188 626612
rect 313240 626600 313246 626612
rect 580166 626600 580172 626612
rect 313240 626572 580172 626600
rect 313240 626560 313246 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 387794 623812 387800 623824
rect 3476 623784 387800 623812
rect 3476 623772 3482 623784
rect 387794 623772 387800 623784
rect 387852 623772 387858 623824
rect 364521 618239 364579 618245
rect 364521 618205 364533 618239
rect 364567 618236 364579 618239
rect 364610 618236 364616 618248
rect 364567 618208 364616 618236
rect 364567 618205 364579 618208
rect 364521 618199 364579 618205
rect 364610 618196 364616 618208
rect 364668 618196 364674 618248
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 429286 611328 429292 611380
rect 429344 611368 429350 611380
rect 429470 611368 429476 611380
rect 429344 611340 429476 611368
rect 429344 611328 429350 611340
rect 429470 611328 429476 611340
rect 429528 611328 429534 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 391934 610008 391940 610020
rect 3476 609980 391940 610008
rect 3476 609968 3482 609980
rect 391934 609968 391940 609980
rect 391992 609968 391998 610020
rect 364518 608648 364524 608660
rect 364479 608620 364524 608648
rect 364518 608608 364524 608620
rect 364576 608608 364582 608660
rect 429378 608580 429384 608592
rect 429339 608552 429384 608580
rect 429378 608540 429384 608552
rect 429436 608540 429442 608592
rect 559098 608580 559104 608592
rect 559059 608552 559104 608580
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 309042 603100 309048 603152
rect 309100 603140 309106 603152
rect 580166 603140 580172 603152
rect 309100 603112 580172 603140
rect 309100 603100 309106 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 429381 601715 429439 601721
rect 429381 601681 429393 601715
rect 429427 601712 429439 601715
rect 429562 601712 429568 601724
rect 429427 601684 429568 601712
rect 429427 601681 429439 601684
rect 429381 601675 429439 601681
rect 429562 601672 429568 601684
rect 429620 601672 429626 601724
rect 559101 601715 559159 601721
rect 559101 601681 559113 601715
rect 559147 601712 559159 601715
rect 559282 601712 559288 601724
rect 559147 601684 559288 601712
rect 559147 601681 559159 601684
rect 559101 601675 559159 601681
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 364610 598924 364616 598936
rect 364571 598896 364616 598924
rect 364610 598884 364616 598896
rect 364668 598884 364674 598936
rect 429562 598924 429568 598936
rect 429523 598896 429568 598924
rect 429562 598884 429568 598896
rect 429620 598884 429626 598936
rect 559282 598924 559288 598936
rect 559243 598896 559288 598924
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 390554 594844 390560 594856
rect 3292 594816 390560 594844
rect 3292 594804 3298 594816
rect 390554 594804 390560 594816
rect 390612 594804 390618 594856
rect 311802 592016 311808 592068
rect 311860 592056 311866 592068
rect 580166 592056 580172 592068
rect 311860 592028 580172 592056
rect 311860 592016 311866 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 364613 589339 364671 589345
rect 364613 589305 364625 589339
rect 364659 589336 364671 589339
rect 364702 589336 364708 589348
rect 364659 589308 364708 589336
rect 364659 589305 364671 589308
rect 364613 589299 364671 589305
rect 364702 589296 364708 589308
rect 364760 589296 364766 589348
rect 429565 589339 429623 589345
rect 429565 589305 429577 589339
rect 429611 589336 429623 589339
rect 429654 589336 429660 589348
rect 429611 589308 429660 589336
rect 429611 589305 429623 589308
rect 429565 589299 429623 589305
rect 429654 589296 429660 589308
rect 429712 589296 429718 589348
rect 559285 589339 559343 589345
rect 559285 589305 559297 589339
rect 559331 589336 559343 589339
rect 559374 589336 559380 589348
rect 559331 589308 559380 589336
rect 559331 589305 559343 589308
rect 559285 589299 559343 589305
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 344462 584672 344468 584724
rect 344520 584712 344526 584724
rect 364702 584712 364708 584724
rect 344520 584684 364708 584712
rect 344520 584672 344526 584684
rect 364702 584672 364708 584684
rect 364760 584672 364766 584724
rect 300762 584604 300768 584656
rect 300820 584644 300826 584656
rect 350810 584644 350816 584656
rect 300820 584616 350816 584644
rect 300820 584604 300826 584616
rect 350810 584604 350816 584616
rect 350868 584604 350874 584656
rect 338206 584536 338212 584588
rect 338264 584576 338270 584588
rect 429654 584576 429660 584588
rect 338264 584548 429660 584576
rect 338264 584536 338270 584548
rect 429654 584536 429660 584548
rect 429712 584536 429718 584588
rect 331858 584468 331864 584520
rect 331916 584508 331922 584520
rect 494238 584508 494244 584520
rect 331916 584480 494244 584508
rect 331916 584468 331922 584480
rect 494238 584468 494244 584480
rect 494296 584468 494302 584520
rect 325510 584400 325516 584452
rect 325568 584440 325574 584452
rect 559374 584440 559380 584452
rect 325568 584412 559380 584440
rect 325568 584400 325574 584412
rect 559374 584400 559380 584412
rect 559432 584400 559438 584452
rect 298186 583652 298192 583704
rect 298244 583692 298250 583704
rect 471238 583692 471244 583704
rect 298244 583664 471244 583692
rect 298244 583652 298250 583664
rect 471238 583652 471244 583664
rect 471296 583652 471302 583704
rect 256050 583584 256056 583636
rect 256108 583624 256114 583636
rect 580534 583624 580540 583636
rect 256108 583596 580540 583624
rect 256108 583584 256114 583596
rect 580534 583584 580540 583596
rect 580592 583584 580598 583636
rect 245562 583516 245568 583568
rect 245620 583556 245626 583568
rect 580258 583556 580264 583568
rect 245620 583528 580264 583556
rect 245620 583516 245626 583528
rect 580258 583516 580264 583528
rect 580316 583516 580322 583568
rect 6638 583448 6644 583500
rect 6696 583488 6702 583500
rect 399202 583488 399208 583500
rect 6696 583460 399208 583488
rect 6696 583448 6702 583460
rect 399202 583448 399208 583460
rect 399260 583448 399266 583500
rect 4706 583380 4712 583432
rect 4764 583420 4770 583432
rect 405550 583420 405556 583432
rect 4764 583392 405556 583420
rect 4764 583380 4770 583392
rect 405550 583380 405556 583392
rect 405608 583380 405614 583432
rect 10318 583312 10324 583364
rect 10376 583352 10382 583364
rect 411898 583352 411904 583364
rect 10376 583324 411904 583352
rect 10376 583312 10382 583324
rect 411898 583312 411904 583324
rect 411956 583312 411962 583364
rect 6270 583244 6276 583296
rect 6328 583284 6334 583296
rect 409782 583284 409788 583296
rect 6328 583256 409788 583284
rect 6328 583244 6334 583256
rect 409782 583244 409788 583256
rect 409840 583244 409846 583296
rect 3142 583176 3148 583228
rect 3200 583216 3206 583228
rect 407666 583216 407672 583228
rect 3200 583188 407672 583216
rect 3200 583176 3206 583188
rect 407666 583176 407672 583188
rect 407724 583176 407730 583228
rect 13078 583108 13084 583160
rect 13136 583148 13142 583160
rect 418154 583148 418160 583160
rect 13136 583120 418160 583148
rect 13136 583108 13142 583120
rect 418154 583108 418160 583120
rect 418212 583108 418218 583160
rect 14458 583040 14464 583092
rect 14516 583080 14522 583092
rect 424502 583080 424508 583092
rect 14516 583052 424508 583080
rect 14516 583040 14522 583052
rect 424502 583040 424508 583052
rect 424560 583040 424566 583092
rect 3234 582972 3240 583024
rect 3292 583012 3298 583024
rect 414014 583012 414020 583024
rect 3292 582984 414020 583012
rect 3292 582972 3298 582984
rect 414014 582972 414020 582984
rect 414072 582972 414078 583024
rect 5442 582904 5448 582956
rect 5500 582944 5506 582956
rect 422386 582944 422392 582956
rect 5500 582916 422392 582944
rect 5500 582904 5506 582916
rect 422386 582904 422392 582916
rect 422444 582904 422450 582956
rect 15838 582836 15844 582888
rect 15896 582876 15902 582888
rect 437106 582876 437112 582888
rect 15896 582848 437112 582876
rect 15896 582836 15902 582848
rect 437106 582836 437112 582848
rect 437164 582836 437170 582888
rect 4062 582768 4068 582820
rect 4120 582808 4126 582820
rect 430850 582808 430856 582820
rect 4120 582780 430856 582808
rect 4120 582768 4126 582780
rect 430850 582768 430856 582780
rect 430908 582768 430914 582820
rect 5350 582700 5356 582752
rect 5408 582740 5414 582752
rect 432966 582740 432972 582752
rect 5408 582712 432972 582740
rect 5408 582700 5414 582712
rect 432966 582700 432972 582712
rect 433024 582700 433030 582752
rect 3878 582632 3884 582684
rect 3936 582672 3942 582684
rect 434990 582672 434996 582684
rect 3936 582644 434996 582672
rect 3936 582632 3942 582644
rect 434990 582632 434996 582644
rect 435048 582632 435054 582684
rect 17218 582564 17224 582616
rect 17276 582604 17282 582616
rect 449802 582604 449808 582616
rect 17276 582576 449808 582604
rect 17276 582564 17282 582576
rect 449802 582564 449808 582576
rect 449860 582564 449866 582616
rect 5258 582496 5264 582548
rect 5316 582536 5322 582548
rect 445570 582536 445576 582548
rect 5316 582508 445576 582536
rect 5316 582496 5322 582508
rect 445570 582496 445576 582508
rect 445628 582496 445634 582548
rect 3694 582428 3700 582480
rect 3752 582468 3758 582480
rect 443454 582468 443460 582480
rect 3752 582440 443460 582468
rect 3752 582428 3758 582440
rect 443454 582428 443460 582440
rect 443512 582428 443518 582480
rect 5166 582360 5172 582412
rect 5224 582400 5230 582412
rect 447686 582400 447692 582412
rect 5224 582372 447692 582400
rect 5224 582360 5230 582372
rect 447686 582360 447692 582372
rect 447744 582360 447750 582412
rect 302418 581680 302424 581732
rect 302476 581720 302482 581732
rect 469582 581720 469588 581732
rect 302476 581692 469588 581720
rect 302476 581680 302482 581692
rect 469582 581680 469588 581692
rect 469640 581680 469646 581732
rect 296070 581612 296076 581664
rect 296128 581652 296134 581664
rect 469766 581652 469772 581664
rect 296128 581624 469772 581652
rect 296128 581612 296134 581624
rect 469766 581612 469772 581624
rect 469824 581612 469830 581664
rect 289722 581544 289728 581596
rect 289780 581584 289786 581596
rect 470502 581584 470508 581596
rect 289780 581556 470508 581584
rect 289780 581544 289786 581556
rect 470502 581544 470508 581556
rect 470560 581544 470566 581596
rect 287606 581476 287612 581528
rect 287664 581516 287670 581528
rect 470410 581516 470416 581528
rect 287664 581488 470416 581516
rect 287664 581476 287670 581488
rect 470410 581476 470416 581488
rect 470468 581476 470474 581528
rect 283466 581408 283472 581460
rect 283524 581448 283530 581460
rect 470318 581448 470324 581460
rect 283524 581420 470324 581448
rect 283524 581408 283530 581420
rect 470318 581408 470324 581420
rect 470376 581408 470382 581460
rect 281350 581340 281356 581392
rect 281408 581380 281414 581392
rect 470226 581380 470232 581392
rect 281408 581352 470232 581380
rect 281408 581340 281414 581352
rect 470226 581340 470232 581352
rect 470284 581340 470290 581392
rect 275002 581272 275008 581324
rect 275060 581312 275066 581324
rect 470134 581312 470140 581324
rect 275060 581284 470140 581312
rect 275060 581272 275066 581284
rect 470134 581272 470140 581284
rect 470192 581272 470198 581324
rect 268654 581204 268660 581256
rect 268712 581244 268718 581256
rect 469950 581244 469956 581256
rect 268712 581216 469956 581244
rect 268712 581204 268718 581216
rect 469950 581204 469956 581216
rect 470008 581204 470014 581256
rect 304534 581136 304540 581188
rect 304592 581176 304598 581188
rect 552658 581176 552664 581188
rect 304592 581148 552664 581176
rect 304592 581136 304598 581148
rect 552658 581136 552664 581148
rect 552716 581136 552722 581188
rect 264514 581068 264520 581120
rect 264572 581108 264578 581120
rect 580902 581108 580908 581120
rect 264572 581080 580908 581108
rect 264572 581068 264578 581080
rect 580902 581068 580908 581080
rect 580960 581068 580966 581120
rect 4798 581000 4804 581052
rect 4856 581040 4862 581052
rect 466638 581040 466644 581052
rect 4856 581012 466644 581040
rect 4856 581000 4862 581012
rect 466638 581000 466644 581012
rect 466696 581000 466702 581052
rect 300302 580320 300308 580372
rect 300360 580360 300366 580372
rect 469674 580360 469680 580372
rect 300360 580332 469680 580360
rect 300360 580320 300366 580332
rect 469674 580320 469680 580332
rect 469732 580320 469738 580372
rect 262398 580252 262404 580304
rect 262456 580292 262462 580304
rect 469858 580292 469864 580304
rect 262456 580264 469864 580292
rect 262456 580252 262462 580264
rect 469858 580252 469864 580264
rect 469916 580252 469922 580304
rect 306558 580184 306564 580236
rect 306616 580224 306622 580236
rect 580166 580224 580172 580236
rect 306616 580196 580172 580224
rect 306616 580184 306622 580196
rect 580166 580184 580172 580196
rect 580224 580184 580230 580236
rect 6730 580116 6736 580168
rect 6788 580156 6794 580168
rect 395062 580156 395068 580168
rect 6788 580128 395068 580156
rect 6788 580116 6794 580128
rect 395062 580116 395068 580128
rect 395120 580116 395126 580168
rect 6546 580048 6552 580100
rect 6604 580088 6610 580100
rect 397086 580088 397092 580100
rect 6604 580060 397092 580088
rect 6604 580048 6610 580060
rect 397086 580048 397092 580060
rect 397144 580048 397150 580100
rect 6454 579980 6460 580032
rect 6512 580020 6518 580032
rect 400950 580020 400956 580032
rect 6512 579992 400956 580020
rect 6512 579980 6518 579992
rect 400950 579980 400956 579992
rect 401008 579980 401014 580032
rect 6362 579912 6368 579964
rect 6420 579952 6426 579964
rect 403158 579952 403164 579964
rect 6420 579924 403164 579952
rect 6420 579912 6426 579924
rect 403158 579912 403164 579924
rect 403216 579912 403222 579964
rect 3786 579844 3792 579896
rect 3844 579884 3850 579896
rect 438854 579884 438860 579896
rect 3844 579856 438860 579884
rect 3844 579844 3850 579856
rect 438854 579844 438860 579856
rect 438912 579844 438918 579896
rect 5074 579776 5080 579828
rect 5132 579816 5138 579828
rect 451550 579816 451556 579828
rect 5132 579788 451556 579816
rect 5132 579776 5138 579788
rect 451550 579776 451556 579788
rect 451608 579776 451614 579828
rect 4982 579708 4988 579760
rect 5040 579748 5046 579760
rect 458266 579748 458272 579760
rect 5040 579720 458272 579748
rect 5040 579708 5046 579720
rect 458266 579708 458272 579720
rect 458324 579708 458330 579760
rect 6178 579640 6184 579692
rect 6236 579680 6242 579692
rect 464246 579680 464252 579692
rect 6236 579652 464252 579680
rect 6236 579640 6242 579652
rect 464246 579640 464252 579652
rect 464304 579640 464310 579692
rect 289725 579615 289783 579621
rect 289725 579612 289737 579615
rect 282196 579584 289737 579612
rect 282196 579476 282224 579584
rect 289725 579581 289737 579584
rect 289771 579581 289783 579615
rect 289725 579575 289783 579581
rect 454037 579615 454095 579621
rect 454037 579581 454049 579615
rect 454083 579612 454095 579615
rect 463605 579615 463663 579621
rect 463605 579612 463617 579615
rect 454083 579584 463617 579612
rect 454083 579581 454095 579584
rect 454037 579575 454095 579581
rect 463605 579581 463617 579584
rect 463651 579581 463663 579615
rect 463605 579575 463663 579581
rect 289909 579547 289967 579553
rect 289909 579513 289921 579547
rect 289955 579544 289967 579547
rect 289955 579516 294552 579544
rect 289955 579513 289967 579516
rect 289909 579507 289967 579513
rect 275480 579448 282224 579476
rect 289725 579479 289783 579485
rect 271138 579368 271144 579420
rect 271196 579408 271202 579420
rect 271196 579380 273208 579408
rect 271196 579368 271202 579380
rect 252094 579340 252100 579352
rect 252055 579312 252100 579340
rect 252094 579300 252100 579312
rect 252152 579300 252158 579352
rect 254210 579340 254216 579352
rect 254171 579312 254216 579340
rect 254210 579300 254216 579312
rect 254268 579300 254274 579352
rect 258442 579300 258448 579352
rect 258500 579300 258506 579352
rect 260650 579300 260656 579352
rect 260708 579300 260714 579352
rect 266906 579300 266912 579352
rect 266964 579300 266970 579352
rect 273070 579300 273076 579352
rect 273128 579300 273134 579352
rect 273180 579340 273208 579380
rect 275480 579340 275508 579448
rect 289725 579445 289737 579479
rect 289771 579476 289783 579479
rect 289817 579479 289875 579485
rect 289817 579476 289829 579479
rect 289771 579448 289829 579476
rect 289771 579445 289783 579448
rect 289725 579439 289783 579445
rect 289817 579445 289829 579448
rect 289863 579445 289875 579479
rect 289817 579439 289875 579445
rect 273180 579312 275508 579340
rect 277302 579300 277308 579352
rect 277360 579300 277366 579352
rect 279602 579300 279608 579352
rect 279660 579300 279666 579352
rect 285674 579300 285680 579352
rect 285732 579300 285738 579352
rect 292114 579300 292120 579352
rect 292172 579300 292178 579352
rect 258460 578728 258488 579300
rect 260668 578796 260696 579300
rect 266924 578864 266952 579300
rect 273088 578932 273116 579300
rect 277320 579000 277348 579300
rect 279620 579068 279648 579300
rect 285692 579136 285720 579300
rect 292132 579204 292160 579300
rect 294524 579272 294552 579516
rect 318797 579479 318855 579485
rect 318797 579445 318809 579479
rect 318843 579476 318855 579479
rect 328365 579479 328423 579485
rect 328365 579476 328377 579479
rect 318843 579448 328377 579476
rect 318843 579445 318855 579448
rect 318797 579439 318855 579445
rect 328365 579445 328377 579448
rect 328411 579445 328423 579479
rect 328365 579439 328423 579445
rect 338117 579479 338175 579485
rect 338117 579445 338129 579479
rect 338163 579476 338175 579479
rect 347685 579479 347743 579485
rect 347685 579476 347697 579479
rect 338163 579448 347697 579476
rect 338163 579445 338175 579448
rect 338117 579439 338175 579445
rect 347685 579445 347697 579448
rect 347731 579445 347743 579479
rect 347685 579439 347743 579445
rect 357437 579479 357495 579485
rect 357437 579445 357449 579479
rect 357483 579476 357495 579479
rect 367005 579479 367063 579485
rect 367005 579476 367017 579479
rect 357483 579448 367017 579476
rect 357483 579445 357495 579448
rect 357437 579439 357495 579445
rect 367005 579445 367017 579448
rect 367051 579445 367063 579479
rect 367005 579439 367063 579445
rect 376757 579479 376815 579485
rect 376757 579445 376769 579479
rect 376803 579476 376815 579479
rect 386325 579479 386383 579485
rect 386325 579476 386337 579479
rect 376803 579448 386337 579476
rect 376803 579445 376815 579448
rect 376757 579439 376815 579445
rect 386325 579445 386337 579448
rect 386371 579445 386383 579479
rect 386325 579439 386383 579445
rect 396077 579479 396135 579485
rect 396077 579445 396089 579479
rect 396123 579476 396135 579479
rect 405645 579479 405703 579485
rect 405645 579476 405657 579479
rect 396123 579448 405657 579476
rect 396123 579445 396135 579448
rect 396077 579439 396135 579445
rect 405645 579445 405657 579448
rect 405691 579445 405703 579479
rect 405645 579439 405703 579445
rect 408497 579479 408555 579485
rect 408497 579445 408509 579479
rect 408543 579476 408555 579479
rect 415305 579479 415363 579485
rect 415305 579476 415317 579479
rect 408543 579448 415317 579476
rect 408543 579445 408555 579448
rect 408497 579439 408555 579445
rect 415305 579445 415317 579448
rect 415351 579445 415363 579479
rect 444285 579479 444343 579485
rect 444285 579476 444297 579479
rect 415305 579439 415363 579445
rect 435744 579448 444297 579476
rect 415670 579408 415676 579420
rect 415631 579380 415676 579408
rect 415670 579368 415676 579380
rect 415728 579368 415734 579420
rect 428366 579408 428372 579420
rect 428327 579380 428372 579408
rect 428366 579368 428372 579380
rect 428424 579368 428430 579420
rect 294601 579343 294659 579349
rect 294601 579309 294613 579343
rect 294647 579340 294659 579343
rect 299293 579343 299351 579349
rect 299293 579340 299305 579343
rect 294647 579312 299305 579340
rect 294647 579309 294659 579312
rect 294601 579303 294659 579309
rect 299293 579309 299305 579312
rect 299339 579309 299351 579343
rect 299293 579303 299351 579309
rect 311989 579343 312047 579349
rect 311989 579309 312001 579343
rect 312035 579340 312047 579343
rect 318797 579343 318855 579349
rect 318797 579340 318809 579343
rect 312035 579312 318809 579340
rect 312035 579309 312047 579312
rect 311989 579303 312047 579309
rect 318797 579309 318809 579312
rect 318843 579309 318855 579343
rect 318797 579303 318855 579309
rect 331309 579343 331367 579349
rect 331309 579309 331321 579343
rect 331355 579340 331367 579343
rect 338117 579343 338175 579349
rect 338117 579340 338129 579343
rect 331355 579312 338129 579340
rect 331355 579309 331367 579312
rect 331309 579303 331367 579309
rect 338117 579309 338129 579312
rect 338163 579309 338175 579343
rect 338117 579303 338175 579309
rect 350629 579343 350687 579349
rect 350629 579309 350641 579343
rect 350675 579340 350687 579343
rect 357437 579343 357495 579349
rect 357437 579340 357449 579343
rect 350675 579312 357449 579340
rect 350675 579309 350687 579312
rect 350629 579303 350687 579309
rect 357437 579309 357449 579312
rect 357483 579309 357495 579343
rect 357437 579303 357495 579309
rect 369949 579343 370007 579349
rect 369949 579309 369961 579343
rect 369995 579340 370007 579343
rect 376757 579343 376815 579349
rect 376757 579340 376769 579343
rect 369995 579312 376769 579340
rect 369995 579309 370007 579312
rect 369949 579303 370007 579309
rect 376757 579309 376769 579312
rect 376803 579309 376815 579343
rect 376757 579303 376815 579309
rect 389269 579343 389327 579349
rect 389269 579309 389281 579343
rect 389315 579340 389327 579343
rect 396077 579343 396135 579349
rect 396077 579340 396089 579343
rect 389315 579312 396089 579340
rect 389315 579309 389327 579312
rect 389269 579303 389327 579309
rect 396077 579309 396089 579312
rect 396123 579309 396135 579343
rect 396077 579303 396135 579309
rect 415305 579343 415363 579349
rect 415305 579309 415317 579343
rect 415351 579340 415363 579343
rect 435744 579340 435772 579448
rect 444285 579445 444297 579448
rect 444331 579445 444343 579479
rect 444285 579439 444343 579445
rect 444377 579479 444435 579485
rect 444377 579445 444389 579479
rect 444423 579476 444435 579479
rect 454037 579479 454095 579485
rect 454037 579476 454049 579479
rect 444423 579448 454049 579476
rect 444423 579445 444435 579448
rect 444377 579439 444435 579445
rect 454037 579445 454049 579448
rect 454083 579445 454095 579479
rect 454037 579439 454095 579445
rect 453574 579408 453580 579420
rect 453535 579380 453580 579408
rect 453574 579368 453580 579380
rect 453632 579368 453638 579420
rect 455782 579408 455788 579420
rect 455743 579380 455788 579408
rect 455782 579368 455788 579380
rect 455840 579368 455846 579420
rect 441062 579340 441068 579352
rect 415351 579312 418200 579340
rect 415351 579309 415363 579312
rect 415305 579303 415363 579309
rect 311805 579275 311863 579281
rect 311805 579272 311817 579275
rect 294524 579244 311817 579272
rect 311805 579241 311817 579244
rect 311851 579241 311863 579275
rect 311805 579235 311863 579241
rect 328365 579275 328423 579281
rect 328365 579241 328377 579275
rect 328411 579272 328423 579275
rect 331125 579275 331183 579281
rect 331125 579272 331137 579275
rect 328411 579244 331137 579272
rect 328411 579241 328423 579244
rect 328365 579235 328423 579241
rect 331125 579241 331137 579244
rect 331171 579241 331183 579275
rect 331125 579235 331183 579241
rect 347685 579275 347743 579281
rect 347685 579241 347697 579275
rect 347731 579272 347743 579275
rect 350445 579275 350503 579281
rect 350445 579272 350457 579275
rect 347731 579244 350457 579272
rect 347731 579241 347743 579244
rect 347685 579235 347743 579241
rect 350445 579241 350457 579244
rect 350491 579241 350503 579275
rect 350445 579235 350503 579241
rect 367005 579275 367063 579281
rect 367005 579241 367017 579275
rect 367051 579272 367063 579275
rect 369765 579275 369823 579281
rect 369765 579272 369777 579275
rect 367051 579244 369777 579272
rect 367051 579241 367063 579244
rect 367005 579235 367063 579241
rect 369765 579241 369777 579244
rect 369811 579241 369823 579275
rect 369765 579235 369823 579241
rect 386325 579275 386383 579281
rect 386325 579241 386337 579275
rect 386371 579272 386383 579275
rect 389085 579275 389143 579281
rect 389085 579272 389097 579275
rect 386371 579244 389097 579272
rect 386371 579241 386383 579244
rect 386325 579235 386383 579241
rect 389085 579241 389097 579244
rect 389131 579241 389143 579275
rect 389085 579235 389143 579241
rect 405645 579275 405703 579281
rect 405645 579241 405657 579275
rect 405691 579272 405703 579275
rect 408497 579275 408555 579281
rect 408497 579272 408509 579275
rect 405691 579244 408509 579272
rect 405691 579241 405703 579244
rect 405645 579235 405703 579241
rect 408497 579241 408509 579244
rect 408543 579241 408555 579275
rect 418172 579272 418200 579312
rect 427832 579312 435772 579340
rect 441023 579312 441068 579340
rect 427832 579272 427860 579312
rect 441062 579300 441068 579312
rect 441120 579300 441126 579352
rect 463605 579343 463663 579349
rect 463605 579309 463617 579343
rect 463651 579340 463663 579343
rect 464433 579343 464491 579349
rect 464433 579340 464445 579343
rect 463651 579312 464445 579340
rect 463651 579309 463663 579312
rect 463605 579303 463663 579309
rect 464433 579309 464445 579312
rect 464479 579309 464491 579343
rect 464433 579303 464491 579309
rect 418172 579244 427860 579272
rect 444285 579275 444343 579281
rect 408497 579235 408555 579241
rect 444285 579241 444297 579275
rect 444331 579272 444343 579275
rect 444377 579275 444435 579281
rect 444377 579272 444389 579275
rect 444331 579244 444389 579272
rect 444331 579241 444343 579244
rect 444285 579235 444343 579241
rect 444377 579241 444389 579244
rect 444423 579241 444435 579275
rect 444377 579235 444435 579241
rect 579798 579204 579804 579216
rect 292132 579176 579804 579204
rect 579798 579164 579804 579176
rect 579856 579164 579862 579216
rect 579890 579136 579896 579148
rect 285692 579108 579896 579136
rect 579890 579096 579896 579108
rect 579948 579096 579954 579148
rect 580074 579068 580080 579080
rect 279620 579040 580080 579068
rect 580074 579028 580080 579040
rect 580132 579028 580138 579080
rect 294601 579003 294659 579009
rect 294601 579000 294613 579003
rect 277320 578972 294613 579000
rect 294601 578969 294613 578972
rect 294647 578969 294659 579003
rect 299293 579003 299351 579009
rect 294601 578963 294659 578969
rect 294708 578972 299244 579000
rect 294708 578932 294736 578972
rect 273088 578904 294736 578932
rect 299216 578932 299244 578972
rect 299293 578969 299305 579003
rect 299339 579000 299351 579003
rect 579982 579000 579988 579012
rect 299339 578972 579988 579000
rect 299339 578969 299351 578972
rect 299293 578963 299351 578969
rect 579982 578960 579988 578972
rect 580040 578960 580046 579012
rect 580166 578932 580172 578944
rect 299216 578904 580172 578932
rect 580166 578892 580172 578904
rect 580224 578892 580230 578944
rect 299109 578867 299167 578873
rect 299109 578864 299121 578867
rect 266924 578836 299121 578864
rect 299109 578833 299121 578836
rect 299155 578833 299167 578867
rect 299109 578827 299167 578833
rect 299385 578867 299443 578873
rect 299385 578833 299397 578867
rect 299431 578864 299443 578867
rect 580810 578864 580816 578876
rect 299431 578836 580816 578864
rect 299431 578833 299443 578836
rect 299385 578827 299443 578833
rect 580810 578824 580816 578836
rect 580868 578824 580874 578876
rect 299201 578799 299259 578805
rect 299201 578796 299213 578799
rect 260668 578768 299213 578796
rect 299201 578765 299213 578768
rect 299247 578765 299259 578799
rect 299201 578759 299259 578765
rect 299293 578799 299351 578805
rect 299293 578765 299305 578799
rect 299339 578796 299351 578799
rect 580626 578796 580632 578808
rect 299339 578768 580632 578796
rect 299339 578765 299351 578768
rect 299293 578759 299351 578765
rect 580626 578756 580632 578768
rect 580684 578756 580690 578808
rect 580718 578728 580724 578740
rect 258460 578700 580724 578728
rect 580718 578688 580724 578700
rect 580776 578688 580782 578740
rect 254213 578663 254271 578669
rect 254213 578629 254225 578663
rect 254259 578660 254271 578663
rect 299109 578663 299167 578669
rect 299109 578660 299121 578663
rect 254259 578632 299121 578660
rect 254259 578629 254271 578632
rect 254213 578623 254271 578629
rect 299109 578629 299121 578632
rect 299155 578629 299167 578663
rect 299109 578623 299167 578629
rect 299293 578663 299351 578669
rect 299293 578629 299305 578663
rect 299339 578660 299351 578663
rect 580350 578660 580356 578672
rect 299339 578632 580356 578660
rect 299339 578629 299351 578632
rect 299293 578623 299351 578629
rect 580350 578620 580356 578632
rect 580408 578620 580414 578672
rect 252097 578595 252155 578601
rect 252097 578561 252109 578595
rect 252143 578592 252155 578595
rect 299017 578595 299075 578601
rect 299017 578592 299029 578595
rect 252143 578564 299029 578592
rect 252143 578561 252155 578564
rect 252097 578555 252155 578561
rect 299017 578561 299029 578564
rect 299063 578561 299075 578595
rect 299017 578555 299075 578561
rect 299201 578595 299259 578601
rect 299201 578561 299213 578595
rect 299247 578592 299259 578595
rect 580442 578592 580448 578604
rect 299247 578564 580448 578592
rect 299247 578561 299259 578564
rect 299201 578555 299259 578561
rect 580442 578552 580448 578564
rect 580500 578552 580506 578604
rect 3326 578484 3332 578536
rect 3384 578524 3390 578536
rect 298925 578527 298983 578533
rect 298925 578524 298937 578527
rect 3384 578496 298937 578524
rect 3384 578484 3390 578496
rect 298925 578493 298937 578496
rect 298971 578493 298983 578527
rect 298925 578487 298983 578493
rect 299109 578527 299167 578533
rect 299109 578493 299121 578527
rect 299155 578524 299167 578527
rect 415673 578527 415731 578533
rect 415673 578524 415685 578527
rect 299155 578496 415685 578524
rect 299155 578493 299167 578496
rect 299109 578487 299167 578493
rect 415673 578493 415685 578496
rect 415719 578493 415731 578527
rect 415673 578487 415731 578493
rect 3970 578416 3976 578468
rect 4028 578456 4034 578468
rect 428369 578459 428427 578465
rect 428369 578456 428381 578459
rect 4028 578428 428381 578456
rect 4028 578416 4034 578428
rect 428369 578425 428381 578428
rect 428415 578425 428427 578459
rect 428369 578419 428427 578425
rect 3602 578348 3608 578400
rect 3660 578388 3666 578400
rect 441065 578391 441123 578397
rect 441065 578388 441077 578391
rect 3660 578360 441077 578388
rect 3660 578348 3666 578360
rect 441065 578357 441077 578360
rect 441111 578357 441123 578391
rect 441065 578351 441123 578357
rect 3418 578280 3424 578332
rect 3476 578320 3482 578332
rect 453577 578323 453635 578329
rect 453577 578320 453589 578323
rect 3476 578292 453589 578320
rect 3476 578280 3482 578292
rect 453577 578289 453589 578292
rect 453623 578289 453635 578323
rect 453577 578283 453635 578289
rect 3510 578212 3516 578264
rect 3568 578252 3574 578264
rect 455785 578255 455843 578261
rect 455785 578252 455797 578255
rect 3568 578224 455797 578252
rect 3568 578212 3574 578224
rect 455785 578221 455797 578224
rect 455831 578221 455843 578255
rect 455785 578215 455843 578221
rect 464433 577915 464491 577921
rect 464433 577881 464445 577915
rect 464479 577912 464491 577915
rect 470042 577912 470048 577924
rect 464479 577884 470048 577912
rect 464479 577881 464491 577884
rect 464433 577875 464491 577881
rect 470042 577872 470048 577884
rect 470100 577872 470106 577924
rect 3050 568284 3056 568336
rect 3108 568324 3114 568336
rect 6730 568324 6736 568336
rect 3108 568296 6736 568324
rect 3108 568284 3114 568296
rect 6730 568284 6736 568296
rect 6788 568284 6794 568336
rect 579706 567128 579712 567180
rect 579764 567168 579770 567180
rect 580902 567168 580908 567180
rect 579764 567140 580908 567168
rect 579764 567128 579770 567140
rect 580902 567128 580908 567140
rect 580960 567128 580966 567180
rect 579706 557608 579712 557660
rect 579764 557648 579770 557660
rect 579764 557620 580948 557648
rect 579764 557608 579770 557620
rect 580920 557592 580948 557620
rect 580902 557540 580908 557592
rect 580960 557540 580966 557592
rect 469582 557472 469588 557524
rect 469640 557512 469646 557524
rect 579706 557512 579712 557524
rect 469640 557484 579712 557512
rect 469640 557472 469646 557484
rect 579706 557472 579712 557484
rect 579764 557472 579770 557524
rect 3050 553324 3056 553376
rect 3108 553364 3114 553376
rect 6638 553364 6644 553376
rect 3108 553336 6644 553364
rect 3108 553324 3114 553336
rect 6638 553324 6644 553336
rect 6696 553324 6702 553376
rect 579614 547816 579620 547868
rect 579672 547856 579678 547868
rect 580902 547856 580908 547868
rect 579672 547828 580908 547856
rect 579672 547816 579678 547828
rect 580902 547816 580908 547828
rect 580960 547816 580966 547868
rect 552658 546388 552664 546440
rect 552716 546428 552722 546440
rect 579706 546428 579712 546440
rect 552716 546400 579712 546428
rect 552716 546388 552722 546400
rect 579706 546388 579712 546400
rect 579764 546388 579770 546440
rect 3050 538636 3056 538688
rect 3108 538676 3114 538688
rect 6546 538676 6552 538688
rect 3108 538648 6552 538676
rect 3108 538636 3114 538648
rect 6546 538636 6552 538648
rect 6604 538636 6610 538688
rect 579614 538228 579620 538280
rect 579672 538268 579678 538280
rect 580902 538268 580908 538280
rect 579672 538240 580908 538268
rect 579672 538228 579678 538240
rect 580902 538228 580908 538240
rect 580960 538228 580966 538280
rect 469674 534012 469680 534064
rect 469732 534052 469738 534064
rect 579706 534052 579712 534064
rect 469732 534024 579712 534052
rect 469732 534012 469738 534024
rect 579706 534012 579712 534024
rect 579764 534012 579770 534064
rect 579706 528504 579712 528556
rect 579764 528544 579770 528556
rect 580902 528544 580908 528556
rect 579764 528516 580908 528544
rect 579764 528504 579770 528516
rect 580902 528504 580908 528516
rect 580960 528504 580966 528556
rect 579706 518916 579712 518968
rect 579764 518956 579770 518968
rect 580902 518956 580908 518968
rect 579764 518928 580908 518956
rect 579764 518916 579770 518928
rect 580902 518916 580908 518928
rect 580960 518916 580966 518968
rect 469766 510552 469772 510604
rect 469824 510592 469830 510604
rect 579706 510592 579712 510604
rect 469824 510564 579712 510592
rect 469824 510552 469830 510564
rect 579706 510552 579712 510564
rect 579764 510552 579770 510604
rect 3050 510212 3056 510264
rect 3108 510252 3114 510264
rect 6454 510252 6460 510264
rect 3108 510224 6460 510252
rect 3108 510212 3114 510224
rect 6454 510212 6460 510224
rect 6512 510212 6518 510264
rect 579706 509192 579712 509244
rect 579764 509232 579770 509244
rect 580902 509232 580908 509244
rect 579764 509204 580908 509232
rect 579764 509192 579770 509204
rect 580902 509192 580908 509204
rect 580960 509192 580966 509244
rect 579706 499604 579712 499656
rect 579764 499644 579770 499656
rect 579764 499616 580948 499644
rect 579764 499604 579770 499616
rect 580920 499588 580948 499616
rect 580902 499536 580908 499588
rect 580960 499536 580966 499588
rect 471238 499468 471244 499520
rect 471296 499508 471302 499520
rect 579706 499508 579712 499520
rect 471296 499480 579712 499508
rect 471296 499468 471302 499480
rect 579706 499468 579712 499480
rect 579764 499468 579770 499520
rect 2774 495524 2780 495576
rect 2832 495564 2838 495576
rect 4706 495564 4712 495576
rect 2832 495536 4712 495564
rect 2832 495524 2838 495536
rect 4706 495524 4712 495536
rect 4764 495524 4770 495576
rect 579706 489812 579712 489864
rect 579764 489852 579770 489864
rect 580902 489852 580908 489864
rect 579764 489824 580908 489852
rect 579764 489812 579770 489824
rect 580902 489812 580908 489824
rect 580960 489812 580966 489864
rect 2958 481108 2964 481160
rect 3016 481148 3022 481160
rect 6362 481148 6368 481160
rect 3016 481120 6368 481148
rect 3016 481108 3022 481120
rect 6362 481108 6368 481120
rect 6420 481108 6426 481160
rect 579706 480224 579712 480276
rect 579764 480264 579770 480276
rect 580902 480264 580908 480276
rect 579764 480236 580908 480264
rect 579764 480224 579770 480236
rect 580902 480224 580908 480236
rect 580960 480224 580966 480276
rect 579614 470500 579620 470552
rect 579672 470540 579678 470552
rect 580902 470540 580908 470552
rect 579672 470512 580908 470540
rect 579672 470500 579678 470512
rect 580902 470500 580908 470512
rect 580960 470500 580966 470552
rect 470502 463632 470508 463684
rect 470560 463672 470566 463684
rect 579706 463672 579712 463684
rect 470560 463644 579712 463672
rect 470560 463632 470566 463644
rect 579706 463632 579712 463644
rect 579764 463632 579770 463684
rect 579614 460912 579620 460964
rect 579672 460952 579678 460964
rect 580902 460952 580908 460964
rect 579672 460924 580908 460952
rect 579672 460912 579678 460924
rect 580902 460912 580908 460924
rect 580960 460912 580966 460964
rect 579798 451188 579804 451240
rect 579856 451228 579862 451240
rect 580902 451228 580908 451240
rect 579856 451200 580908 451228
rect 579856 451188 579862 451200
rect 580902 451188 580908 451200
rect 580960 451188 580966 451240
rect 579798 441600 579804 441652
rect 579856 441640 579862 441652
rect 580902 441640 580908 441652
rect 579856 441612 580908 441640
rect 579856 441600 579862 441612
rect 580902 441600 580908 441612
rect 580960 441600 580966 441652
rect 470410 440172 470416 440224
rect 470468 440212 470474 440224
rect 579798 440212 579804 440224
rect 470468 440184 579804 440212
rect 470468 440172 470474 440184
rect 579798 440172 579804 440184
rect 579856 440172 579862 440224
rect 3142 438812 3148 438864
rect 3200 438852 3206 438864
rect 10318 438852 10324 438864
rect 3200 438824 10324 438852
rect 3200 438812 3206 438824
rect 10318 438812 10324 438824
rect 10376 438812 10382 438864
rect 579798 431876 579804 431928
rect 579856 431916 579862 431928
rect 580902 431916 580908 431928
rect 579856 431888 580908 431916
rect 579856 431876 579862 431888
rect 580902 431876 580908 431888
rect 580960 431876 580966 431928
rect 3142 424056 3148 424108
rect 3200 424096 3206 424108
rect 6270 424096 6276 424108
rect 3200 424068 6276 424096
rect 3200 424056 3206 424068
rect 6270 424056 6276 424068
rect 6328 424056 6334 424108
rect 579798 422288 579804 422340
rect 579856 422328 579862 422340
rect 580902 422328 580908 422340
rect 579856 422300 580908 422328
rect 579856 422288 579862 422300
rect 580902 422288 580908 422300
rect 580960 422288 580966 422340
rect 470318 416712 470324 416764
rect 470376 416752 470382 416764
rect 579798 416752 579804 416764
rect 470376 416724 579804 416752
rect 470376 416712 470382 416724
rect 579798 416712 579804 416724
rect 579856 416712 579862 416764
rect 579798 412564 579804 412616
rect 579856 412604 579862 412616
rect 580902 412604 580908 412616
rect 579856 412576 580908 412604
rect 579856 412564 579862 412576
rect 580902 412564 580908 412576
rect 580960 412564 580966 412616
rect 579798 402976 579804 403028
rect 579856 403016 579862 403028
rect 580902 403016 580908 403028
rect 579856 402988 580908 403016
rect 579856 402976 579862 402988
rect 580902 402976 580908 402988
rect 580960 402976 580966 403028
rect 470226 393252 470232 393304
rect 470284 393292 470290 393304
rect 579890 393292 579896 393304
rect 470284 393264 579896 393292
rect 470284 393252 470290 393264
rect 579890 393252 579896 393264
rect 579948 393252 579954 393304
rect 580902 393292 580908 393304
rect 580000 393264 580908 393292
rect 579798 393184 579804 393236
rect 579856 393224 579862 393236
rect 580000 393224 580028 393264
rect 580902 393252 580908 393264
rect 580960 393252 580966 393304
rect 579856 393196 580028 393224
rect 579856 393184 579862 393196
rect 579798 384276 579804 384328
rect 579856 384316 579862 384328
rect 580902 384316 580908 384328
rect 579856 384288 580908 384316
rect 579856 384276 579862 384288
rect 580902 384276 580908 384288
rect 580960 384276 580966 384328
rect 3234 380808 3240 380860
rect 3292 380848 3298 380860
rect 13078 380848 13084 380860
rect 3292 380820 13084 380848
rect 3292 380808 3298 380820
rect 13078 380808 13084 380820
rect 13136 380808 13142 380860
rect 579982 361224 579988 361276
rect 580040 361264 580046 361276
rect 580902 361264 580908 361276
rect 580040 361236 580908 361264
rect 580040 361224 580046 361236
rect 580902 361224 580908 361236
rect 580960 361224 580966 361276
rect 579798 360136 579804 360188
rect 579856 360176 579862 360188
rect 579982 360176 579988 360188
rect 579856 360148 579988 360176
rect 579856 360136 579862 360148
rect 579982 360136 579988 360148
rect 580040 360136 580046 360188
rect 470134 346332 470140 346384
rect 470192 346372 470198 346384
rect 579798 346372 579804 346384
rect 470192 346344 579804 346372
rect 470192 346332 470198 346344
rect 579798 346332 579804 346344
rect 579856 346332 579862 346384
rect 580074 345040 580080 345092
rect 580132 345080 580138 345092
rect 580902 345080 580908 345092
rect 580132 345052 580908 345080
rect 580132 345040 580138 345052
rect 580902 345040 580908 345052
rect 580960 345040 580966 345092
rect 580074 344904 580080 344956
rect 580132 344944 580138 344956
rect 580902 344944 580908 344956
rect 580132 344916 580908 344944
rect 580132 344904 580138 344916
rect 580902 344904 580908 344916
rect 580960 344904 580966 344956
rect 460569 338147 460627 338153
rect 460569 338113 460581 338147
rect 460615 338144 460627 338147
rect 466365 338147 466423 338153
rect 466365 338144 466377 338147
rect 460615 338116 466377 338144
rect 460615 338113 460627 338116
rect 460569 338107 460627 338113
rect 466365 338113 466377 338116
rect 466411 338113 466423 338147
rect 466365 338107 466423 338113
rect 71038 338036 71044 338088
rect 71096 338076 71102 338088
rect 254946 338076 254952 338088
rect 71096 338048 254952 338076
rect 71096 338036 71102 338048
rect 254946 338036 254952 338048
rect 255004 338036 255010 338088
rect 284386 338076 284392 338088
rect 284347 338048 284392 338076
rect 284386 338036 284392 338048
rect 284444 338036 284450 338088
rect 316681 338079 316739 338085
rect 316681 338045 316693 338079
rect 316727 338076 316739 338079
rect 354398 338076 354404 338088
rect 316727 338048 354404 338076
rect 316727 338045 316739 338048
rect 316681 338039 316739 338045
rect 354398 338036 354404 338048
rect 354456 338036 354462 338088
rect 358078 338036 358084 338088
rect 358136 338076 358142 338088
rect 371510 338076 371516 338088
rect 358136 338048 371516 338076
rect 358136 338036 358142 338048
rect 371510 338036 371516 338048
rect 371568 338036 371574 338088
rect 376662 338036 376668 338088
rect 376720 338076 376726 338088
rect 379425 338079 379483 338085
rect 379425 338076 379437 338079
rect 376720 338048 379437 338076
rect 376720 338036 376726 338048
rect 379425 338045 379437 338048
rect 379471 338045 379483 338079
rect 379425 338039 379483 338045
rect 379517 338079 379575 338085
rect 379517 338045 379529 338079
rect 379563 338076 379575 338079
rect 380342 338076 380348 338088
rect 379563 338048 380348 338076
rect 379563 338045 379575 338048
rect 379517 338039 379575 338045
rect 380342 338036 380348 338048
rect 380400 338036 380406 338088
rect 406286 338036 406292 338088
rect 406344 338076 406350 338088
rect 417418 338076 417424 338088
rect 406344 338048 417424 338076
rect 406344 338036 406350 338048
rect 417418 338036 417424 338048
rect 417476 338036 417482 338088
rect 419074 338036 419080 338088
rect 419132 338076 419138 338088
rect 431402 338076 431408 338088
rect 419132 338048 431408 338076
rect 419132 338036 419138 338048
rect 431402 338036 431408 338048
rect 431460 338036 431466 338088
rect 435726 338036 435732 338088
rect 435784 338076 435790 338088
rect 499574 338076 499580 338088
rect 435784 338048 499580 338076
rect 435784 338036 435790 338048
rect 499574 338036 499580 338048
rect 499632 338036 499638 338088
rect 66898 337968 66904 338020
rect 66956 338008 66962 338020
rect 252002 338008 252008 338020
rect 66956 337980 252008 338008
rect 66956 337968 66962 337980
rect 252002 337968 252008 337980
rect 252060 337968 252066 338020
rect 306190 337968 306196 338020
rect 306248 338008 306254 338020
rect 355870 338008 355876 338020
rect 306248 337980 355876 338008
rect 306248 337968 306254 337980
rect 355870 337968 355876 337980
rect 355928 337968 355934 338020
rect 364242 337968 364248 338020
rect 364300 338008 364306 338020
rect 376754 338008 376760 338020
rect 364300 337980 376760 338008
rect 364300 337968 364306 337980
rect 376754 337968 376760 337980
rect 376812 337968 376818 338020
rect 382274 338008 382280 338020
rect 379440 337980 382280 338008
rect 61378 337900 61384 337952
rect 61436 337940 61442 337952
rect 247586 337940 247592 337952
rect 61436 337912 247592 337940
rect 61436 337900 61442 337912
rect 247586 337900 247592 337912
rect 247644 337900 247650 337952
rect 303154 337900 303160 337952
rect 303212 337940 303218 337952
rect 352926 337940 352932 337952
rect 303212 337912 352932 337940
rect 303212 337900 303218 337912
rect 352926 337900 352932 337912
rect 352984 337900 352990 337952
rect 355318 337900 355324 337952
rect 355376 337940 355382 337952
rect 370038 337940 370044 337952
rect 355376 337912 370044 337940
rect 355376 337900 355382 337912
rect 370038 337900 370044 337912
rect 370096 337900 370102 337952
rect 371142 337900 371148 337952
rect 371200 337940 371206 337952
rect 379440 337940 379468 337980
rect 382274 337968 382280 337980
rect 382332 337968 382338 338020
rect 404354 337968 404360 338020
rect 404412 338008 404418 338020
rect 412545 338011 412603 338017
rect 412545 338008 412557 338011
rect 404412 337980 412557 338008
rect 404412 337968 404418 337980
rect 412545 337977 412557 337980
rect 412591 337977 412603 338011
rect 412545 337971 412603 337977
rect 414658 337968 414664 338020
rect 414716 338008 414722 338020
rect 429746 338008 429752 338020
rect 414716 337980 429752 338008
rect 414716 337968 414722 337980
rect 429746 337968 429752 337980
rect 429804 337968 429810 338020
rect 437198 337968 437204 338020
rect 437256 338008 437262 338020
rect 442350 338008 442356 338020
rect 437256 337980 442356 338008
rect 437256 337968 437262 337980
rect 442350 337968 442356 337980
rect 442408 337968 442414 338020
rect 446030 337968 446036 338020
rect 446088 338008 446094 338020
rect 451185 338011 451243 338017
rect 451185 338008 451197 338011
rect 446088 337980 451197 338008
rect 446088 337968 446094 337980
rect 451185 337977 451197 337980
rect 451231 337977 451243 338011
rect 451185 337971 451243 337977
rect 451826 337968 451832 338020
rect 451884 338008 451890 338020
rect 461581 338011 461639 338017
rect 461581 338008 461593 338011
rect 451884 337980 461593 338008
rect 451884 337968 451890 337980
rect 461581 337977 461593 337980
rect 461627 337977 461639 338011
rect 461581 337971 461639 337977
rect 461670 337968 461676 338020
rect 461728 338008 461734 338020
rect 466273 338011 466331 338017
rect 466273 338008 466285 338011
rect 461728 337980 466285 338008
rect 461728 337968 461734 337980
rect 466273 337977 466285 337980
rect 466319 337977 466331 338011
rect 525058 338008 525064 338020
rect 466273 337971 466331 337977
rect 466380 337980 525064 338008
rect 371200 337912 379468 337940
rect 371200 337900 371206 337912
rect 400398 337900 400404 337952
rect 400456 337940 400462 337952
rect 413278 337940 413284 337952
rect 400456 337912 413284 337940
rect 400456 337900 400462 337912
rect 413278 337900 413284 337912
rect 413336 337900 413342 337952
rect 413646 337900 413652 337952
rect 413704 337940 413710 337952
rect 420178 337940 420184 337952
rect 413704 337912 420184 337940
rect 413704 337900 413710 337912
rect 420178 337900 420184 337912
rect 420236 337900 420242 337952
rect 420546 337900 420552 337952
rect 420604 337940 420610 337952
rect 454681 337943 454739 337949
rect 454681 337940 454693 337943
rect 420604 337912 454693 337940
rect 420604 337900 420610 337912
rect 454681 337909 454693 337912
rect 454727 337909 454739 337943
rect 454681 337903 454739 337909
rect 454770 337900 454776 337952
rect 454828 337940 454834 337952
rect 460569 337943 460627 337949
rect 460569 337940 460581 337943
rect 454828 337912 460581 337940
rect 454828 337900 454834 337912
rect 460569 337909 460581 337912
rect 460615 337909 460627 337943
rect 460569 337903 460627 337909
rect 460658 337900 460664 337952
rect 460716 337940 460722 337952
rect 466380 337940 466408 337980
rect 525058 337968 525064 337980
rect 525116 337968 525122 338020
rect 460716 337912 466408 337940
rect 460716 337900 460722 337912
rect 467098 337900 467104 337952
rect 467156 337940 467162 337952
rect 467742 337940 467748 337952
rect 467156 337912 467748 337940
rect 467156 337900 467162 337912
rect 467742 337900 467748 337912
rect 467800 337900 467806 337952
rect 468018 337900 468024 337952
rect 468076 337940 468082 337952
rect 469122 337940 469128 337952
rect 468076 337912 469128 337940
rect 468076 337900 468082 337912
rect 469122 337900 469128 337912
rect 469180 337900 469186 337952
rect 469217 337943 469275 337949
rect 469217 337909 469229 337943
rect 469263 337940 469275 337943
rect 527818 337940 527824 337952
rect 469263 337912 527824 337940
rect 469263 337909 469275 337912
rect 469217 337903 469275 337909
rect 527818 337900 527824 337912
rect 527876 337900 527882 337952
rect 57238 337832 57244 337884
rect 57296 337872 57302 337884
rect 247126 337872 247132 337884
rect 57296 337844 247132 337872
rect 57296 337832 57302 337844
rect 247126 337832 247132 337844
rect 247184 337832 247190 337884
rect 290458 337832 290464 337884
rect 290516 337872 290522 337884
rect 335909 337875 335967 337881
rect 335909 337872 335921 337875
rect 290516 337844 335921 337872
rect 290516 337832 290522 337844
rect 335909 337841 335921 337844
rect 335955 337841 335967 337875
rect 335909 337835 335967 337841
rect 336001 337875 336059 337881
rect 336001 337841 336013 337875
rect 336047 337872 336059 337875
rect 347038 337872 347044 337884
rect 336047 337844 347044 337872
rect 336047 337841 336059 337844
rect 336001 337835 336059 337841
rect 347038 337832 347044 337844
rect 347096 337832 347102 337884
rect 348418 337832 348424 337884
rect 348476 337872 348482 337884
rect 365622 337872 365628 337884
rect 348476 337844 365628 337872
rect 348476 337832 348482 337844
rect 365622 337832 365628 337844
rect 365680 337832 365686 337884
rect 365717 337875 365775 337881
rect 365717 337841 365729 337875
rect 365763 337872 365775 337875
rect 377398 337872 377404 337884
rect 365763 337844 377404 337872
rect 365763 337841 365775 337844
rect 365717 337835 365775 337841
rect 377398 337832 377404 337844
rect 377456 337832 377462 337884
rect 398466 337832 398472 337884
rect 398524 337872 398530 337884
rect 408770 337872 408776 337884
rect 398524 337844 408776 337872
rect 398524 337832 398530 337844
rect 408770 337832 408776 337844
rect 408828 337832 408834 337884
rect 414198 337832 414204 337884
rect 414256 337872 414262 337884
rect 415302 337872 415308 337884
rect 414256 337844 415308 337872
rect 414256 337832 414262 337844
rect 415302 337832 415308 337844
rect 415360 337832 415366 337884
rect 416056 337844 416820 337872
rect 50338 337764 50344 337816
rect 50396 337804 50402 337816
rect 244182 337804 244188 337816
rect 50396 337776 244188 337804
rect 50396 337764 50402 337776
rect 244182 337764 244188 337776
rect 244240 337764 244246 337816
rect 259638 337764 259644 337816
rect 259696 337804 259702 337816
rect 260098 337804 260104 337816
rect 259696 337776 260104 337804
rect 259696 337764 259702 337776
rect 260098 337764 260104 337776
rect 260156 337764 260162 337816
rect 288250 337764 288256 337816
rect 288308 337804 288314 337816
rect 302237 337807 302295 337813
rect 288308 337776 297404 337804
rect 288308 337764 288314 337776
rect 32398 337696 32404 337748
rect 32456 337736 32462 337748
rect 237834 337736 237840 337748
rect 32456 337708 237840 337736
rect 32456 337696 32462 337708
rect 237834 337696 237840 337708
rect 237892 337696 237898 337748
rect 248506 337696 248512 337748
rect 248564 337736 248570 337748
rect 249518 337736 249524 337748
rect 248564 337708 249524 337736
rect 248564 337696 248570 337708
rect 249518 337696 249524 337708
rect 249576 337696 249582 337748
rect 251450 337696 251456 337748
rect 251508 337736 251514 337748
rect 252462 337736 252468 337748
rect 251508 337708 252468 337736
rect 251508 337696 251514 337708
rect 252462 337696 252468 337708
rect 252520 337696 252526 337748
rect 254578 337696 254584 337748
rect 254636 337736 254642 337748
rect 262306 337736 262312 337748
rect 254636 337708 262312 337736
rect 254636 337696 254642 337708
rect 262306 337696 262312 337708
rect 262364 337696 262370 337748
rect 297376 337736 297404 337776
rect 302237 337773 302249 337807
rect 302283 337804 302295 337807
rect 351914 337804 351920 337816
rect 302283 337776 351920 337804
rect 302283 337773 302295 337776
rect 302237 337767 302295 337773
rect 351914 337764 351920 337776
rect 351972 337764 351978 337816
rect 358722 337764 358728 337816
rect 358780 337804 358786 337816
rect 358780 337776 362816 337804
rect 358780 337764 358786 337776
rect 348510 337736 348516 337748
rect 297376 337708 348516 337736
rect 348510 337696 348516 337708
rect 348568 337696 348574 337748
rect 348973 337739 349031 337745
rect 348973 337705 348985 337739
rect 349019 337736 349031 337739
rect 360105 337739 360163 337745
rect 360105 337736 360117 337739
rect 349019 337708 360117 337736
rect 349019 337705 349031 337708
rect 348973 337699 349031 337705
rect 360105 337705 360117 337708
rect 360151 337705 360163 337739
rect 360105 337699 360163 337705
rect 39298 337628 39304 337680
rect 39356 337668 39362 337680
rect 244642 337668 244648 337680
rect 39356 337640 244648 337668
rect 39356 337628 39362 337640
rect 244642 337628 244648 337640
rect 244700 337628 244706 337680
rect 260098 337628 260104 337680
rect 260156 337668 260162 337680
rect 277026 337668 277032 337680
rect 260156 337640 277032 337668
rect 260156 337628 260162 337640
rect 277026 337628 277032 337640
rect 277084 337628 277090 337680
rect 285582 337628 285588 337680
rect 285640 337668 285646 337680
rect 336001 337671 336059 337677
rect 336001 337668 336013 337671
rect 285640 337640 336013 337668
rect 285640 337628 285646 337640
rect 336001 337637 336013 337640
rect 336047 337637 336059 337671
rect 336001 337631 336059 337637
rect 336090 337628 336096 337680
rect 336148 337668 336154 337680
rect 344554 337668 344560 337680
rect 336148 337640 344560 337668
rect 336148 337628 336154 337640
rect 344554 337628 344560 337640
rect 344612 337628 344618 337680
rect 344649 337671 344707 337677
rect 344649 337637 344661 337671
rect 344695 337668 344707 337671
rect 349982 337668 349988 337680
rect 344695 337640 349988 337668
rect 344695 337637 344707 337640
rect 344649 337631 344707 337637
rect 349982 337628 349988 337640
rect 350040 337628 350046 337680
rect 354858 337668 354864 337680
rect 350276 337640 354864 337668
rect 35158 337560 35164 337612
rect 35216 337600 35222 337612
rect 241698 337600 241704 337612
rect 35216 337572 241704 337600
rect 35216 337560 35222 337572
rect 241698 337560 241704 337572
rect 241756 337560 241762 337612
rect 255958 337560 255964 337612
rect 256016 337600 256022 337612
rect 260469 337603 260527 337609
rect 260469 337600 260481 337603
rect 256016 337572 260481 337600
rect 256016 337560 256022 337572
rect 260469 337569 260481 337572
rect 260515 337569 260527 337603
rect 260469 337563 260527 337569
rect 261386 337560 261392 337612
rect 261444 337600 261450 337612
rect 279970 337600 279976 337612
rect 261444 337572 279976 337600
rect 261444 337560 261450 337572
rect 279970 337560 279976 337572
rect 280028 337560 280034 337612
rect 281442 337560 281448 337612
rect 281500 337600 281506 337612
rect 345566 337600 345572 337612
rect 281500 337572 345572 337600
rect 281500 337560 281506 337572
rect 345566 337560 345572 337572
rect 345624 337560 345630 337612
rect 345661 337603 345719 337609
rect 345661 337569 345673 337603
rect 345707 337600 345719 337603
rect 350166 337600 350172 337612
rect 345707 337572 350172 337600
rect 345707 337569 345719 337572
rect 345661 337563 345719 337569
rect 350166 337560 350172 337572
rect 350224 337560 350230 337612
rect 28258 337492 28264 337544
rect 28316 337532 28322 337544
rect 28316 337504 234476 337532
rect 28316 337492 28322 337504
rect 19978 337424 19984 337476
rect 20036 337464 20042 337476
rect 234338 337464 234344 337476
rect 20036 337436 234344 337464
rect 20036 337424 20042 337436
rect 234338 337424 234344 337436
rect 234396 337424 234402 337476
rect 234448 337464 234476 337504
rect 253198 337492 253204 337544
rect 253256 337532 253262 337544
rect 259362 337532 259368 337544
rect 253256 337504 259368 337532
rect 253256 337492 253262 337504
rect 259362 337492 259368 337504
rect 259420 337492 259426 337544
rect 275554 337532 275560 337544
rect 260300 337504 275560 337532
rect 238294 337464 238300 337476
rect 234448 337436 238300 337464
rect 238294 337424 238300 337436
rect 238352 337424 238358 337476
rect 258718 337424 258724 337476
rect 258776 337464 258782 337476
rect 260300 337464 260328 337504
rect 275554 337492 275560 337504
rect 275612 337492 275618 337544
rect 275922 337492 275928 337544
rect 275980 337532 275986 337544
rect 335817 337535 335875 337541
rect 335817 337532 335829 337535
rect 275980 337504 335829 337532
rect 275980 337492 275986 337504
rect 335817 337501 335829 337504
rect 335863 337501 335875 337535
rect 341610 337532 341616 337544
rect 335817 337495 335875 337501
rect 336016 337504 341616 337532
rect 269666 337464 269672 337476
rect 258776 337436 260328 337464
rect 260392 337436 269672 337464
rect 258776 337424 258782 337436
rect 13078 337356 13084 337408
rect 13136 337396 13142 337408
rect 233510 337396 233516 337408
rect 13136 337368 233516 337396
rect 13136 337356 13142 337368
rect 233510 337356 233516 337368
rect 233568 337356 233574 337408
rect 233878 337356 233884 337408
rect 233936 337396 233942 337408
rect 241238 337396 241244 337408
rect 233936 337368 241244 337396
rect 233936 337356 233942 337368
rect 241238 337356 241244 337368
rect 241296 337356 241302 337408
rect 250438 337356 250444 337408
rect 250496 337396 250502 337408
rect 253474 337396 253480 337408
rect 250496 337368 253480 337396
rect 250496 337356 250502 337368
rect 253474 337356 253480 337368
rect 253532 337356 253538 337408
rect 257338 337356 257344 337408
rect 257396 337396 257402 337408
rect 260392 337396 260420 337436
rect 269666 337424 269672 337436
rect 269724 337424 269730 337476
rect 271782 337424 271788 337476
rect 271840 337464 271846 337476
rect 336016 337464 336044 337504
rect 341610 337492 341616 337504
rect 341668 337492 341674 337544
rect 342809 337535 342867 337541
rect 342809 337501 342821 337535
rect 342855 337532 342867 337535
rect 344281 337535 344339 337541
rect 344281 337532 344293 337535
rect 342855 337504 344293 337532
rect 342855 337501 342867 337504
rect 342809 337495 342867 337501
rect 344281 337501 344293 337504
rect 344327 337501 344339 337535
rect 344281 337495 344339 337501
rect 344370 337492 344376 337544
rect 344428 337532 344434 337544
rect 350276 337532 350304 337640
rect 354858 337628 354864 337640
rect 354916 337628 354922 337680
rect 356698 337628 356704 337680
rect 356756 337668 356762 337680
rect 360746 337668 360752 337680
rect 356756 337640 360752 337668
rect 356756 337628 356762 337640
rect 360746 337628 360752 337640
rect 360804 337628 360810 337680
rect 362788 337668 362816 337776
rect 362862 337764 362868 337816
rect 362920 337804 362926 337816
rect 378870 337804 378876 337816
rect 362920 337776 378876 337804
rect 362920 337764 362926 337776
rect 378870 337764 378876 337776
rect 378928 337764 378934 337816
rect 388438 337764 388444 337816
rect 388496 337804 388502 337816
rect 389174 337804 389180 337816
rect 388496 337776 389180 337804
rect 388496 337764 388502 337776
rect 389174 337764 389180 337776
rect 389232 337764 389238 337816
rect 407298 337764 407304 337816
rect 407356 337804 407362 337816
rect 412453 337807 412511 337813
rect 412453 337804 412465 337807
rect 407356 337776 412465 337804
rect 407356 337764 407362 337776
rect 412453 337773 412465 337776
rect 412499 337773 412511 337807
rect 412453 337767 412511 337773
rect 412545 337807 412603 337813
rect 412545 337773 412557 337807
rect 412591 337804 412603 337807
rect 416056 337804 416084 337844
rect 412591 337776 416084 337804
rect 412591 337773 412603 337776
rect 412545 337767 412603 337773
rect 416130 337764 416136 337816
rect 416188 337804 416194 337816
rect 416682 337804 416688 337816
rect 416188 337776 416688 337804
rect 416188 337764 416194 337776
rect 416682 337764 416688 337776
rect 416740 337764 416746 337816
rect 416792 337804 416820 337844
rect 417602 337832 417608 337884
rect 417660 337872 417666 337884
rect 455598 337872 455604 337884
rect 417660 337844 455604 337872
rect 417660 337832 417666 337844
rect 455598 337832 455604 337844
rect 455656 337832 455662 337884
rect 457714 337832 457720 337884
rect 457772 337872 457778 337884
rect 523678 337872 523684 337884
rect 457772 337844 523684 337872
rect 457772 337832 457778 337844
rect 523678 337832 523684 337844
rect 523736 337832 523742 337884
rect 420270 337804 420276 337816
rect 416792 337776 420276 337804
rect 420270 337764 420276 337776
rect 420328 337764 420334 337816
rect 422018 337764 422024 337816
rect 422076 337804 422082 337816
rect 438118 337804 438124 337816
rect 422076 337776 438124 337804
rect 422076 337764 422082 337776
rect 438118 337764 438124 337776
rect 438176 337764 438182 337816
rect 438670 337764 438676 337816
rect 438728 337804 438734 337816
rect 438728 337776 440280 337804
rect 438728 337764 438734 337776
rect 364337 337739 364395 337745
rect 364337 337705 364349 337739
rect 364383 337736 364395 337739
rect 369578 337736 369584 337748
rect 364383 337708 369584 337736
rect 364383 337705 364395 337708
rect 364337 337699 364395 337705
rect 369578 337696 369584 337708
rect 369636 337696 369642 337748
rect 375926 337736 375932 337748
rect 372908 337708 375932 337736
rect 364981 337671 365039 337677
rect 362788 337640 364748 337668
rect 351178 337560 351184 337612
rect 351236 337600 351242 337612
rect 364720 337600 364748 337640
rect 364981 337637 364993 337671
rect 365027 337668 365039 337671
rect 372908 337668 372936 337708
rect 375926 337696 375932 337708
rect 375984 337696 375990 337748
rect 380158 337696 380164 337748
rect 380216 337736 380222 337748
rect 381354 337736 381360 337748
rect 380216 337708 381360 337736
rect 380216 337696 380222 337708
rect 381354 337696 381360 337708
rect 381412 337696 381418 337748
rect 381538 337696 381544 337748
rect 381596 337736 381602 337748
rect 382826 337736 382832 337748
rect 381596 337708 382832 337736
rect 381596 337696 381602 337708
rect 382826 337696 382832 337708
rect 382884 337696 382890 337748
rect 384942 337696 384948 337748
rect 385000 337736 385006 337748
rect 388162 337736 388168 337748
rect 385000 337708 388168 337736
rect 385000 337696 385006 337708
rect 388162 337696 388168 337708
rect 388220 337696 388226 337748
rect 398926 337696 398932 337748
rect 398984 337736 398990 337748
rect 398984 337708 400996 337736
rect 398984 337696 398990 337708
rect 376570 337668 376576 337680
rect 365027 337640 372936 337668
rect 373092 337640 376576 337668
rect 365027 337637 365039 337640
rect 364981 337631 365039 337637
rect 365717 337603 365775 337609
rect 365717 337600 365729 337603
rect 351236 337572 364656 337600
rect 364720 337572 365729 337600
rect 351236 337560 351242 337572
rect 344428 337504 350304 337532
rect 344428 337492 344434 337504
rect 351822 337492 351828 337544
rect 351880 337532 351886 337544
rect 364429 337535 364487 337541
rect 364429 337532 364441 337535
rect 351880 337504 364441 337532
rect 351880 337492 351886 337504
rect 364429 337501 364441 337504
rect 364475 337501 364487 337535
rect 364429 337495 364487 337501
rect 271840 337436 336044 337464
rect 336093 337467 336151 337473
rect 271840 337424 271846 337436
rect 336093 337433 336105 337467
rect 336139 337464 336151 337467
rect 344094 337464 344100 337476
rect 336139 337436 344100 337464
rect 336139 337433 336151 337436
rect 336093 337427 336151 337433
rect 344094 337424 344100 337436
rect 344152 337424 344158 337476
rect 347777 337467 347835 337473
rect 347777 337433 347789 337467
rect 347823 337464 347835 337467
rect 348973 337467 349031 337473
rect 348973 337464 348985 337467
rect 347823 337436 348985 337464
rect 347823 337433 347835 337436
rect 347777 337427 347835 337433
rect 348973 337433 348985 337436
rect 349019 337433 349031 337467
rect 348973 337427 349031 337433
rect 349062 337424 349068 337476
rect 349120 337464 349126 337476
rect 364628 337464 364656 337572
rect 365717 337569 365729 337572
rect 365763 337569 365775 337603
rect 365717 337563 365775 337569
rect 366910 337560 366916 337612
rect 366968 337600 366974 337612
rect 373092 337600 373120 337640
rect 376570 337628 376576 337640
rect 376628 337628 376634 337680
rect 384298 337628 384304 337680
rect 384356 337668 384362 337680
rect 387702 337668 387708 337680
rect 384356 337640 387708 337668
rect 384356 337628 384362 337640
rect 387702 337628 387708 337640
rect 387760 337628 387766 337680
rect 398006 337628 398012 337680
rect 398064 337668 398070 337680
rect 399478 337668 399484 337680
rect 398064 337640 399484 337668
rect 398064 337628 398070 337640
rect 399478 337628 399484 337640
rect 399536 337628 399542 337680
rect 400968 337668 400996 337708
rect 403342 337696 403348 337748
rect 403400 337736 403406 337748
rect 403400 337708 410196 337736
rect 403400 337696 403406 337708
rect 406378 337668 406384 337680
rect 400968 337640 406384 337668
rect 406378 337628 406384 337640
rect 406436 337628 406442 337680
rect 410168 337668 410196 337708
rect 410242 337696 410248 337748
rect 410300 337736 410306 337748
rect 411070 337736 411076 337748
rect 410300 337708 411076 337736
rect 410300 337696 410306 337708
rect 411070 337696 411076 337708
rect 411128 337696 411134 337748
rect 411180 337708 414244 337736
rect 411180 337668 411208 337708
rect 410168 337640 411208 337668
rect 411254 337628 411260 337680
rect 411312 337668 411318 337680
rect 412358 337668 412364 337680
rect 411312 337640 412364 337668
rect 411312 337628 411318 337640
rect 412358 337628 412364 337640
rect 412416 337628 412422 337680
rect 412453 337671 412511 337677
rect 412453 337637 412465 337671
rect 412499 337668 412511 337671
rect 413925 337671 413983 337677
rect 413925 337668 413937 337671
rect 412499 337640 413937 337668
rect 412499 337637 412511 337640
rect 412453 337631 412511 337637
rect 413925 337637 413937 337640
rect 413971 337637 413983 337671
rect 413925 337631 413983 337637
rect 383286 337600 383292 337612
rect 366968 337572 373120 337600
rect 374748 337572 383292 337600
rect 366968 337560 366974 337572
rect 364705 337535 364763 337541
rect 364705 337501 364717 337535
rect 364751 337532 364763 337535
rect 364751 337504 372200 337532
rect 364751 337501 364763 337504
rect 364705 337495 364763 337501
rect 372062 337464 372068 337476
rect 349120 337436 364564 337464
rect 364628 337436 372068 337464
rect 349120 337424 349126 337436
rect 257396 337368 260420 337396
rect 260469 337399 260527 337405
rect 257396 337356 257402 337368
rect 260469 337365 260481 337399
rect 260515 337396 260527 337399
rect 266722 337396 266728 337408
rect 260515 337368 266728 337396
rect 260515 337365 260527 337368
rect 260469 337359 260527 337365
rect 266722 337356 266728 337368
rect 266780 337356 266786 337408
rect 269022 337356 269028 337408
rect 269080 337396 269086 337408
rect 340230 337396 340236 337408
rect 269080 337368 340236 337396
rect 269080 337356 269086 337368
rect 340230 337356 340236 337368
rect 340288 337356 340294 337408
rect 340782 337356 340788 337408
rect 340840 337396 340846 337408
rect 364337 337399 364395 337405
rect 364337 337396 364349 337399
rect 340840 337368 364349 337396
rect 340840 337356 340846 337368
rect 364337 337365 364349 337368
rect 364383 337365 364395 337399
rect 364337 337359 364395 337365
rect 79318 337288 79324 337340
rect 79376 337328 79382 337340
rect 260834 337328 260840 337340
rect 79376 337300 260840 337328
rect 79376 337288 79382 337300
rect 260834 337288 260840 337300
rect 260892 337288 260898 337340
rect 271322 337288 271328 337340
rect 271380 337328 271386 337340
rect 271380 337300 303660 337328
rect 271380 337288 271386 337300
rect 103425 337263 103483 337269
rect 103425 337229 103437 337263
rect 103471 337260 103483 337263
rect 113177 337263 113235 337269
rect 113177 337260 113189 337263
rect 103471 337232 113189 337260
rect 103471 337229 103483 337232
rect 103425 337223 103483 337229
rect 113177 337229 113189 337232
rect 113223 337229 113235 337263
rect 113177 337223 113235 337229
rect 122745 337263 122803 337269
rect 122745 337229 122757 337263
rect 122791 337260 122803 337263
rect 132494 337260 132500 337272
rect 122791 337232 132500 337260
rect 122791 337229 122803 337232
rect 122745 337223 122803 337229
rect 132494 337220 132500 337232
rect 132552 337220 132558 337272
rect 142062 337220 142068 337272
rect 142120 337260 142126 337272
rect 151814 337260 151820 337272
rect 142120 337232 151820 337260
rect 142120 337220 142126 337232
rect 151814 337220 151820 337232
rect 151872 337220 151878 337272
rect 161382 337220 161388 337272
rect 161440 337260 161446 337272
rect 171134 337260 171140 337272
rect 161440 337232 171140 337260
rect 161440 337220 161446 337232
rect 171134 337220 171140 337232
rect 171192 337220 171198 337272
rect 180702 337220 180708 337272
rect 180760 337260 180766 337272
rect 190454 337260 190460 337272
rect 180760 337232 190460 337260
rect 180760 337220 180766 337232
rect 190454 337220 190460 337232
rect 190512 337220 190518 337272
rect 200022 337220 200028 337272
rect 200080 337260 200086 337272
rect 209774 337260 209780 337272
rect 200080 337232 209780 337260
rect 200080 337220 200086 337232
rect 209774 337220 209780 337232
rect 209832 337220 209838 337272
rect 219342 337220 219348 337272
rect 219400 337260 219406 337272
rect 229186 337260 229192 337272
rect 219400 337232 229192 337260
rect 219400 337220 219406 337232
rect 229186 337220 229192 337232
rect 229244 337220 229250 337272
rect 234614 337220 234620 337272
rect 234672 337260 234678 337272
rect 257890 337260 257896 337272
rect 234672 337232 257896 337260
rect 234672 337220 234678 337232
rect 257890 337220 257896 337232
rect 257948 337220 257954 337272
rect 258810 337220 258816 337272
rect 258868 337260 258874 337272
rect 272610 337260 272616 337272
rect 258868 337232 272616 337260
rect 258868 337220 258874 337232
rect 272610 337220 272616 337232
rect 272668 337220 272674 337272
rect 272794 337220 272800 337272
rect 272852 337260 272858 337272
rect 303632 337260 303660 337300
rect 309778 337288 309784 337340
rect 309836 337328 309842 337340
rect 316681 337331 316739 337337
rect 316681 337328 316693 337331
rect 309836 337300 316693 337328
rect 309836 337288 309842 337300
rect 316681 337297 316693 337300
rect 316727 337297 316739 337331
rect 347777 337331 347835 337337
rect 347777 337328 347789 337331
rect 316681 337291 316739 337297
rect 333164 337300 347789 337328
rect 312722 337260 312728 337272
rect 272852 337232 302372 337260
rect 303632 337232 312728 337260
rect 272852 337220 272858 337232
rect 84838 337152 84844 337204
rect 84896 337192 84902 337204
rect 263778 337192 263784 337204
rect 84896 337164 263784 337192
rect 84896 337152 84902 337164
rect 263778 337152 263784 337164
rect 263836 337152 263842 337204
rect 297910 337152 297916 337204
rect 297968 337192 297974 337204
rect 302237 337195 302295 337201
rect 302237 337192 302249 337195
rect 297968 337164 302249 337192
rect 297968 337152 297974 337164
rect 302237 337161 302249 337164
rect 302283 337161 302295 337195
rect 302237 337155 302295 337161
rect 86957 337127 87015 337133
rect 86957 337093 86969 337127
rect 87003 337124 87015 337127
rect 87003 337096 93900 337124
rect 87003 337093 87015 337096
rect 86957 337087 87015 337093
rect 77938 336948 77944 337000
rect 77996 336988 78002 337000
rect 86957 336991 87015 336997
rect 86957 336988 86969 336991
rect 77996 336960 86969 336988
rect 77996 336948 78002 336960
rect 86957 336957 86969 336960
rect 87003 336957 87015 336991
rect 93872 336988 93900 337096
rect 100662 337084 100668 337136
rect 100720 337124 100726 337136
rect 271138 337124 271144 337136
rect 100720 337096 271144 337124
rect 100720 337084 100726 337096
rect 271138 337084 271144 337096
rect 271196 337084 271202 337136
rect 302344 337124 302372 337232
rect 312722 337220 312728 337232
rect 312780 337220 312786 337272
rect 321833 337263 321891 337269
rect 321833 337229 321845 337263
rect 321879 337260 321891 337263
rect 333164 337260 333192 337300
rect 347777 337297 347789 337300
rect 347823 337297 347835 337331
rect 347777 337291 347835 337297
rect 360105 337331 360163 337337
rect 360105 337297 360117 337331
rect 360151 337328 360163 337331
rect 361758 337328 361764 337340
rect 360151 337300 361764 337328
rect 360151 337297 360163 337300
rect 360105 337291 360163 337297
rect 361758 337288 361764 337300
rect 361816 337288 361822 337340
rect 364536 337328 364564 337436
rect 372062 337424 372068 337436
rect 372120 337424 372126 337476
rect 372172 337464 372200 337504
rect 373902 337492 373908 337544
rect 373960 337532 373966 337544
rect 374748 337532 374776 337572
rect 383286 337560 383292 337572
rect 383344 337560 383350 337612
rect 404814 337560 404820 337612
rect 404872 337600 404878 337612
rect 412637 337603 412695 337609
rect 412637 337600 412649 337603
rect 404872 337572 412649 337600
rect 404872 337560 404878 337572
rect 412637 337569 412649 337572
rect 412683 337569 412695 337603
rect 412637 337563 412695 337569
rect 412726 337560 412732 337612
rect 412784 337600 412790 337612
rect 413830 337600 413836 337612
rect 412784 337572 413836 337600
rect 412784 337560 412790 337572
rect 413830 337560 413836 337572
rect 413888 337560 413894 337612
rect 414216 337600 414244 337708
rect 415578 337696 415584 337748
rect 415636 337736 415642 337748
rect 416498 337736 416504 337748
rect 415636 337708 416504 337736
rect 415636 337696 415642 337708
rect 416498 337696 416504 337708
rect 416556 337696 416562 337748
rect 417050 337696 417056 337748
rect 417108 337736 417114 337748
rect 417970 337736 417976 337748
rect 417108 337708 417976 337736
rect 417108 337696 417114 337708
rect 417970 337696 417976 337708
rect 418028 337696 418034 337748
rect 418522 337696 418528 337748
rect 418580 337736 418586 337748
rect 419442 337736 419448 337748
rect 418580 337708 419448 337736
rect 418580 337696 418586 337708
rect 419442 337696 419448 337708
rect 419500 337696 419506 337748
rect 419534 337696 419540 337748
rect 419592 337736 419598 337748
rect 420822 337736 420828 337748
rect 419592 337708 420828 337736
rect 419592 337696 419598 337708
rect 420822 337696 420828 337708
rect 420880 337696 420886 337748
rect 421466 337696 421472 337748
rect 421524 337736 421530 337748
rect 422202 337736 422208 337748
rect 421524 337708 422208 337736
rect 421524 337696 421530 337708
rect 422202 337696 422208 337708
rect 422260 337696 422266 337748
rect 422478 337696 422484 337748
rect 422536 337736 422542 337748
rect 424410 337736 424416 337748
rect 422536 337708 424416 337736
rect 422536 337696 422542 337708
rect 424410 337696 424416 337708
rect 424468 337696 424474 337748
rect 425422 337696 425428 337748
rect 425480 337736 425486 337748
rect 428458 337736 428464 337748
rect 425480 337708 428464 337736
rect 425480 337696 425486 337708
rect 428458 337696 428464 337708
rect 428516 337696 428522 337748
rect 429378 337696 429384 337748
rect 429436 337736 429442 337748
rect 430482 337736 430488 337748
rect 429436 337708 430488 337736
rect 429436 337696 429442 337708
rect 430482 337696 430488 337708
rect 430540 337696 430546 337748
rect 432233 337739 432291 337745
rect 432233 337736 432245 337739
rect 430592 337708 432245 337736
rect 414293 337671 414351 337677
rect 414293 337637 414305 337671
rect 414339 337668 414351 337671
rect 427078 337668 427084 337680
rect 414339 337640 427084 337668
rect 414339 337637 414351 337640
rect 414293 337631 414351 337637
rect 427078 337628 427084 337640
rect 427136 337628 427142 337680
rect 430592 337668 430620 337708
rect 432233 337705 432245 337708
rect 432279 337705 432291 337739
rect 432233 337699 432291 337705
rect 432322 337696 432328 337748
rect 432380 337736 432386 337748
rect 433150 337736 433156 337748
rect 432380 337708 433156 337736
rect 432380 337696 432386 337708
rect 433150 337696 433156 337708
rect 433208 337696 433214 337748
rect 433702 337696 433708 337748
rect 433760 337736 433766 337748
rect 434622 337736 434628 337748
rect 433760 337708 434628 337736
rect 433760 337696 433766 337708
rect 434622 337696 434628 337708
rect 434680 337696 434686 337748
rect 435174 337696 435180 337748
rect 435232 337736 435238 337748
rect 436002 337736 436008 337748
rect 435232 337708 436008 337736
rect 435232 337696 435238 337708
rect 436002 337696 436008 337708
rect 436060 337696 436066 337748
rect 436186 337696 436192 337748
rect 436244 337736 436250 337748
rect 437382 337736 437388 337748
rect 436244 337708 437388 337736
rect 436244 337696 436250 337708
rect 437382 337696 437388 337708
rect 437440 337696 437446 337748
rect 439130 337696 439136 337748
rect 439188 337736 439194 337748
rect 440142 337736 440148 337748
rect 439188 337708 440148 337736
rect 439188 337696 439194 337708
rect 440142 337696 440148 337708
rect 440200 337696 440206 337748
rect 440252 337736 440280 337776
rect 440602 337764 440608 337816
rect 440660 337804 440666 337816
rect 441522 337804 441528 337816
rect 440660 337776 441528 337804
rect 440660 337764 440666 337776
rect 441522 337764 441528 337776
rect 441580 337764 441586 337816
rect 442074 337764 442080 337816
rect 442132 337804 442138 337816
rect 442902 337804 442908 337816
rect 442132 337776 442908 337804
rect 442132 337764 442138 337776
rect 442902 337764 442908 337776
rect 442960 337764 442966 337816
rect 444558 337764 444564 337816
rect 444616 337804 444622 337816
rect 445662 337804 445668 337816
rect 444616 337776 445668 337804
rect 444616 337764 444622 337776
rect 445662 337764 445668 337776
rect 445720 337764 445726 337816
rect 448974 337764 448980 337816
rect 449032 337804 449038 337816
rect 451093 337807 451151 337813
rect 451093 337804 451105 337807
rect 449032 337776 451105 337804
rect 449032 337764 449038 337776
rect 451093 337773 451105 337776
rect 451139 337773 451151 337807
rect 451093 337767 451151 337773
rect 451185 337807 451243 337813
rect 451185 337773 451197 337807
rect 451231 337804 451243 337807
rect 451277 337807 451335 337813
rect 451277 337804 451289 337807
rect 451231 337776 451289 337804
rect 451231 337773 451243 337776
rect 451185 337767 451243 337773
rect 451277 337773 451289 337776
rect 451323 337773 451335 337807
rect 451277 337767 451335 337773
rect 451366 337764 451372 337816
rect 451424 337804 451430 337816
rect 452470 337804 452476 337816
rect 451424 337776 452476 337804
rect 451424 337764 451430 337776
rect 452470 337764 452476 337776
rect 452528 337764 452534 337816
rect 452838 337764 452844 337816
rect 452896 337804 452902 337816
rect 453758 337804 453764 337816
rect 452896 337776 453764 337804
rect 452896 337764 452902 337776
rect 453758 337764 453764 337776
rect 453816 337764 453822 337816
rect 454310 337764 454316 337816
rect 454368 337804 454374 337816
rect 455230 337804 455236 337816
rect 454368 337776 455236 337804
rect 454368 337764 454374 337776
rect 455230 337764 455236 337776
rect 455288 337764 455294 337816
rect 455782 337764 455788 337816
rect 455840 337804 455846 337816
rect 456610 337804 456616 337816
rect 455840 337776 456616 337804
rect 455840 337764 455846 337776
rect 456610 337764 456616 337776
rect 456668 337764 456674 337816
rect 460198 337764 460204 337816
rect 460256 337804 460262 337816
rect 460750 337804 460756 337816
rect 460256 337776 460756 337804
rect 460256 337764 460262 337776
rect 460750 337764 460756 337776
rect 460808 337764 460814 337816
rect 466365 337807 466423 337813
rect 466365 337773 466377 337807
rect 466411 337804 466423 337807
rect 520918 337804 520924 337816
rect 466411 337776 520924 337804
rect 466411 337773 466423 337776
rect 466365 337767 466423 337773
rect 520918 337764 520924 337776
rect 520976 337764 520982 337816
rect 506474 337736 506480 337748
rect 440252 337708 506480 337736
rect 506474 337696 506480 337708
rect 506532 337696 506538 337748
rect 428292 337640 430620 337668
rect 421190 337600 421196 337612
rect 414216 337572 421196 337600
rect 421190 337560 421196 337572
rect 421248 337560 421254 337612
rect 426802 337560 426808 337612
rect 426860 337600 426866 337612
rect 428292 337600 428320 337640
rect 430850 337628 430856 337680
rect 430908 337668 430914 337680
rect 431862 337668 431868 337680
rect 430908 337640 431868 337668
rect 430908 337628 430914 337640
rect 431862 337628 431868 337640
rect 431920 337628 431926 337680
rect 434714 337628 434720 337680
rect 434772 337668 434778 337680
rect 435910 337668 435916 337680
rect 434772 337640 435916 337668
rect 434772 337628 434778 337640
rect 435910 337628 435916 337640
rect 435968 337628 435974 337680
rect 436646 337628 436652 337680
rect 436704 337668 436710 337680
rect 437290 337668 437296 337680
rect 436704 337640 437296 337668
rect 436704 337628 436710 337640
rect 437290 337628 437296 337640
rect 437348 337628 437354 337680
rect 440234 337628 440240 337680
rect 440292 337668 440298 337680
rect 443457 337671 443515 337677
rect 443457 337668 443469 337671
rect 440292 337640 443469 337668
rect 440292 337628 440298 337640
rect 443457 337637 443469 337640
rect 443503 337637 443515 337671
rect 443457 337631 443515 337637
rect 443546 337628 443552 337680
rect 443604 337668 443610 337680
rect 444282 337668 444288 337680
rect 443604 337640 444288 337668
rect 443604 337628 443610 337640
rect 444282 337628 444288 337640
rect 444340 337628 444346 337680
rect 445018 337628 445024 337680
rect 445076 337668 445082 337680
rect 445570 337668 445576 337680
rect 445076 337640 445576 337668
rect 445076 337628 445082 337640
rect 445570 337628 445576 337640
rect 445628 337628 445634 337680
rect 446490 337628 446496 337680
rect 446548 337668 446554 337680
rect 447042 337668 447048 337680
rect 446548 337640 447048 337668
rect 446548 337628 446554 337640
rect 447042 337628 447048 337640
rect 447100 337628 447106 337680
rect 448238 337628 448244 337680
rect 448296 337668 448302 337680
rect 448422 337668 448428 337680
rect 448296 337640 448428 337668
rect 448296 337628 448302 337640
rect 448422 337628 448428 337640
rect 448480 337628 448486 337680
rect 449894 337628 449900 337680
rect 449952 337668 449958 337680
rect 450998 337668 451004 337680
rect 449952 337640 451004 337668
rect 449952 337628 449958 337640
rect 450998 337628 451004 337640
rect 451056 337628 451062 337680
rect 451093 337671 451151 337677
rect 451093 337637 451105 337671
rect 451139 337668 451151 337671
rect 518158 337668 518164 337680
rect 451139 337640 518164 337668
rect 451139 337637 451151 337640
rect 451093 337631 451151 337637
rect 518158 337628 518164 337640
rect 518216 337628 518222 337680
rect 426860 337572 428320 337600
rect 426860 337560 426866 337572
rect 428366 337560 428372 337612
rect 428424 337600 428430 337612
rect 431218 337600 431224 337612
rect 428424 337572 431224 337600
rect 428424 337560 428430 337572
rect 431218 337560 431224 337572
rect 431276 337560 431282 337612
rect 431310 337560 431316 337612
rect 431368 337600 431374 337612
rect 449158 337600 449164 337612
rect 431368 337572 449164 337600
rect 431368 337560 431374 337572
rect 449158 337560 449164 337572
rect 449216 337560 449222 337612
rect 450446 337560 450452 337612
rect 450504 337600 450510 337612
rect 451182 337600 451188 337612
rect 450504 337572 451188 337600
rect 450504 337560 450510 337572
rect 451182 337560 451188 337572
rect 451240 337560 451246 337612
rect 453298 337560 453304 337612
rect 453356 337600 453362 337612
rect 453942 337600 453948 337612
rect 453356 337572 453948 337600
rect 453356 337560 453362 337572
rect 453942 337560 453948 337572
rect 454000 337560 454006 337612
rect 456981 337603 457039 337609
rect 456981 337569 456993 337603
rect 457027 337600 457039 337603
rect 460385 337603 460443 337609
rect 460385 337600 460397 337603
rect 457027 337572 460397 337600
rect 457027 337569 457039 337572
rect 456981 337563 457039 337569
rect 460385 337569 460397 337572
rect 460431 337569 460443 337603
rect 460385 337563 460443 337569
rect 461581 337603 461639 337609
rect 461581 337569 461593 337603
rect 461627 337600 461639 337603
rect 521010 337600 521016 337612
rect 461627 337572 521016 337600
rect 461627 337569 461639 337572
rect 461581 337563 461639 337569
rect 521010 337560 521016 337572
rect 521068 337560 521074 337612
rect 373960 337504 374776 337532
rect 373960 337492 373966 337504
rect 375282 337492 375288 337544
rect 375340 337532 375346 337544
rect 383746 337532 383752 337544
rect 375340 337504 383752 337532
rect 375340 337492 375346 337504
rect 383746 337492 383752 337504
rect 383804 337492 383810 337544
rect 405826 337492 405832 337544
rect 405884 337532 405890 337544
rect 426434 337532 426440 337544
rect 405884 337504 426440 337532
rect 405884 337492 405890 337504
rect 426434 337492 426440 337504
rect 426492 337492 426498 337544
rect 431865 337535 431923 337541
rect 431865 337501 431877 337535
rect 431911 337532 431923 337535
rect 442258 337532 442264 337544
rect 431911 337504 442264 337532
rect 431911 337501 431923 337504
rect 431865 337495 431923 337501
rect 442258 337492 442264 337504
rect 442316 337492 442322 337544
rect 447502 337492 447508 337544
rect 447560 337532 447566 337544
rect 448422 337532 448428 337544
rect 447560 337504 448428 337532
rect 447560 337492 447566 337504
rect 448422 337492 448428 337504
rect 448480 337492 448486 337544
rect 451277 337535 451335 337541
rect 451277 337501 451289 337535
rect 451323 337532 451335 337535
rect 516778 337532 516784 337544
rect 451323 337504 516784 337532
rect 451323 337501 451335 337504
rect 451277 337495 451335 337501
rect 516778 337492 516784 337504
rect 516836 337492 516842 337544
rect 374454 337464 374460 337476
rect 372172 337436 374460 337464
rect 374454 337424 374460 337436
rect 374512 337424 374518 337476
rect 374641 337467 374699 337473
rect 374641 337433 374653 337467
rect 374687 337464 374699 337467
rect 381814 337464 381820 337476
rect 374687 337436 381820 337464
rect 374687 337433 374699 337436
rect 374641 337427 374699 337433
rect 381814 337424 381820 337436
rect 381872 337424 381878 337476
rect 387058 337424 387064 337476
rect 387116 337464 387122 337476
rect 388714 337464 388720 337476
rect 387116 337436 388720 337464
rect 387116 337424 387122 337436
rect 388714 337424 388720 337436
rect 388772 337424 388778 337476
rect 396994 337424 397000 337476
rect 397052 337464 397058 337476
rect 405918 337464 405924 337476
rect 397052 337436 405924 337464
rect 397052 337424 397058 337436
rect 405918 337424 405924 337436
rect 405976 337424 405982 337476
rect 409138 337424 409144 337476
rect 409196 337464 409202 337476
rect 433518 337464 433524 337476
rect 409196 337436 433524 337464
rect 409196 337424 409202 337436
rect 433518 337424 433524 337436
rect 433576 337424 433582 337476
rect 437658 337424 437664 337476
rect 437716 337464 437722 337476
rect 438670 337464 438676 337476
rect 437716 337436 438676 337464
rect 437716 337424 437722 337436
rect 438670 337424 438676 337436
rect 438728 337424 438734 337476
rect 443086 337424 443092 337476
rect 443144 337464 443150 337476
rect 514018 337464 514024 337476
rect 443144 337436 514024 337464
rect 443144 337424 443150 337436
rect 514018 337424 514024 337436
rect 514076 337424 514082 337476
rect 369762 337356 369768 337408
rect 369820 337396 369826 337408
rect 369857 337399 369915 337405
rect 369857 337396 369869 337399
rect 369820 337368 369869 337396
rect 369820 337356 369826 337368
rect 369857 337365 369869 337368
rect 369903 337365 369915 337399
rect 369857 337359 369915 337365
rect 382182 337356 382188 337408
rect 382240 337396 382246 337408
rect 386690 337396 386696 337408
rect 382240 337368 386696 337396
rect 382240 337356 382246 337368
rect 386690 337356 386696 337368
rect 386748 337356 386754 337408
rect 400950 337356 400956 337408
rect 401008 337396 401014 337408
rect 402238 337396 402244 337408
rect 401008 337368 402244 337396
rect 401008 337356 401014 337368
rect 402238 337356 402244 337368
rect 402296 337356 402302 337408
rect 409230 337356 409236 337408
rect 409288 337396 409294 337408
rect 433978 337396 433984 337408
rect 409288 337368 433984 337396
rect 409288 337356 409294 337368
rect 433978 337356 433984 337368
rect 434036 337356 434042 337408
rect 434254 337356 434260 337408
rect 434312 337396 434318 337408
rect 439498 337396 439504 337408
rect 434312 337368 439504 337396
rect 434312 337356 434318 337368
rect 439498 337356 439504 337368
rect 439556 337356 439562 337408
rect 443457 337399 443515 337405
rect 443457 337365 443469 337399
rect 443503 337396 443515 337399
rect 510614 337396 510620 337408
rect 443503 337368 510620 337396
rect 443503 337365 443515 337368
rect 443457 337359 443515 337365
rect 510614 337356 510620 337368
rect 510672 337356 510678 337408
rect 364536 337300 365024 337328
rect 321879 337232 333192 337260
rect 321879 337229 321891 337232
rect 321833 337223 321891 337229
rect 333238 337220 333244 337272
rect 333296 337260 333302 337272
rect 364996 337260 365024 337300
rect 367002 337288 367008 337340
rect 367060 337328 367066 337340
rect 380802 337328 380808 337340
rect 367060 337300 380808 337328
rect 367060 337288 367066 337300
rect 380802 337288 380808 337300
rect 380860 337288 380866 337340
rect 412637 337331 412695 337337
rect 412637 337297 412649 337331
rect 412683 337328 412695 337331
rect 412683 337300 417096 337328
rect 412683 337297 412695 337300
rect 412637 337291 412695 337297
rect 372982 337260 372988 337272
rect 333296 337232 363828 337260
rect 364996 337232 372988 337260
rect 333296 337220 333302 337232
rect 312538 337152 312544 337204
rect 312596 337192 312602 337204
rect 341705 337195 341763 337201
rect 341705 337192 341717 337195
rect 312596 337164 341717 337192
rect 312596 337152 312602 337164
rect 341705 337161 341717 337164
rect 341751 337161 341763 337195
rect 341705 337155 341763 337161
rect 341794 337152 341800 337204
rect 341852 337192 341858 337204
rect 348970 337192 348976 337204
rect 341852 337164 348976 337192
rect 341852 337152 341858 337164
rect 348970 337152 348976 337164
rect 349028 337152 349034 337204
rect 359458 337152 359464 337204
rect 359516 337192 359522 337204
rect 363690 337192 363696 337204
rect 359516 337164 363696 337192
rect 359516 337152 359522 337164
rect 363690 337152 363696 337164
rect 363748 337152 363754 337204
rect 363800 337192 363828 337232
rect 372982 337220 372988 337232
rect 373040 337220 373046 337272
rect 366634 337192 366640 337204
rect 363800 337164 366640 337192
rect 366634 337152 366640 337164
rect 366692 337152 366698 337204
rect 369857 337195 369915 337201
rect 369857 337161 369869 337195
rect 369903 337192 369915 337195
rect 374641 337195 374699 337201
rect 374641 337192 374653 337195
rect 369903 337164 374653 337192
rect 369903 337161 369915 337164
rect 369857 337155 369915 337161
rect 374641 337161 374653 337164
rect 374687 337161 374699 337195
rect 374641 337155 374699 337161
rect 401870 337152 401876 337204
rect 401928 337192 401934 337204
rect 416958 337192 416964 337204
rect 401928 337164 416964 337192
rect 401928 337152 401934 337164
rect 416958 337152 416964 337164
rect 417016 337152 417022 337204
rect 417068 337192 417096 337300
rect 419994 337288 420000 337340
rect 420052 337328 420058 337340
rect 420730 337328 420736 337340
rect 420052 337300 420736 337328
rect 420052 337288 420058 337300
rect 420730 337288 420736 337300
rect 420788 337288 420794 337340
rect 421006 337288 421012 337340
rect 421064 337328 421070 337340
rect 456981 337331 457039 337337
rect 456981 337328 456993 337331
rect 421064 337300 456993 337328
rect 421064 337288 421070 337300
rect 456981 337297 456993 337300
rect 457027 337297 457039 337331
rect 461581 337331 461639 337337
rect 461581 337328 461593 337331
rect 456981 337291 457039 337297
rect 457088 337300 461593 337328
rect 423490 337220 423496 337272
rect 423548 337260 423554 337272
rect 457088 337260 457116 337300
rect 461581 337297 461593 337300
rect 461627 337297 461639 337331
rect 463878 337328 463884 337340
rect 461581 337291 461639 337297
rect 461688 337300 463884 337328
rect 423548 337232 457116 337260
rect 457165 337263 457223 337269
rect 423548 337220 423554 337232
rect 457165 337229 457177 337263
rect 457211 337260 457223 337263
rect 460290 337260 460296 337272
rect 457211 337232 460296 337260
rect 457211 337229 457223 337232
rect 457165 337223 457223 337229
rect 460290 337220 460296 337232
rect 460348 337220 460354 337272
rect 460385 337263 460443 337269
rect 460385 337229 460397 337263
rect 460431 337260 460443 337263
rect 461688 337260 461716 337300
rect 463878 337288 463884 337300
rect 463936 337288 463942 337340
rect 465074 337288 465080 337340
rect 465132 337328 465138 337340
rect 466362 337328 466368 337340
rect 465132 337300 466368 337328
rect 465132 337288 465138 337300
rect 466362 337288 466368 337300
rect 466420 337288 466426 337340
rect 466457 337331 466515 337337
rect 466457 337297 466469 337331
rect 466503 337328 466515 337331
rect 470594 337328 470600 337340
rect 466503 337300 470600 337328
rect 466503 337297 466515 337300
rect 466457 337291 466515 337297
rect 470594 337288 470600 337300
rect 470652 337288 470658 337340
rect 470686 337288 470692 337340
rect 470744 337328 470750 337340
rect 529198 337328 529204 337340
rect 470744 337300 529204 337328
rect 470744 337288 470750 337300
rect 529198 337288 529204 337300
rect 529256 337288 529262 337340
rect 460431 337232 461716 337260
rect 460431 337229 460443 337232
rect 460385 337223 460443 337229
rect 463602 337220 463608 337272
rect 463660 337260 463666 337272
rect 469217 337263 469275 337269
rect 469217 337260 469229 337263
rect 463660 337232 469229 337260
rect 463660 337220 463666 337232
rect 469217 337229 469229 337232
rect 469263 337229 469275 337263
rect 469217 337223 469275 337229
rect 469490 337220 469496 337272
rect 469548 337260 469554 337272
rect 530578 337260 530584 337272
rect 469548 337232 530584 337260
rect 469548 337220 469554 337232
rect 530578 337220 530584 337232
rect 530636 337220 530642 337272
rect 424318 337192 424324 337204
rect 417068 337164 424324 337192
rect 424318 337152 424324 337164
rect 424376 337152 424382 337204
rect 427906 337152 427912 337204
rect 427964 337192 427970 337204
rect 431865 337195 431923 337201
rect 431865 337192 431877 337195
rect 427964 337164 431877 337192
rect 427964 337152 427970 337164
rect 431865 337161 431877 337164
rect 431911 337161 431923 337195
rect 431865 337155 431923 337161
rect 432782 337152 432788 337204
rect 432840 337192 432846 337204
rect 492674 337192 492680 337204
rect 432840 337164 492680 337192
rect 432840 337152 432846 337164
rect 492674 337152 492680 337164
rect 492732 337152 492738 337204
rect 314194 337124 314200 337136
rect 302344 337096 314200 337124
rect 314194 337084 314200 337096
rect 314252 337084 314258 337136
rect 316678 337084 316684 337136
rect 316736 337124 316742 337136
rect 342809 337127 342867 337133
rect 342809 337124 342821 337127
rect 316736 337096 342821 337124
rect 316736 337084 316742 337096
rect 342809 337093 342821 337096
rect 342855 337093 342867 337127
rect 342809 337087 342867 337093
rect 342898 337084 342904 337136
rect 342956 337124 342962 337136
rect 345845 337127 345903 337133
rect 345845 337124 345857 337127
rect 342956 337096 345857 337124
rect 342956 337084 342962 337096
rect 345845 337093 345857 337096
rect 345891 337093 345903 337127
rect 345845 337087 345903 337093
rect 355962 337084 355968 337136
rect 356020 337124 356026 337136
rect 364981 337127 365039 337133
rect 364981 337124 364993 337127
rect 356020 337096 364993 337124
rect 356020 337084 356026 337096
rect 364981 337093 364993 337096
rect 365027 337093 365039 337127
rect 364981 337087 365039 337093
rect 369118 337084 369124 337136
rect 369176 337124 369182 337136
rect 371050 337124 371056 337136
rect 369176 337096 371056 337124
rect 369176 337084 369182 337096
rect 371050 337084 371056 337096
rect 371108 337084 371114 337136
rect 415118 337084 415124 337136
rect 415176 337124 415182 337136
rect 421558 337124 421564 337136
rect 415176 337096 421564 337124
rect 415176 337084 415182 337096
rect 421558 337084 421564 337096
rect 421616 337084 421622 337136
rect 429838 337084 429844 337136
rect 429896 337124 429902 337136
rect 485774 337124 485780 337136
rect 429896 337096 485780 337124
rect 429896 337084 429902 337096
rect 485774 337084 485780 337096
rect 485832 337084 485838 337136
rect 95878 337016 95884 337068
rect 95936 337056 95942 337068
rect 265250 337056 265256 337068
rect 95936 337028 265256 337056
rect 95936 337016 95942 337028
rect 265250 337016 265256 337028
rect 265308 337016 265314 337068
rect 335262 337016 335268 337068
rect 335320 337056 335326 337068
rect 367646 337056 367652 337068
rect 335320 337028 367652 337056
rect 335320 337016 335326 337028
rect 367646 337016 367652 337028
rect 367704 337016 367710 337068
rect 397454 337016 397460 337068
rect 397512 337056 397518 337068
rect 403618 337056 403624 337068
rect 397512 337028 403624 337056
rect 397512 337016 397518 337028
rect 403618 337016 403624 337028
rect 403676 337016 403682 337068
rect 407758 337016 407764 337068
rect 407816 337056 407822 337068
rect 409138 337056 409144 337068
rect 407816 337028 409144 337056
rect 407816 337016 407822 337028
rect 409138 337016 409144 337028
rect 409196 337016 409202 337068
rect 426894 337016 426900 337068
rect 426952 337056 426958 337068
rect 477586 337056 477592 337068
rect 426952 337028 477592 337056
rect 426952 337016 426958 337028
rect 477586 337016 477592 337028
rect 477644 337016 477650 337068
rect 103425 336991 103483 336997
rect 103425 336988 103437 336991
rect 93872 336960 103437 336988
rect 86957 336951 87015 336957
rect 103425 336957 103437 336960
rect 103471 336957 103483 336991
rect 103425 336951 103483 336957
rect 107562 336948 107568 337000
rect 107620 336988 107626 337000
rect 274082 336988 274088 337000
rect 107620 336960 274088 336988
rect 107620 336948 107626 336960
rect 274082 336948 274088 336960
rect 274140 336948 274146 337000
rect 319438 336948 319444 337000
rect 319496 336988 319502 337000
rect 345753 336991 345811 336997
rect 345753 336988 345765 336991
rect 319496 336960 345765 336988
rect 319496 336948 319502 336960
rect 345753 336957 345765 336960
rect 345799 336957 345811 336991
rect 345753 336951 345811 336957
rect 345845 336991 345903 336997
rect 345845 336957 345857 336991
rect 345891 336988 345903 336991
rect 353386 336988 353392 337000
rect 345891 336960 353392 336988
rect 345891 336957 345903 336960
rect 345845 336951 345903 336957
rect 353386 336948 353392 336960
rect 353444 336948 353450 337000
rect 378042 336948 378048 337000
rect 378100 336988 378106 337000
rect 385218 336988 385224 337000
rect 378100 336960 385224 336988
rect 378100 336948 378106 336960
rect 385218 336948 385224 336960
rect 385276 336948 385282 337000
rect 401410 336948 401416 337000
rect 401468 336988 401474 337000
rect 404998 336988 405004 337000
rect 401468 336960 405004 336988
rect 401468 336948 401474 336960
rect 404998 336948 405004 336960
rect 405056 336948 405062 337000
rect 432233 336991 432291 336997
rect 432233 336957 432245 336991
rect 432279 336988 432291 336991
rect 475378 336988 475384 337000
rect 432279 336960 475384 336988
rect 432279 336957 432291 336960
rect 432233 336951 432291 336957
rect 475378 336948 475384 336960
rect 475436 336948 475442 337000
rect 102778 336880 102784 336932
rect 102836 336920 102842 336932
rect 268194 336920 268200 336932
rect 102836 336892 268200 336920
rect 102836 336880 102842 336892
rect 268194 336880 268200 336892
rect 268252 336880 268258 336932
rect 345474 336920 345480 336932
rect 335740 336892 345480 336920
rect 118602 336812 118608 336864
rect 118660 336852 118666 336864
rect 278498 336852 278504 336864
rect 118660 336824 278504 336852
rect 118660 336812 118666 336824
rect 278498 336812 278504 336824
rect 278556 336812 278562 336864
rect 113177 336787 113235 336793
rect 113177 336753 113189 336787
rect 113223 336784 113235 336787
rect 122745 336787 122803 336793
rect 122745 336784 122757 336787
rect 113223 336756 122757 336784
rect 113223 336753 113235 336756
rect 113177 336747 113235 336753
rect 122745 336753 122757 336756
rect 122791 336753 122803 336787
rect 122745 336747 122803 336753
rect 125502 336744 125508 336796
rect 125560 336784 125566 336796
rect 281166 336784 281172 336796
rect 125560 336756 281172 336784
rect 125560 336744 125566 336756
rect 281166 336744 281172 336756
rect 281224 336744 281230 336796
rect 327718 336744 327724 336796
rect 327776 336784 327782 336796
rect 335740 336784 335768 336892
rect 345474 336880 345480 336892
rect 345532 336880 345538 336932
rect 345934 336880 345940 336932
rect 345992 336920 345998 336932
rect 360286 336920 360292 336932
rect 345992 336892 360292 336920
rect 345992 336880 345998 336892
rect 360286 336880 360292 336892
rect 360344 336880 360350 336932
rect 380802 336880 380808 336932
rect 380860 336920 380866 336932
rect 386230 336920 386236 336932
rect 380860 336892 386236 336920
rect 380860 336880 380866 336892
rect 386230 336880 386236 336892
rect 386288 336880 386294 336932
rect 392118 336880 392124 336932
rect 392176 336920 392182 336932
rect 393590 336920 393596 336932
rect 392176 336892 393596 336920
rect 392176 336880 392182 336892
rect 393590 336880 393596 336892
rect 393648 336880 393654 336932
rect 393866 336880 393872 336932
rect 393924 336920 393930 336932
rect 397454 336920 397460 336932
rect 393924 336892 397460 336920
rect 393924 336880 393930 336892
rect 397454 336880 397460 336892
rect 397512 336880 397518 336932
rect 423950 336880 423956 336932
rect 424008 336920 424014 336932
rect 466457 336923 466515 336929
rect 466457 336920 466469 336923
rect 424008 336892 466469 336920
rect 424008 336880 424014 336892
rect 466457 336889 466469 336892
rect 466503 336889 466515 336923
rect 466457 336883 466515 336889
rect 466546 336880 466552 336932
rect 466604 336920 466610 336932
rect 470502 336920 470508 336932
rect 466604 336892 470508 336920
rect 466604 336880 466610 336892
rect 470502 336880 470508 336892
rect 470560 336880 470566 336932
rect 344278 336812 344284 336864
rect 344336 336852 344342 336864
rect 357342 336852 357348 336864
rect 344336 336824 357348 336852
rect 344336 336812 344342 336824
rect 357342 336812 357348 336824
rect 357400 336812 357406 336864
rect 362218 336812 362224 336864
rect 362276 336852 362282 336864
rect 365162 336852 365168 336864
rect 362276 336824 365168 336852
rect 362276 336812 362282 336824
rect 365162 336812 365168 336824
rect 365220 336812 365226 336864
rect 381630 336812 381636 336864
rect 381688 336852 381694 336864
rect 384758 336852 384764 336864
rect 381688 336824 384764 336852
rect 381688 336812 381694 336824
rect 384758 336812 384764 336824
rect 384816 336812 384822 336864
rect 396074 336812 396080 336864
rect 396132 336852 396138 336864
rect 398190 336852 398196 336864
rect 396132 336824 398196 336852
rect 396132 336812 396138 336824
rect 398190 336812 398196 336824
rect 398248 336812 398254 336864
rect 424962 336812 424968 336864
rect 425020 336852 425026 336864
rect 439590 336852 439596 336864
rect 425020 336824 439596 336852
rect 425020 336812 425026 336824
rect 439590 336812 439596 336824
rect 439648 336812 439654 336864
rect 441614 336812 441620 336864
rect 441672 336852 441678 336864
rect 443638 336852 443644 336864
rect 441672 336824 443644 336852
rect 441672 336812 441678 336824
rect 443638 336812 443644 336824
rect 443696 336812 443702 336864
rect 456794 336812 456800 336864
rect 456852 336852 456858 336864
rect 458082 336852 458088 336864
rect 456852 336824 458088 336852
rect 456852 336812 456858 336824
rect 458082 336812 458088 336824
rect 458140 336812 458146 336864
rect 459186 336812 459192 336864
rect 459244 336852 459250 336864
rect 460198 336852 460204 336864
rect 459244 336824 460204 336852
rect 459244 336812 459250 336824
rect 460198 336812 460204 336824
rect 460256 336812 460262 336864
rect 461581 336855 461639 336861
rect 461581 336821 461593 336855
rect 461627 336852 461639 336855
rect 469214 336852 469220 336864
rect 461627 336824 469220 336852
rect 461627 336821 461639 336824
rect 461581 336815 461639 336821
rect 469214 336812 469220 336824
rect 469272 336812 469278 336864
rect 509878 336852 509884 336864
rect 469324 336824 509884 336852
rect 327776 336756 335768 336784
rect 335817 336787 335875 336793
rect 327776 336744 327782 336756
rect 335817 336753 335829 336787
rect 335863 336784 335875 336787
rect 343082 336784 343088 336796
rect 335863 336756 343088 336784
rect 335863 336753 335875 336756
rect 335817 336747 335875 336753
rect 343082 336744 343088 336756
rect 343140 336744 343146 336796
rect 345569 336787 345627 336793
rect 345569 336784 345581 336787
rect 343192 336756 345581 336784
rect 251818 336676 251824 336728
rect 251876 336716 251882 336728
rect 256418 336716 256424 336728
rect 251876 336688 256424 336716
rect 251876 336676 251882 336688
rect 256418 336676 256424 336688
rect 256476 336676 256482 336728
rect 330205 336719 330263 336725
rect 330205 336685 330217 336719
rect 330251 336716 330263 336719
rect 330570 336716 330576 336728
rect 330251 336688 330576 336716
rect 330251 336685 330263 336688
rect 330205 336679 330263 336685
rect 330570 336676 330576 336688
rect 330628 336676 330634 336728
rect 341705 336719 341763 336725
rect 341705 336685 341717 336719
rect 341751 336716 341763 336719
rect 343192 336716 343220 336756
rect 345569 336753 345581 336756
rect 345615 336753 345627 336787
rect 345569 336747 345627 336753
rect 345753 336787 345811 336793
rect 345753 336753 345765 336787
rect 345799 336784 345811 336787
rect 351454 336784 351460 336796
rect 345799 336756 351460 336784
rect 345799 336753 345811 336756
rect 345753 336747 345811 336753
rect 351454 336744 351460 336756
rect 351512 336744 351518 336796
rect 352558 336744 352564 336796
rect 352616 336784 352622 336796
rect 357802 336784 357808 336796
rect 352616 336756 357808 336784
rect 352616 336744 352622 336756
rect 357802 336744 357808 336756
rect 357860 336744 357866 336796
rect 363598 336744 363604 336796
rect 363656 336784 363662 336796
rect 364702 336784 364708 336796
rect 363656 336756 364708 336784
rect 363656 336744 363662 336756
rect 364702 336744 364708 336756
rect 364760 336744 364766 336796
rect 370498 336744 370504 336796
rect 370556 336784 370562 336796
rect 372522 336784 372528 336796
rect 370556 336756 372528 336784
rect 370556 336744 370562 336756
rect 372522 336744 372528 336756
rect 372580 336744 372586 336796
rect 376018 336744 376024 336796
rect 376076 336784 376082 336796
rect 376938 336784 376944 336796
rect 376076 336756 376944 336784
rect 376076 336744 376082 336756
rect 376938 336744 376944 336756
rect 376996 336744 377002 336796
rect 377674 336744 377680 336796
rect 377732 336784 377738 336796
rect 378410 336784 378416 336796
rect 377732 336756 378416 336784
rect 377732 336744 377738 336756
rect 378410 336744 378416 336756
rect 378468 336744 378474 336796
rect 394050 336744 394056 336796
rect 394108 336784 394114 336796
rect 394602 336784 394608 336796
rect 394108 336756 394608 336784
rect 394108 336744 394114 336756
rect 394602 336744 394608 336756
rect 394660 336744 394666 336796
rect 395062 336744 395068 336796
rect 395120 336784 395126 336796
rect 395890 336784 395896 336796
rect 395120 336756 395896 336784
rect 395120 336744 395126 336756
rect 395890 336744 395896 336756
rect 395948 336744 395954 336796
rect 396534 336744 396540 336796
rect 396592 336784 396598 336796
rect 398098 336784 398104 336796
rect 396592 336756 398104 336784
rect 396592 336744 396598 336756
rect 398098 336744 398104 336756
rect 398156 336744 398162 336796
rect 424594 336744 424600 336796
rect 424652 336784 424658 336796
rect 454681 336787 454739 336793
rect 424652 336756 425008 336784
rect 424652 336744 424658 336756
rect 424980 336728 425008 336756
rect 454681 336753 454693 336787
rect 454727 336784 454739 336787
rect 457165 336787 457223 336793
rect 457165 336784 457177 336787
rect 454727 336756 457177 336784
rect 454727 336753 454739 336756
rect 454681 336747 454739 336753
rect 457165 336753 457177 336756
rect 457211 336753 457223 336787
rect 457165 336747 457223 336753
rect 457254 336744 457260 336796
rect 457312 336784 457318 336796
rect 457990 336784 457996 336796
rect 457312 336756 457996 336784
rect 457312 336744 457318 336756
rect 457990 336744 457996 336756
rect 458048 336744 458054 336796
rect 458266 336744 458272 336796
rect 458324 336784 458330 336796
rect 459462 336784 459468 336796
rect 458324 336756 459468 336784
rect 458324 336744 458330 336756
rect 459462 336744 459468 336756
rect 459520 336744 459526 336796
rect 459738 336744 459744 336796
rect 459796 336784 459802 336796
rect 460842 336784 460848 336796
rect 459796 336756 460848 336784
rect 459796 336744 459802 336756
rect 460842 336744 460848 336756
rect 460900 336744 460906 336796
rect 461210 336744 461216 336796
rect 461268 336784 461274 336796
rect 462130 336784 462136 336796
rect 461268 336756 462136 336784
rect 461268 336744 461274 336756
rect 462130 336744 462136 336756
rect 462188 336744 462194 336796
rect 462682 336744 462688 336796
rect 462740 336784 462746 336796
rect 463510 336784 463516 336796
rect 462740 336756 463516 336784
rect 462740 336744 462746 336756
rect 463510 336744 463516 336756
rect 463568 336744 463574 336796
rect 464154 336744 464160 336796
rect 464212 336784 464218 336796
rect 464982 336784 464988 336796
rect 464212 336756 464988 336784
rect 464212 336744 464218 336756
rect 464982 336744 464988 336756
rect 465040 336744 465046 336796
rect 465074 336744 465080 336796
rect 465132 336784 465138 336796
rect 469324 336784 469352 336824
rect 509878 336812 509884 336824
rect 509936 336812 509942 336864
rect 505738 336784 505744 336796
rect 465132 336756 469352 336784
rect 469416 336756 505744 336784
rect 465132 336744 465138 336756
rect 341751 336688 343220 336716
rect 374457 336719 374515 336725
rect 341751 336685 341763 336688
rect 341705 336679 341763 336685
rect 374457 336685 374469 336719
rect 374503 336716 374515 336719
rect 374546 336716 374552 336728
rect 374503 336688 374552 336716
rect 374503 336685 374515 336688
rect 374457 336679 374515 336685
rect 374546 336676 374552 336688
rect 374604 336676 374610 336728
rect 375834 336716 375840 336728
rect 375795 336688 375840 336716
rect 375834 336676 375840 336688
rect 375892 336676 375898 336728
rect 424962 336676 424968 336728
rect 425020 336676 425026 336728
rect 466273 336719 466331 336725
rect 466273 336685 466285 336719
rect 466319 336716 466331 336719
rect 469416 336716 469444 336756
rect 505738 336744 505744 336756
rect 505796 336744 505802 336796
rect 466319 336688 469444 336716
rect 466319 336685 466331 336688
rect 466273 336679 466331 336685
rect 247678 336472 247684 336524
rect 247736 336512 247742 336524
rect 248598 336512 248604 336524
rect 247736 336484 248604 336512
rect 247736 336472 247742 336484
rect 248598 336472 248604 336484
rect 248656 336472 248662 336524
rect 249058 336200 249064 336252
rect 249116 336240 249122 336252
rect 250530 336240 250536 336252
rect 249116 336212 250536 336240
rect 249116 336200 249122 336212
rect 250530 336200 250536 336212
rect 250588 336200 250594 336252
rect 331398 336104 331404 336116
rect 331359 336076 331404 336104
rect 331398 336064 331404 336076
rect 331456 336064 331462 336116
rect 331214 335860 331220 335912
rect 331272 335900 331278 335912
rect 331490 335900 331496 335912
rect 331272 335872 331496 335900
rect 331272 335860 331278 335872
rect 331490 335860 331496 335872
rect 331548 335860 331554 335912
rect 236178 335656 236184 335708
rect 236236 335696 236242 335708
rect 237006 335696 237012 335708
rect 236236 335668 237012 335696
rect 236236 335656 236242 335668
rect 237006 335656 237012 335668
rect 237064 335656 237070 335708
rect 302234 335656 302240 335708
rect 302292 335696 302298 335708
rect 302694 335696 302700 335708
rect 302292 335668 302700 335696
rect 302292 335656 302298 335668
rect 302694 335656 302700 335668
rect 302752 335656 302758 335708
rect 316034 335656 316040 335708
rect 316092 335696 316098 335708
rect 316862 335696 316868 335708
rect 316092 335668 316868 335696
rect 316092 335656 316098 335668
rect 316862 335656 316868 335668
rect 316920 335656 316926 335708
rect 318794 335656 318800 335708
rect 318852 335696 318858 335708
rect 319806 335696 319812 335708
rect 318852 335668 319812 335696
rect 318852 335656 318858 335668
rect 319806 335656 319812 335668
rect 319864 335656 319870 335708
rect 332686 335656 332692 335708
rect 332744 335696 332750 335708
rect 333422 335696 333428 335708
rect 332744 335668 333428 335696
rect 332744 335656 332750 335668
rect 333422 335656 333428 335668
rect 333480 335656 333486 335708
rect 334066 335656 334072 335708
rect 334124 335696 334130 335708
rect 334894 335696 334900 335708
rect 334124 335668 334900 335696
rect 334124 335656 334130 335668
rect 334894 335656 334900 335668
rect 334952 335656 334958 335708
rect 236086 335588 236092 335640
rect 236144 335628 236150 335640
rect 236546 335628 236552 335640
rect 236144 335600 236552 335628
rect 236144 335588 236150 335600
rect 236546 335588 236552 335600
rect 236604 335588 236610 335640
rect 241606 335588 241612 335640
rect 241664 335628 241670 335640
rect 242342 335628 242348 335640
rect 241664 335600 242348 335628
rect 241664 335588 241670 335600
rect 242342 335588 242348 335600
rect 242400 335588 242406 335640
rect 260926 335588 260932 335640
rect 260984 335628 260990 335640
rect 261478 335628 261484 335640
rect 260984 335600 261484 335628
rect 260984 335588 260990 335600
rect 261478 335588 261484 335600
rect 261536 335588 261542 335640
rect 263686 335588 263692 335640
rect 263744 335628 263750 335640
rect 264422 335628 264428 335640
rect 263744 335600 264428 335628
rect 263744 335588 263750 335600
rect 264422 335588 264428 335600
rect 264480 335588 264486 335640
rect 265066 335588 265072 335640
rect 265124 335628 265130 335640
rect 265894 335628 265900 335640
rect 265124 335600 265900 335628
rect 265124 335588 265130 335600
rect 265894 335588 265900 335600
rect 265952 335588 265958 335640
rect 266446 335588 266452 335640
rect 266504 335628 266510 335640
rect 267366 335628 267372 335640
rect 266504 335600 267372 335628
rect 266504 335588 266510 335600
rect 267366 335588 267372 335600
rect 267424 335588 267430 335640
rect 280246 335588 280252 335640
rect 280304 335628 280310 335640
rect 280614 335628 280620 335640
rect 280304 335600 280620 335628
rect 280304 335588 280310 335600
rect 280614 335588 280620 335600
rect 280672 335588 280678 335640
rect 281534 335588 281540 335640
rect 281592 335628 281598 335640
rect 282086 335628 282092 335640
rect 281592 335600 282092 335628
rect 281592 335588 281598 335600
rect 282086 335588 282092 335600
rect 282144 335588 282150 335640
rect 283006 335588 283012 335640
rect 283064 335628 283070 335640
rect 283558 335628 283564 335640
rect 283064 335600 283564 335628
rect 283064 335588 283070 335600
rect 283558 335588 283564 335600
rect 283616 335588 283622 335640
rect 285674 335588 285680 335640
rect 285732 335628 285738 335640
rect 285950 335628 285956 335640
rect 285732 335600 285956 335628
rect 285732 335588 285738 335600
rect 285950 335588 285956 335600
rect 286008 335588 286014 335640
rect 286042 335588 286048 335640
rect 286100 335628 286106 335640
rect 286594 335628 286600 335640
rect 286100 335600 286600 335628
rect 286100 335588 286106 335600
rect 286594 335588 286600 335600
rect 286652 335588 286658 335640
rect 287054 335588 287060 335640
rect 287112 335628 287118 335640
rect 287974 335628 287980 335640
rect 287112 335600 287980 335628
rect 287112 335588 287118 335600
rect 287974 335588 287980 335600
rect 288032 335588 288038 335640
rect 288434 335588 288440 335640
rect 288492 335628 288498 335640
rect 289446 335628 289452 335640
rect 288492 335600 289452 335628
rect 288492 335588 288498 335600
rect 289446 335588 289452 335600
rect 289504 335588 289510 335640
rect 292758 335588 292764 335640
rect 292816 335628 292822 335640
rect 293310 335628 293316 335640
rect 292816 335600 293316 335628
rect 292816 335588 292822 335600
rect 293310 335588 293316 335600
rect 293368 335588 293374 335640
rect 298278 335588 298284 335640
rect 298336 335628 298342 335640
rect 298646 335628 298652 335640
rect 298336 335600 298652 335628
rect 298336 335588 298342 335600
rect 298646 335588 298652 335600
rect 298704 335588 298710 335640
rect 300854 335588 300860 335640
rect 300912 335628 300918 335640
rect 301222 335628 301228 335640
rect 300912 335600 301228 335628
rect 300912 335588 300918 335600
rect 301222 335588 301228 335600
rect 301280 335588 301286 335640
rect 303614 335588 303620 335640
rect 303672 335628 303678 335640
rect 304166 335628 304172 335640
rect 303672 335600 304172 335628
rect 303672 335588 303678 335600
rect 304166 335588 304172 335600
rect 304224 335588 304230 335640
rect 307754 335588 307760 335640
rect 307812 335628 307818 335640
rect 308582 335628 308588 335640
rect 307812 335600 308588 335628
rect 307812 335588 307818 335600
rect 308582 335588 308588 335600
rect 308640 335588 308646 335640
rect 309134 335588 309140 335640
rect 309192 335628 309198 335640
rect 310054 335628 310060 335640
rect 309192 335600 310060 335628
rect 309192 335588 309198 335600
rect 310054 335588 310060 335600
rect 310112 335588 310118 335640
rect 310514 335588 310520 335640
rect 310572 335628 310578 335640
rect 311526 335628 311532 335640
rect 310572 335600 311532 335628
rect 310572 335588 310578 335600
rect 311526 335588 311532 335600
rect 311584 335588 311590 335640
rect 314654 335588 314660 335640
rect 314712 335628 314718 335640
rect 315390 335628 315396 335640
rect 314712 335600 315396 335628
rect 314712 335588 314718 335600
rect 315390 335588 315396 335600
rect 315448 335588 315454 335640
rect 316126 335588 316132 335640
rect 316184 335628 316190 335640
rect 316310 335628 316316 335640
rect 316184 335600 316316 335628
rect 316184 335588 316190 335600
rect 316310 335588 316316 335600
rect 316368 335588 316374 335640
rect 317414 335588 317420 335640
rect 317472 335628 317478 335640
rect 318334 335628 318340 335640
rect 317472 335600 318340 335628
rect 317472 335588 317478 335600
rect 318334 335588 318340 335600
rect 318392 335588 318398 335640
rect 318886 335588 318892 335640
rect 318944 335628 318950 335640
rect 319254 335628 319260 335640
rect 318944 335600 319260 335628
rect 318944 335588 318950 335600
rect 319254 335588 319260 335600
rect 319312 335588 319318 335640
rect 320174 335588 320180 335640
rect 320232 335628 320238 335640
rect 320726 335628 320732 335640
rect 320232 335600 320732 335628
rect 320232 335588 320238 335600
rect 320726 335588 320732 335600
rect 320784 335588 320790 335640
rect 321646 335588 321652 335640
rect 321704 335628 321710 335640
rect 322198 335628 322204 335640
rect 321704 335600 322204 335628
rect 321704 335588 321710 335600
rect 322198 335588 322204 335600
rect 322256 335588 322262 335640
rect 329834 335588 329840 335640
rect 329892 335628 329898 335640
rect 330110 335628 330116 335640
rect 329892 335600 330116 335628
rect 329892 335588 329898 335600
rect 330110 335588 330116 335600
rect 330168 335588 330174 335640
rect 332594 335588 332600 335640
rect 332652 335628 332658 335640
rect 333054 335628 333060 335640
rect 332652 335600 333060 335628
rect 332652 335588 332658 335600
rect 333054 335588 333060 335600
rect 333112 335588 333118 335640
rect 333974 335588 333980 335640
rect 334032 335628 334038 335640
rect 334526 335628 334532 335640
rect 334032 335600 334532 335628
rect 334032 335588 334038 335600
rect 334526 335588 334532 335600
rect 334584 335588 334590 335640
rect 338114 335588 338120 335640
rect 338172 335628 338178 335640
rect 338942 335628 338948 335640
rect 338172 335600 338948 335628
rect 338172 335588 338178 335600
rect 338942 335588 338948 335600
rect 339000 335588 339006 335640
rect 356146 335588 356152 335640
rect 356204 335628 356210 335640
rect 356606 335628 356612 335640
rect 356204 335600 356612 335628
rect 356204 335588 356210 335600
rect 356606 335588 356612 335600
rect 356664 335588 356670 335640
rect 358998 335588 359004 335640
rect 359056 335628 359062 335640
rect 359366 335628 359372 335640
rect 359056 335600 359372 335628
rect 359056 335588 359062 335600
rect 359366 335588 359372 335600
rect 359424 335588 359430 335640
rect 363046 335588 363052 335640
rect 363104 335628 363110 335640
rect 363782 335628 363788 335640
rect 363104 335600 363788 335628
rect 363104 335588 363110 335600
rect 363782 335588 363788 335600
rect 363840 335588 363846 335640
rect 367278 335588 367284 335640
rect 367336 335628 367342 335640
rect 367922 335628 367928 335640
rect 367336 335600 367928 335628
rect 367336 335588 367342 335600
rect 367922 335588 367928 335600
rect 367980 335588 367986 335640
rect 458910 335588 458916 335640
rect 458968 335628 458974 335640
rect 459370 335628 459376 335640
rect 458968 335600 459376 335628
rect 458968 335588 458974 335600
rect 459370 335588 459376 335600
rect 459428 335588 459434 335640
rect 341702 335560 341708 335572
rect 341663 335532 341708 335560
rect 341702 335520 341708 335532
rect 341760 335520 341766 335572
rect 235074 335452 235080 335504
rect 235132 335492 235138 335504
rect 235626 335492 235632 335504
rect 235132 335464 235632 335492
rect 235132 335452 235138 335464
rect 235626 335452 235632 335464
rect 235684 335452 235690 335504
rect 245838 335452 245844 335504
rect 245896 335492 245902 335504
rect 246666 335492 246672 335504
rect 245896 335464 246672 335492
rect 245896 335452 245902 335464
rect 246666 335452 246672 335464
rect 246724 335452 246730 335504
rect 331306 335452 331312 335504
rect 331364 335492 331370 335504
rect 331950 335492 331956 335504
rect 331364 335464 331956 335492
rect 331364 335452 331370 335464
rect 331950 335452 331956 335464
rect 332008 335452 332014 335504
rect 580074 335384 580080 335436
rect 580132 335424 580138 335436
rect 580994 335424 581000 335436
rect 580132 335396 581000 335424
rect 580132 335384 580138 335396
rect 580994 335384 581000 335396
rect 581052 335384 581058 335436
rect 580074 335248 580080 335300
rect 580132 335288 580138 335300
rect 580994 335288 581000 335300
rect 580132 335260 581000 335288
rect 580132 335248 580138 335260
rect 580994 335248 581000 335260
rect 581052 335248 581058 335300
rect 284389 335223 284447 335229
rect 284389 335189 284401 335223
rect 284435 335220 284447 335223
rect 284478 335220 284484 335232
rect 284435 335192 284484 335220
rect 284435 335189 284447 335192
rect 284389 335183 284447 335189
rect 284478 335180 284484 335192
rect 284536 335180 284542 335232
rect 278774 334772 278780 334824
rect 278832 334812 278838 334824
rect 278958 334812 278964 334824
rect 278832 334784 278964 334812
rect 278832 334772 278838 334784
rect 278958 334772 278964 334784
rect 279016 334772 279022 334824
rect 302513 334747 302571 334753
rect 302513 334713 302525 334747
rect 302559 334744 302571 334747
rect 303062 334744 303068 334756
rect 302559 334716 303068 334744
rect 302559 334713 302571 334716
rect 302513 334707 302571 334713
rect 303062 334704 303068 334716
rect 303120 334704 303126 334756
rect 258166 334568 258172 334620
rect 258224 334608 258230 334620
rect 258534 334608 258540 334620
rect 258224 334580 258540 334608
rect 258224 334568 258230 334580
rect 258534 334568 258540 334580
rect 258592 334568 258598 334620
rect 328546 334500 328552 334552
rect 328604 334540 328610 334552
rect 329006 334540 329012 334552
rect 328604 334512 329012 334540
rect 328604 334500 328610 334512
rect 329006 334500 329012 334512
rect 329064 334500 329070 334552
rect 250165 334475 250223 334481
rect 250165 334441 250177 334475
rect 250211 334472 250223 334475
rect 250622 334472 250628 334484
rect 250211 334444 250628 334472
rect 250211 334441 250223 334444
rect 250165 334435 250223 334441
rect 250622 334432 250628 334444
rect 250680 334432 250686 334484
rect 270770 334296 270776 334348
rect 270828 334336 270834 334348
rect 271230 334336 271236 334348
rect 270828 334308 271236 334336
rect 270828 334296 270834 334308
rect 271230 334296 271236 334308
rect 271288 334296 271294 334348
rect 272242 334296 272248 334348
rect 272300 334336 272306 334348
rect 272702 334336 272708 334348
rect 272300 334308 272708 334336
rect 272300 334296 272306 334308
rect 272702 334296 272708 334308
rect 272760 334296 272766 334348
rect 247126 334160 247132 334212
rect 247184 334200 247190 334212
rect 248138 334200 248144 334212
rect 247184 334172 248144 334200
rect 247184 334160 247190 334172
rect 248138 334160 248144 334172
rect 248196 334160 248202 334212
rect 335354 334160 335360 334212
rect 335412 334200 335418 334212
rect 335998 334200 336004 334212
rect 335412 334172 336004 334200
rect 335412 334160 335418 334172
rect 335998 334160 336004 334172
rect 336056 334160 336062 334212
rect 304994 333752 305000 333804
rect 305052 333792 305058 333804
rect 305638 333792 305644 333804
rect 305052 333764 305644 333792
rect 305052 333752 305058 333764
rect 305638 333752 305644 333764
rect 305696 333752 305702 333804
rect 301038 333276 301044 333328
rect 301096 333316 301102 333328
rect 301682 333316 301688 333328
rect 301096 333288 301688 333316
rect 301096 333276 301102 333288
rect 301682 333276 301688 333288
rect 301740 333276 301746 333328
rect 325878 333276 325884 333328
rect 325936 333316 325942 333328
rect 326614 333316 326620 333328
rect 325936 333288 326620 333316
rect 325936 333276 325942 333288
rect 326614 333276 326620 333288
rect 326672 333276 326678 333328
rect 361666 333276 361672 333328
rect 361724 333316 361730 333328
rect 362310 333316 362316 333328
rect 361724 333288 362316 333316
rect 361724 333276 361730 333288
rect 362310 333276 362316 333288
rect 362368 333276 362374 333328
rect 306466 333072 306472 333124
rect 306524 333112 306530 333124
rect 306650 333112 306656 333124
rect 306524 333084 306656 333112
rect 306524 333072 306530 333084
rect 306650 333072 306656 333084
rect 306708 333072 306714 333124
rect 262582 333004 262588 333056
rect 262640 333044 262646 333056
rect 263042 333044 263048 333056
rect 262640 333016 263048 333044
rect 262640 333004 262646 333016
rect 263042 333004 263048 333016
rect 263100 333004 263106 333056
rect 284662 332528 284668 332580
rect 284720 332568 284726 332580
rect 285122 332568 285128 332580
rect 284720 332540 285128 332568
rect 284720 332528 284726 332540
rect 285122 332528 285128 332540
rect 285180 332528 285186 332580
rect 242986 332052 242992 332104
rect 243044 332092 243050 332104
rect 243446 332092 243452 332104
rect 243044 332064 243452 332092
rect 243044 332052 243050 332064
rect 243446 332052 243452 332064
rect 243504 332052 243510 332104
rect 336734 331984 336740 332036
rect 336792 332024 336798 332036
rect 336918 332024 336924 332036
rect 336792 331996 336924 332024
rect 336792 331984 336798 331996
rect 336918 331984 336924 331996
rect 336976 331984 336982 332036
rect 284294 331916 284300 331968
rect 284352 331956 284358 331968
rect 284570 331956 284576 331968
rect 284352 331928 284576 331956
rect 284352 331916 284358 331928
rect 284570 331916 284576 331928
rect 284628 331916 284634 331968
rect 357342 331848 357348 331900
rect 357400 331888 357406 331900
rect 357986 331888 357992 331900
rect 357400 331860 357992 331888
rect 357400 331848 357406 331860
rect 357986 331848 357992 331860
rect 358044 331848 358050 331900
rect 299566 331304 299572 331356
rect 299624 331304 299630 331356
rect 336826 331304 336832 331356
rect 336884 331304 336890 331356
rect 259638 331168 259644 331220
rect 259696 331208 259702 331220
rect 259822 331208 259828 331220
rect 259696 331180 259828 331208
rect 259696 331168 259702 331180
rect 259822 331168 259828 331180
rect 259880 331168 259886 331220
rect 262582 331168 262588 331220
rect 262640 331208 262646 331220
rect 262766 331208 262772 331220
rect 262640 331180 262772 331208
rect 262640 331168 262646 331180
rect 262766 331168 262772 331180
rect 262824 331168 262830 331220
rect 299584 331084 299612 331304
rect 336844 331220 336872 331304
rect 389726 331236 389732 331288
rect 389784 331236 389790 331288
rect 336826 331168 336832 331220
rect 336884 331168 336890 331220
rect 389634 331168 389640 331220
rect 389692 331208 389698 331220
rect 389744 331208 389772 331236
rect 389692 331180 389772 331208
rect 389692 331168 389698 331180
rect 299566 331032 299572 331084
rect 299624 331032 299630 331084
rect 299474 330964 299480 331016
rect 299532 331004 299538 331016
rect 299842 331004 299848 331016
rect 299532 330976 299848 331004
rect 299532 330964 299538 330976
rect 299842 330964 299848 330976
rect 299900 330964 299906 331016
rect 321462 329128 321468 329180
rect 321520 329168 321526 329180
rect 321833 329171 321891 329177
rect 321833 329168 321845 329171
rect 321520 329140 321845 329168
rect 321520 329128 321526 329140
rect 321833 329137 321845 329140
rect 321879 329137 321891 329171
rect 321833 329131 321891 329137
rect 347498 328556 347504 328568
rect 338868 328528 347504 328556
rect 338868 328500 338896 328528
rect 347498 328516 347504 328528
rect 347556 328516 347562 328568
rect 250162 328488 250168 328500
rect 250123 328460 250168 328488
rect 250162 328448 250168 328460
rect 250220 328448 250226 328500
rect 278866 328448 278872 328500
rect 278924 328488 278930 328500
rect 279050 328488 279056 328500
rect 278924 328460 279056 328488
rect 278924 328448 278930 328460
rect 279050 328448 279056 328460
rect 279108 328448 279114 328500
rect 288802 328448 288808 328500
rect 288860 328488 288866 328500
rect 289078 328488 289084 328500
rect 288860 328460 289084 328488
rect 288860 328448 288866 328460
rect 289078 328448 289084 328460
rect 289136 328448 289142 328500
rect 302510 328488 302516 328500
rect 302471 328460 302516 328488
rect 302510 328448 302516 328460
rect 302568 328448 302574 328500
rect 303890 328448 303896 328500
rect 303948 328488 303954 328500
rect 304626 328488 304632 328500
rect 303948 328460 304632 328488
rect 303948 328448 303954 328460
rect 304626 328448 304632 328460
rect 304684 328448 304690 328500
rect 323302 328448 323308 328500
rect 323360 328488 323366 328500
rect 323670 328488 323676 328500
rect 323360 328460 323676 328488
rect 323360 328448 323366 328460
rect 323670 328448 323676 328460
rect 323728 328448 323734 328500
rect 324682 328448 324688 328500
rect 324740 328488 324746 328500
rect 325050 328488 325056 328500
rect 324740 328460 325056 328488
rect 324740 328448 324746 328460
rect 325050 328448 325056 328460
rect 325108 328448 325114 328500
rect 338850 328448 338856 328500
rect 338908 328448 338914 328500
rect 339770 328448 339776 328500
rect 339828 328488 339834 328500
rect 340322 328488 340328 328500
rect 339828 328460 340328 328488
rect 339828 328448 339834 328460
rect 340322 328448 340328 328460
rect 340380 328448 340386 328500
rect 341426 328448 341432 328500
rect 341484 328488 341490 328500
rect 341705 328491 341763 328497
rect 341705 328488 341717 328491
rect 341484 328460 341717 328488
rect 341484 328448 341490 328460
rect 341705 328457 341717 328460
rect 341751 328457 341763 328491
rect 341705 328451 341763 328457
rect 372706 328448 372712 328500
rect 372764 328488 372770 328500
rect 373258 328488 373264 328500
rect 372764 328460 373264 328488
rect 372764 328448 372770 328460
rect 373258 328448 373264 328460
rect 373316 328448 373322 328500
rect 259822 328420 259828 328432
rect 259783 328392 259828 328420
rect 259822 328380 259828 328392
rect 259880 328380 259886 328432
rect 295518 328380 295524 328432
rect 295576 328420 295582 328432
rect 295702 328420 295708 328432
rect 295576 328392 295708 328420
rect 295576 328380 295582 328392
rect 295702 328380 295708 328392
rect 295760 328380 295766 328432
rect 296806 328380 296812 328432
rect 296864 328420 296870 328432
rect 296990 328420 296996 328432
rect 296864 328392 296996 328420
rect 296864 328380 296870 328392
rect 296990 328380 296996 328392
rect 297048 328380 297054 328432
rect 389545 328423 389603 328429
rect 389545 328389 389557 328423
rect 389591 328420 389603 328423
rect 389634 328420 389640 328432
rect 389591 328392 389640 328420
rect 389591 328389 389603 328392
rect 389545 328383 389603 328389
rect 389634 328380 389640 328392
rect 389692 328380 389698 328432
rect 470594 328420 470600 328432
rect 470555 328392 470600 328420
rect 470594 328380 470600 328392
rect 470652 328380 470658 328432
rect 330202 327196 330208 327208
rect 330163 327168 330208 327196
rect 330202 327156 330208 327168
rect 330260 327156 330266 327208
rect 327258 327088 327264 327140
rect 327316 327128 327322 327140
rect 327442 327128 327448 327140
rect 327316 327100 327448 327128
rect 327316 327088 327322 327100
rect 327442 327088 327448 327100
rect 327500 327088 327506 327140
rect 331398 327128 331404 327140
rect 331359 327100 331404 327128
rect 331398 327088 331404 327100
rect 331456 327088 331462 327140
rect 374454 327128 374460 327140
rect 374415 327100 374460 327128
rect 374454 327088 374460 327100
rect 374512 327088 374518 327140
rect 375837 327131 375895 327137
rect 375837 327097 375849 327131
rect 375883 327128 375895 327131
rect 375926 327128 375932 327140
rect 375883 327100 375932 327128
rect 375883 327097 375895 327100
rect 375837 327091 375895 327097
rect 375926 327088 375932 327100
rect 375984 327088 375990 327140
rect 302510 327020 302516 327072
rect 302568 327060 302574 327072
rect 302602 327060 302608 327072
rect 302568 327032 302608 327060
rect 302568 327020 302574 327032
rect 302602 327020 302608 327032
rect 302660 327020 302666 327072
rect 357434 327060 357440 327072
rect 357395 327032 357440 327060
rect 357434 327020 357440 327032
rect 357492 327020 357498 327072
rect 360381 327063 360439 327069
rect 360381 327029 360393 327063
rect 360427 327060 360439 327063
rect 360470 327060 360476 327072
rect 360427 327032 360476 327060
rect 360427 327029 360439 327032
rect 360381 327023 360439 327029
rect 360470 327020 360476 327032
rect 360528 327020 360534 327072
rect 463694 325660 463700 325712
rect 463752 325700 463758 325712
rect 463878 325700 463884 325712
rect 463752 325672 463884 325700
rect 463752 325660 463758 325672
rect 463878 325660 463884 325672
rect 463936 325660 463942 325712
rect 580074 325660 580080 325712
rect 580132 325700 580138 325712
rect 580902 325700 580908 325712
rect 580132 325672 580908 325700
rect 580132 325660 580138 325672
rect 580902 325660 580908 325672
rect 580960 325660 580966 325712
rect 3326 324232 3332 324284
rect 3384 324272 3390 324284
rect 14458 324272 14464 324284
rect 3384 324244 14464 324272
rect 3384 324232 3390 324244
rect 14458 324232 14464 324244
rect 14516 324232 14522 324284
rect 376846 323552 376852 323604
rect 376904 323592 376910 323604
rect 377122 323592 377128 323604
rect 376904 323564 377128 323592
rect 376904 323552 376910 323564
rect 377122 323552 377128 323564
rect 377180 323552 377186 323604
rect 470042 322872 470048 322924
rect 470100 322912 470106 322924
rect 580074 322912 580080 322924
rect 470100 322884 580080 322912
rect 470100 322872 470106 322884
rect 580074 322872 580080 322884
rect 580132 322872 580138 322924
rect 239122 321648 239128 321700
rect 239180 321648 239186 321700
rect 235074 321580 235080 321632
rect 235132 321580 235138 321632
rect 230750 321512 230756 321564
rect 230808 321552 230814 321564
rect 230934 321552 230940 321564
rect 230808 321524 230940 321552
rect 230808 321512 230814 321524
rect 230934 321512 230940 321524
rect 230992 321512 230998 321564
rect 232222 321512 232228 321564
rect 232280 321552 232286 321564
rect 232406 321552 232412 321564
rect 232280 321524 232412 321552
rect 232280 321512 232286 321524
rect 232406 321512 232412 321524
rect 232464 321512 232470 321564
rect 235092 321496 235120 321580
rect 239140 321564 239168 321648
rect 251450 321580 251456 321632
rect 251508 321580 251514 321632
rect 286042 321620 286048 321632
rect 285968 321592 286048 321620
rect 239122 321512 239128 321564
rect 239180 321512 239186 321564
rect 235074 321444 235080 321496
rect 235132 321444 235138 321496
rect 251468 321416 251496 321580
rect 285968 321564 285996 321592
rect 286042 321580 286048 321592
rect 286100 321580 286106 321632
rect 310790 321580 310796 321632
rect 310848 321580 310854 321632
rect 337194 321620 337200 321632
rect 337155 321592 337200 321620
rect 337194 321580 337200 321592
rect 337252 321580 337258 321632
rect 341426 321620 341432 321632
rect 341387 321592 341432 321620
rect 341426 321580 341432 321592
rect 341484 321580 341490 321632
rect 285950 321512 285956 321564
rect 286008 321512 286014 321564
rect 310808 321484 310836 321580
rect 310882 321484 310888 321496
rect 310808 321456 310888 321484
rect 310882 321444 310888 321456
rect 310940 321444 310946 321496
rect 251542 321416 251548 321428
rect 251468 321388 251548 321416
rect 251542 321376 251548 321388
rect 251600 321376 251606 321428
rect 337194 320872 337200 320884
rect 337155 320844 337200 320872
rect 337194 320832 337200 320844
rect 337252 320832 337258 320884
rect 259825 318835 259883 318841
rect 259825 318801 259837 318835
rect 259871 318832 259883 318835
rect 259914 318832 259920 318844
rect 259871 318804 259920 318832
rect 259871 318801 259883 318804
rect 259825 318795 259883 318801
rect 259914 318792 259920 318804
rect 259972 318792 259978 318844
rect 294230 318792 294236 318844
rect 294288 318832 294294 318844
rect 294322 318832 294328 318844
rect 294288 318804 294328 318832
rect 294288 318792 294294 318804
rect 294322 318792 294328 318804
rect 294380 318792 294386 318844
rect 306742 318792 306748 318844
rect 306800 318832 306806 318844
rect 306834 318832 306840 318844
rect 306800 318804 306840 318832
rect 306800 318792 306806 318804
rect 306834 318792 306840 318804
rect 306892 318792 306898 318844
rect 341426 318832 341432 318844
rect 341387 318804 341432 318832
rect 341426 318792 341432 318804
rect 341484 318792 341490 318844
rect 374362 318792 374368 318844
rect 374420 318832 374426 318844
rect 374454 318832 374460 318844
rect 374420 318804 374460 318832
rect 374420 318792 374426 318804
rect 374454 318792 374460 318804
rect 374512 318792 374518 318844
rect 375834 318792 375840 318844
rect 375892 318832 375898 318844
rect 375926 318832 375932 318844
rect 375892 318804 375932 318832
rect 375892 318792 375898 318804
rect 375926 318792 375932 318804
rect 375984 318792 375990 318844
rect 389542 318832 389548 318844
rect 389503 318804 389548 318832
rect 389542 318792 389548 318804
rect 389600 318792 389606 318844
rect 470594 318832 470600 318844
rect 470555 318804 470600 318832
rect 470594 318792 470600 318804
rect 470652 318792 470658 318844
rect 230845 318767 230903 318773
rect 230845 318733 230857 318767
rect 230891 318764 230903 318767
rect 230934 318764 230940 318776
rect 230891 318736 230940 318764
rect 230891 318733 230903 318736
rect 230845 318727 230903 318733
rect 230934 318724 230940 318736
rect 230992 318724 230998 318776
rect 236270 318764 236276 318776
rect 236231 318736 236276 318764
rect 236270 318724 236276 318736
rect 236328 318724 236334 318776
rect 239214 318764 239220 318776
rect 239175 318736 239220 318764
rect 239214 318724 239220 318736
rect 239272 318724 239278 318776
rect 284665 318767 284723 318773
rect 284665 318733 284677 318767
rect 284711 318764 284723 318767
rect 284754 318764 284760 318776
rect 284711 318736 284760 318764
rect 284711 318733 284723 318736
rect 284665 318727 284723 318733
rect 284754 318724 284760 318736
rect 284812 318724 284818 318776
rect 285950 318724 285956 318776
rect 286008 318764 286014 318776
rect 286134 318764 286140 318776
rect 286008 318736 286140 318764
rect 286008 318724 286014 318736
rect 286134 318724 286140 318736
rect 286192 318724 286198 318776
rect 357437 317475 357495 317481
rect 357437 317441 357449 317475
rect 357483 317472 357495 317475
rect 357526 317472 357532 317484
rect 357483 317444 357532 317472
rect 357483 317441 357495 317444
rect 357437 317435 357495 317441
rect 357526 317432 357532 317444
rect 357584 317432 357590 317484
rect 360378 317472 360384 317484
rect 360339 317444 360384 317472
rect 360378 317432 360384 317444
rect 360436 317432 360442 317484
rect 291562 317364 291568 317416
rect 291620 317364 291626 317416
rect 299753 317407 299811 317413
rect 299753 317373 299765 317407
rect 299799 317404 299811 317407
rect 299842 317404 299848 317416
rect 299799 317376 299848 317404
rect 299799 317373 299811 317376
rect 299753 317367 299811 317373
rect 299842 317364 299848 317376
rect 299900 317364 299906 317416
rect 325881 317407 325939 317413
rect 325881 317373 325893 317407
rect 325927 317404 325939 317407
rect 325970 317404 325976 317416
rect 325927 317376 325976 317404
rect 325927 317373 325939 317376
rect 325881 317367 325939 317373
rect 325970 317364 325976 317376
rect 326028 317364 326034 317416
rect 337194 317404 337200 317416
rect 337155 317376 337200 317404
rect 337194 317364 337200 317376
rect 337252 317364 337258 317416
rect 375834 317404 375840 317416
rect 375795 317376 375840 317404
rect 375834 317364 375840 317376
rect 375892 317364 375898 317416
rect 377122 317364 377128 317416
rect 377180 317404 377186 317416
rect 377306 317404 377312 317416
rect 377180 317376 377312 317404
rect 377180 317364 377186 317376
rect 377306 317364 377312 317376
rect 377364 317364 377370 317416
rect 291580 317336 291608 317364
rect 291654 317336 291660 317348
rect 291580 317308 291660 317336
rect 291654 317296 291660 317308
rect 291712 317296 291718 317348
rect 579982 316072 579988 316124
rect 580040 316112 580046 316124
rect 580994 316112 581000 316124
rect 580040 316084 581000 316112
rect 580040 316072 580046 316084
rect 580994 316072 581000 316084
rect 581052 316072 581058 316124
rect 262585 315979 262643 315985
rect 262585 315945 262597 315979
rect 262631 315976 262643 315979
rect 262674 315976 262680 315988
rect 262631 315948 262680 315976
rect 262631 315945 262643 315948
rect 262585 315939 262643 315945
rect 262674 315936 262680 315948
rect 262732 315936 262738 315988
rect 580074 315936 580080 315988
rect 580132 315976 580138 315988
rect 580994 315976 581000 315988
rect 580132 315948 581000 315976
rect 580132 315936 580138 315948
rect 580994 315936 581000 315948
rect 581052 315936 581058 315988
rect 284665 314211 284723 314217
rect 284665 314177 284677 314211
rect 284711 314208 284723 314211
rect 284938 314208 284944 314220
rect 284711 314180 284944 314208
rect 284711 314177 284723 314180
rect 284665 314171 284723 314177
rect 284938 314168 284944 314180
rect 284996 314168 285002 314220
rect 250162 313964 250168 314016
rect 250220 313964 250226 314016
rect 250180 313880 250208 313964
rect 288618 313896 288624 313948
rect 288676 313936 288682 313948
rect 288802 313936 288808 313948
rect 288676 313908 288808 313936
rect 288676 313896 288682 313908
rect 288802 313896 288808 313908
rect 288860 313896 288866 313948
rect 250162 313828 250168 313880
rect 250220 313828 250226 313880
rect 273441 313463 273499 313469
rect 273441 313429 273453 313463
rect 273487 313460 273499 313463
rect 273622 313460 273628 313472
rect 273487 313432 273628 313460
rect 273487 313429 273499 313432
rect 273441 313423 273499 313429
rect 273622 313420 273628 313432
rect 273680 313420 273686 313472
rect 272242 311924 272248 311976
rect 272300 311924 272306 311976
rect 306834 311964 306840 311976
rect 306760 311936 306840 311964
rect 259730 311856 259736 311908
rect 259788 311896 259794 311908
rect 259914 311896 259920 311908
rect 259788 311868 259920 311896
rect 259788 311856 259794 311868
rect 259914 311856 259920 311868
rect 259972 311856 259978 311908
rect 272260 311840 272288 311924
rect 273438 311896 273444 311908
rect 273399 311868 273444 311896
rect 273438 311856 273444 311868
rect 273496 311856 273502 311908
rect 306760 311840 306788 311936
rect 306834 311924 306840 311936
rect 306892 311924 306898 311976
rect 310882 311964 310888 311976
rect 310843 311936 310888 311964
rect 310882 311924 310888 311936
rect 310940 311924 310946 311976
rect 323302 311964 323308 311976
rect 323228 311936 323308 311964
rect 323228 311908 323256 311936
rect 323302 311924 323308 311936
rect 323360 311924 323366 311976
rect 374362 311924 374368 311976
rect 374420 311924 374426 311976
rect 323210 311856 323216 311908
rect 323268 311856 323274 311908
rect 341242 311856 341248 311908
rect 341300 311896 341306 311908
rect 341426 311896 341432 311908
rect 341300 311868 341432 311896
rect 341300 311856 341306 311868
rect 341426 311856 341432 311868
rect 341484 311856 341490 311908
rect 244458 311828 244464 311840
rect 244419 311800 244464 311828
rect 244458 311788 244464 311800
rect 244516 311788 244522 311840
rect 272242 311788 272248 311840
rect 272300 311788 272306 311840
rect 306742 311788 306748 311840
rect 306800 311788 306806 311840
rect 337194 311760 337200 311772
rect 337155 311732 337200 311760
rect 337194 311720 337200 311732
rect 337252 311720 337258 311772
rect 374380 311760 374408 311924
rect 374454 311760 374460 311772
rect 374380 311732 374460 311760
rect 374454 311720 374460 311732
rect 374512 311720 374518 311772
rect 236270 309244 236276 309256
rect 236231 309216 236276 309244
rect 236270 309204 236276 309216
rect 236328 309204 236334 309256
rect 295610 309244 295616 309256
rect 295536 309216 295616 309244
rect 230842 309176 230848 309188
rect 230803 309148 230848 309176
rect 230842 309136 230848 309148
rect 230900 309136 230906 309188
rect 239214 309176 239220 309188
rect 239175 309148 239220 309176
rect 239214 309136 239220 309148
rect 239272 309136 239278 309188
rect 244458 309176 244464 309188
rect 244419 309148 244464 309176
rect 244458 309136 244464 309148
rect 244516 309136 244522 309188
rect 267734 309136 267740 309188
rect 267792 309176 267798 309188
rect 267826 309176 267832 309188
rect 267792 309148 267832 309176
rect 267792 309136 267798 309148
rect 267826 309136 267832 309148
rect 267884 309136 267890 309188
rect 295536 309120 295564 309216
rect 295610 309204 295616 309216
rect 295668 309204 295674 309256
rect 296898 309244 296904 309256
rect 296824 309216 296904 309244
rect 296824 309120 296852 309216
rect 296898 309204 296904 309216
rect 296956 309204 296962 309256
rect 389358 309136 389364 309188
rect 389416 309176 389422 309188
rect 389542 309176 389548 309188
rect 389416 309148 389548 309176
rect 389416 309136 389422 309148
rect 389542 309136 389548 309148
rect 389600 309136 389606 309188
rect 236270 309108 236276 309120
rect 236231 309080 236276 309108
rect 236270 309068 236276 309080
rect 236328 309068 236334 309120
rect 259641 309111 259699 309117
rect 259641 309077 259653 309111
rect 259687 309108 259699 309111
rect 259730 309108 259736 309120
rect 259687 309080 259736 309108
rect 259687 309077 259699 309080
rect 259641 309071 259699 309077
rect 259730 309068 259736 309080
rect 259788 309068 259794 309120
rect 295518 309068 295524 309120
rect 295576 309068 295582 309120
rect 296806 309068 296812 309120
rect 296864 309068 296870 309120
rect 327166 309068 327172 309120
rect 327224 309108 327230 309120
rect 327258 309108 327264 309120
rect 327224 309080 327264 309108
rect 327224 309068 327230 309080
rect 327258 309068 327264 309080
rect 327316 309068 327322 309120
rect 341153 309111 341211 309117
rect 341153 309077 341165 309111
rect 341199 309108 341211 309111
rect 341242 309108 341248 309120
rect 341199 309080 341248 309108
rect 341199 309077 341211 309080
rect 341153 309071 341211 309077
rect 341242 309068 341248 309080
rect 341300 309068 341306 309120
rect 357802 309108 357808 309120
rect 357763 309080 357808 309108
rect 357802 309068 357808 309080
rect 357860 309068 357866 309120
rect 358722 309108 358728 309120
rect 358683 309080 358728 309108
rect 358722 309068 358728 309080
rect 358780 309068 358786 309120
rect 470594 309108 470600 309120
rect 470555 309080 470600 309108
rect 470594 309068 470600 309080
rect 470652 309068 470658 309120
rect 389269 309043 389327 309049
rect 389269 309009 389281 309043
rect 389315 309040 389327 309043
rect 389358 309040 389364 309052
rect 389315 309012 389364 309040
rect 389315 309009 389327 309012
rect 389269 309003 389327 309009
rect 389358 309000 389364 309012
rect 389416 309000 389422 309052
rect 2774 308796 2780 308848
rect 2832 308836 2838 308848
rect 5442 308836 5448 308848
rect 2832 308808 5448 308836
rect 2832 308796 2838 308808
rect 5442 308796 5448 308808
rect 5500 308796 5506 308848
rect 310698 307844 310704 307896
rect 310756 307884 310762 307896
rect 310885 307887 310943 307893
rect 310885 307884 310897 307887
rect 310756 307856 310897 307884
rect 310756 307844 310762 307856
rect 310885 307853 310897 307856
rect 310931 307853 310943 307887
rect 310885 307847 310943 307853
rect 325878 307816 325884 307828
rect 325839 307788 325884 307816
rect 325878 307776 325884 307788
rect 325936 307776 325942 307828
rect 375834 307816 375840 307828
rect 375795 307788 375840 307816
rect 375834 307776 375840 307788
rect 375892 307776 375898 307828
rect 310698 307748 310704 307760
rect 310659 307720 310704 307748
rect 310698 307708 310704 307720
rect 310756 307708 310762 307760
rect 327166 307748 327172 307760
rect 327127 307720 327172 307748
rect 327166 307708 327172 307720
rect 327224 307708 327230 307760
rect 337194 307748 337200 307760
rect 337155 307720 337200 307748
rect 337194 307708 337200 307720
rect 337252 307708 337258 307760
rect 374365 307751 374423 307757
rect 374365 307717 374377 307751
rect 374411 307748 374423 307751
rect 374454 307748 374460 307760
rect 374411 307720 374460 307748
rect 374411 307717 374423 307720
rect 374365 307711 374423 307717
rect 374454 307708 374460 307720
rect 374512 307708 374518 307760
rect 301038 306348 301044 306400
rect 301096 306388 301102 306400
rect 301222 306388 301228 306400
rect 301096 306360 301228 306388
rect 301096 306348 301102 306360
rect 301222 306348 301228 306360
rect 301280 306348 301286 306400
rect 317506 306348 317512 306400
rect 317564 306388 317570 306400
rect 317690 306388 317696 306400
rect 317564 306360 317696 306388
rect 317564 306348 317570 306360
rect 317690 306348 317696 306360
rect 317748 306348 317754 306400
rect 463694 306348 463700 306400
rect 463752 306388 463758 306400
rect 463878 306388 463884 306400
rect 463752 306360 463884 306388
rect 463752 306348 463758 306360
rect 463878 306348 463884 306360
rect 463936 306348 463942 306400
rect 580074 306348 580080 306400
rect 580132 306388 580138 306400
rect 580902 306388 580908 306400
rect 580132 306360 580908 306388
rect 580132 306348 580138 306360
rect 580902 306348 580908 306360
rect 580960 306348 580966 306400
rect 294230 304240 294236 304292
rect 294288 304280 294294 304292
rect 294414 304280 294420 304292
rect 294288 304252 294420 304280
rect 294288 304240 294294 304252
rect 294414 304240 294420 304252
rect 294472 304240 294478 304292
rect 338850 302200 338856 302252
rect 338908 302200 338914 302252
rect 338868 302104 338896 302200
rect 338942 302104 338948 302116
rect 338868 302076 338948 302104
rect 338942 302064 338948 302076
rect 339000 302064 339006 302116
rect 377122 302064 377128 302116
rect 377180 302104 377186 302116
rect 377306 302104 377312 302116
rect 377180 302076 377312 302104
rect 377180 302064 377186 302076
rect 377306 302064 377312 302076
rect 377364 302064 377370 302116
rect 236270 299588 236276 299600
rect 236231 299560 236276 299588
rect 236270 299548 236276 299560
rect 236328 299548 236334 299600
rect 259638 299588 259644 299600
rect 259599 299560 259644 299588
rect 259638 299548 259644 299560
rect 259696 299548 259702 299600
rect 267826 299588 267832 299600
rect 267752 299560 267832 299588
rect 267752 299464 267780 299560
rect 267826 299548 267832 299560
rect 267884 299548 267890 299600
rect 288618 299480 288624 299532
rect 288676 299520 288682 299532
rect 288802 299520 288808 299532
rect 288676 299492 288808 299520
rect 288676 299480 288682 299492
rect 288802 299480 288808 299492
rect 288860 299480 288866 299532
rect 299753 299523 299811 299529
rect 299753 299489 299765 299523
rect 299799 299520 299811 299523
rect 299842 299520 299848 299532
rect 299799 299492 299848 299520
rect 299799 299489 299811 299492
rect 299753 299483 299811 299489
rect 299842 299480 299848 299492
rect 299900 299480 299906 299532
rect 306742 299480 306748 299532
rect 306800 299520 306806 299532
rect 306834 299520 306840 299532
rect 306800 299492 306840 299520
rect 306800 299480 306806 299492
rect 306834 299480 306840 299492
rect 306892 299480 306898 299532
rect 341150 299520 341156 299532
rect 341111 299492 341156 299520
rect 341150 299480 341156 299492
rect 341208 299480 341214 299532
rect 357805 299523 357863 299529
rect 357805 299489 357817 299523
rect 357851 299520 357863 299523
rect 357894 299520 357900 299532
rect 357851 299492 357900 299520
rect 357851 299489 357863 299492
rect 357805 299483 357863 299489
rect 357894 299480 357900 299492
rect 357952 299480 357958 299532
rect 358722 299520 358728 299532
rect 358683 299492 358728 299520
rect 358722 299480 358728 299492
rect 358780 299480 358786 299532
rect 389266 299520 389272 299532
rect 389227 299492 389272 299520
rect 389266 299480 389272 299492
rect 389324 299480 389330 299532
rect 470594 299520 470600 299532
rect 470555 299492 470600 299520
rect 470594 299480 470600 299492
rect 470652 299480 470658 299532
rect 235074 299412 235080 299464
rect 235132 299452 235138 299464
rect 235166 299452 235172 299464
rect 235132 299424 235172 299452
rect 235132 299412 235138 299424
rect 235166 299412 235172 299424
rect 235224 299412 235230 299464
rect 236270 299452 236276 299464
rect 236231 299424 236276 299452
rect 236270 299412 236276 299424
rect 236328 299412 236334 299464
rect 259638 299412 259644 299464
rect 259696 299452 259702 299464
rect 259822 299452 259828 299464
rect 259696 299424 259828 299452
rect 259696 299412 259702 299424
rect 259822 299412 259828 299424
rect 259880 299412 259886 299464
rect 267734 299412 267740 299464
rect 267792 299412 267798 299464
rect 323302 299452 323308 299464
rect 323263 299424 323308 299452
rect 323302 299412 323308 299424
rect 323360 299412 323366 299464
rect 324682 299452 324688 299464
rect 324643 299424 324688 299452
rect 324682 299412 324688 299424
rect 324740 299412 324746 299464
rect 325878 299412 325884 299464
rect 325936 299412 325942 299464
rect 338942 299452 338948 299464
rect 338868 299424 338948 299452
rect 325896 299384 325924 299412
rect 338868 299396 338896 299424
rect 338942 299412 338948 299424
rect 339000 299412 339006 299464
rect 372706 299452 372712 299464
rect 372667 299424 372712 299452
rect 372706 299412 372712 299424
rect 372764 299412 372770 299464
rect 375837 299455 375895 299461
rect 375837 299421 375849 299455
rect 375883 299452 375895 299455
rect 375926 299452 375932 299464
rect 375883 299424 375932 299452
rect 375883 299421 375895 299424
rect 375837 299415 375895 299421
rect 375926 299412 375932 299424
rect 375984 299412 375990 299464
rect 469950 299412 469956 299464
rect 470008 299452 470014 299464
rect 580166 299452 580172 299464
rect 470008 299424 580172 299452
rect 470008 299412 470014 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 325970 299384 325976 299396
rect 325896 299356 325976 299384
rect 325970 299344 325976 299356
rect 326028 299344 326034 299396
rect 338850 299344 338856 299396
rect 338908 299344 338914 299396
rect 262582 298228 262588 298240
rect 262543 298200 262588 298228
rect 262582 298188 262588 298200
rect 262640 298188 262646 298240
rect 310701 298163 310759 298169
rect 310701 298129 310713 298163
rect 310747 298160 310759 298163
rect 310882 298160 310888 298172
rect 310747 298132 310888 298160
rect 310747 298129 310759 298132
rect 310701 298123 310759 298129
rect 310882 298120 310888 298132
rect 310940 298120 310946 298172
rect 327169 298163 327227 298169
rect 327169 298129 327181 298163
rect 327215 298160 327227 298163
rect 327258 298160 327264 298172
rect 327215 298132 327264 298160
rect 327215 298129 327227 298132
rect 327169 298123 327227 298129
rect 327258 298120 327264 298132
rect 327316 298120 327322 298172
rect 330110 298120 330116 298172
rect 330168 298160 330174 298172
rect 330202 298160 330208 298172
rect 330168 298132 330208 298160
rect 330168 298120 330174 298132
rect 330202 298120 330208 298132
rect 330260 298120 330266 298172
rect 337197 298163 337255 298169
rect 337197 298129 337209 298163
rect 337243 298160 337255 298163
rect 337286 298160 337292 298172
rect 337243 298132 337292 298160
rect 337243 298129 337255 298132
rect 337197 298123 337255 298129
rect 337286 298120 337292 298132
rect 337344 298120 337350 298172
rect 262582 298052 262588 298104
rect 262640 298052 262646 298104
rect 266722 298092 266728 298104
rect 266683 298064 266728 298092
rect 266722 298052 266728 298064
rect 266780 298052 266786 298104
rect 267734 298092 267740 298104
rect 267695 298064 267740 298092
rect 267734 298052 267740 298064
rect 267792 298052 267798 298104
rect 285950 298092 285956 298104
rect 285911 298064 285956 298092
rect 285950 298052 285956 298064
rect 286008 298052 286014 298104
rect 325970 298052 325976 298104
rect 326028 298092 326034 298104
rect 326062 298092 326068 298104
rect 326028 298064 326068 298092
rect 326028 298052 326034 298064
rect 326062 298052 326068 298064
rect 326120 298052 326126 298104
rect 358722 298092 358728 298104
rect 358683 298064 358728 298092
rect 358722 298052 358728 298064
rect 358780 298052 358786 298104
rect 262600 297968 262628 298052
rect 262582 297916 262588 297968
rect 262640 297916 262646 297968
rect 301038 296760 301044 296812
rect 301096 296800 301102 296812
rect 301406 296800 301412 296812
rect 301096 296772 301412 296800
rect 301096 296760 301102 296772
rect 301406 296760 301412 296772
rect 301464 296760 301470 296812
rect 580074 296760 580080 296812
rect 580132 296800 580138 296812
rect 580994 296800 581000 296812
rect 580132 296772 581000 296800
rect 580132 296760 580138 296772
rect 580994 296760 581000 296772
rect 581052 296760 581058 296812
rect 284754 296692 284760 296744
rect 284812 296732 284818 296744
rect 284846 296732 284852 296744
rect 284812 296704 284852 296732
rect 284812 296692 284818 296704
rect 284846 296692 284852 296704
rect 284904 296692 284910 296744
rect 299842 296624 299848 296676
rect 299900 296664 299906 296676
rect 299934 296664 299940 296676
rect 299900 296636 299940 296664
rect 299900 296624 299906 296636
rect 299934 296624 299940 296636
rect 299992 296624 299998 296676
rect 301038 296624 301044 296676
rect 301096 296664 301102 296676
rect 301130 296664 301136 296676
rect 301096 296636 301136 296664
rect 301096 296624 301102 296636
rect 301130 296624 301136 296636
rect 301188 296624 301194 296676
rect 306834 296624 306840 296676
rect 306892 296664 306898 296676
rect 306926 296664 306932 296676
rect 306892 296636 306932 296664
rect 306892 296624 306898 296636
rect 306926 296624 306932 296636
rect 306984 296624 306990 296676
rect 580166 296624 580172 296676
rect 580224 296664 580230 296676
rect 580994 296664 581000 296676
rect 580224 296636 581000 296664
rect 580224 296624 580230 296636
rect 580994 296624 581000 296636
rect 581052 296624 581058 296676
rect 272334 295440 272340 295452
rect 272260 295412 272340 295440
rect 272260 295316 272288 295412
rect 272334 295400 272340 295412
rect 272392 295400 272398 295452
rect 272242 295264 272248 295316
rect 272300 295264 272306 295316
rect 302510 295264 302516 295316
rect 302568 295304 302574 295316
rect 302694 295304 302700 295316
rect 302568 295276 302700 295304
rect 302568 295264 302574 295276
rect 302694 295264 302700 295276
rect 302752 295264 302758 295316
rect 251453 294695 251511 294701
rect 251453 294661 251465 294695
rect 251499 294692 251511 294695
rect 251542 294692 251548 294704
rect 251499 294664 251548 294692
rect 251499 294661 251511 294664
rect 251453 294655 251511 294661
rect 251542 294652 251548 294664
rect 251600 294652 251606 294704
rect 289998 294584 290004 294636
rect 290056 294624 290062 294636
rect 290182 294624 290188 294636
rect 290056 294596 290188 294624
rect 290056 294584 290062 294596
rect 290182 294584 290188 294596
rect 290240 294584 290246 294636
rect 310882 293060 310888 293072
rect 310843 293032 310888 293060
rect 310882 293020 310888 293032
rect 310940 293020 310946 293072
rect 377122 292612 377128 292664
rect 377180 292612 377186 292664
rect 239214 292584 239220 292596
rect 239175 292556 239220 292584
rect 239214 292544 239220 292556
rect 239272 292544 239278 292596
rect 288710 292544 288716 292596
rect 288768 292584 288774 292596
rect 288768 292556 288848 292584
rect 288768 292544 288774 292556
rect 288820 292528 288848 292556
rect 295518 292544 295524 292596
rect 295576 292544 295582 292596
rect 296806 292544 296812 292596
rect 296864 292544 296870 292596
rect 337102 292544 337108 292596
rect 337160 292584 337166 292596
rect 337286 292584 337292 292596
rect 337160 292556 337292 292584
rect 337160 292544 337166 292556
rect 337286 292544 337292 292556
rect 337344 292544 337350 292596
rect 357434 292544 357440 292596
rect 357492 292584 357498 292596
rect 357894 292584 357900 292596
rect 357492 292556 357900 292584
rect 357492 292544 357498 292556
rect 357894 292544 357900 292556
rect 357952 292544 357958 292596
rect 270770 292516 270776 292528
rect 270731 292488 270776 292516
rect 270770 292476 270776 292488
rect 270828 292476 270834 292528
rect 288802 292476 288808 292528
rect 288860 292476 288866 292528
rect 295536 292516 295564 292544
rect 295610 292516 295616 292528
rect 295536 292488 295616 292516
rect 295610 292476 295616 292488
rect 295668 292476 295674 292528
rect 296824 292516 296852 292544
rect 296898 292516 296904 292528
rect 296824 292488 296904 292516
rect 296898 292476 296904 292488
rect 296956 292476 296962 292528
rect 377140 292460 377168 292612
rect 377122 292408 377128 292460
rect 377180 292408 377186 292460
rect 236270 289864 236276 289876
rect 236231 289836 236276 289864
rect 236270 289824 236276 289836
rect 236328 289824 236334 289876
rect 239214 289864 239220 289876
rect 239175 289836 239220 289864
rect 239214 289824 239220 289836
rect 239272 289824 239278 289876
rect 251450 289864 251456 289876
rect 251411 289836 251456 289864
rect 251450 289824 251456 289836
rect 251508 289824 251514 289876
rect 294233 289867 294291 289873
rect 294233 289833 294245 289867
rect 294279 289864 294291 289867
rect 294322 289864 294328 289876
rect 294279 289836 294328 289864
rect 294279 289833 294291 289836
rect 294233 289827 294291 289833
rect 294322 289824 294328 289836
rect 294380 289824 294386 289876
rect 324682 289864 324688 289876
rect 324643 289836 324688 289864
rect 324682 289824 324688 289836
rect 324740 289824 324746 289876
rect 372706 289864 372712 289876
rect 372667 289836 372712 289864
rect 372706 289824 372712 289836
rect 372764 289824 372770 289876
rect 374362 289864 374368 289876
rect 374323 289836 374368 289864
rect 374362 289824 374368 289836
rect 374420 289824 374426 289876
rect 375834 289864 375840 289876
rect 375795 289836 375840 289864
rect 375834 289824 375840 289836
rect 375892 289824 375898 289876
rect 244458 289796 244464 289808
rect 244419 289768 244464 289796
rect 244458 289756 244464 289768
rect 244516 289756 244522 289808
rect 250070 289756 250076 289808
rect 250128 289796 250134 289808
rect 250346 289796 250352 289808
rect 250128 289768 250352 289796
rect 250128 289756 250134 289768
rect 250346 289756 250352 289768
rect 250404 289756 250410 289808
rect 259730 289756 259736 289808
rect 259788 289796 259794 289808
rect 259914 289796 259920 289808
rect 259788 289768 259920 289796
rect 259788 289756 259794 289768
rect 259914 289756 259920 289768
rect 259972 289756 259978 289808
rect 289998 289756 290004 289808
rect 290056 289796 290062 289808
rect 290182 289796 290188 289808
rect 290056 289768 290188 289796
rect 290056 289756 290062 289768
rect 290182 289756 290188 289768
rect 290240 289756 290246 289808
rect 327169 289799 327227 289805
rect 327169 289765 327181 289799
rect 327215 289796 327227 289799
rect 327258 289796 327264 289808
rect 327215 289768 327264 289796
rect 327215 289765 327227 289768
rect 327169 289759 327227 289765
rect 327258 289756 327264 289768
rect 327316 289756 327322 289808
rect 357434 289756 357440 289808
rect 357492 289796 357498 289808
rect 389361 289799 389419 289805
rect 357492 289768 357537 289796
rect 357492 289756 357498 289768
rect 389361 289765 389373 289799
rect 389407 289796 389419 289799
rect 389450 289796 389456 289808
rect 389407 289768 389456 289796
rect 389407 289765 389419 289768
rect 389361 289759 389419 289765
rect 389450 289756 389456 289768
rect 389508 289756 389514 289808
rect 470594 289796 470600 289808
rect 470555 289768 470600 289796
rect 470594 289756 470600 289768
rect 470652 289756 470658 289808
rect 236270 289728 236276 289740
rect 236231 289700 236276 289728
rect 236270 289688 236276 289700
rect 236328 289688 236334 289740
rect 266722 288436 266728 288448
rect 266683 288408 266728 288436
rect 266722 288396 266728 288408
rect 266780 288396 266786 288448
rect 267734 288436 267740 288448
rect 267695 288408 267740 288436
rect 267734 288396 267740 288408
rect 267792 288396 267798 288448
rect 285950 288436 285956 288448
rect 285911 288408 285956 288436
rect 285950 288396 285956 288408
rect 286008 288396 286014 288448
rect 323302 288436 323308 288448
rect 323263 288408 323308 288436
rect 323302 288396 323308 288408
rect 323360 288396 323366 288448
rect 358722 288436 358728 288448
rect 358683 288408 358728 288436
rect 358722 288396 358728 288408
rect 358780 288396 358786 288448
rect 291562 287036 291568 287088
rect 291620 287076 291626 287088
rect 291654 287076 291660 287088
rect 291620 287048 291660 287076
rect 291620 287036 291626 287048
rect 291654 287036 291660 287048
rect 291712 287036 291718 287088
rect 294230 287076 294236 287088
rect 294191 287048 294236 287076
rect 294230 287036 294236 287048
rect 294288 287036 294294 287088
rect 330478 287036 330484 287088
rect 330536 287076 330542 287088
rect 330662 287076 330668 287088
rect 330536 287048 330668 287076
rect 330536 287036 330542 287048
rect 330662 287036 330668 287048
rect 330720 287036 330726 287088
rect 463694 287036 463700 287088
rect 463752 287076 463758 287088
rect 463878 287076 463884 287088
rect 463752 287048 463884 287076
rect 463752 287036 463758 287048
rect 463878 287036 463884 287048
rect 463936 287036 463942 287088
rect 580166 287036 580172 287088
rect 580224 287076 580230 287088
rect 580902 287076 580908 287088
rect 580224 287048 580908 287076
rect 580224 287036 580230 287048
rect 580902 287036 580908 287048
rect 580960 287036 580966 287088
rect 270770 285648 270776 285660
rect 270731 285620 270776 285648
rect 270770 285608 270776 285620
rect 270828 285608 270834 285660
rect 337197 285651 337255 285657
rect 337197 285617 337209 285651
rect 337243 285648 337255 285651
rect 337286 285648 337292 285660
rect 337243 285620 337292 285648
rect 337243 285617 337255 285620
rect 337197 285611 337255 285617
rect 337286 285608 337292 285620
rect 337344 285608 337350 285660
rect 284386 283568 284392 283620
rect 284444 283608 284450 283620
rect 284846 283608 284852 283620
rect 284444 283580 284852 283608
rect 284444 283568 284450 283580
rect 284846 283568 284852 283580
rect 284904 283568 284910 283620
rect 323394 283568 323400 283620
rect 323452 283608 323458 283620
rect 323489 283611 323547 283617
rect 323489 283608 323501 283611
rect 323452 283580 323501 283608
rect 323452 283568 323458 283580
rect 323489 283577 323501 283580
rect 323535 283577 323547 283611
rect 323489 283571 323547 283577
rect 327169 283611 327227 283617
rect 327169 283577 327181 283611
rect 327215 283608 327227 283611
rect 327258 283608 327264 283620
rect 327215 283580 327264 283608
rect 327215 283577 327227 283580
rect 327169 283571 327227 283577
rect 327258 283568 327264 283580
rect 327316 283568 327322 283620
rect 296898 282996 296904 283008
rect 296824 282968 296904 282996
rect 296824 282872 296852 282968
rect 296898 282956 296904 282968
rect 296956 282956 296962 283008
rect 341150 282928 341156 282940
rect 341111 282900 341156 282928
rect 341150 282888 341156 282900
rect 341208 282888 341214 282940
rect 360286 282888 360292 282940
rect 360344 282928 360350 282940
rect 360470 282928 360476 282940
rect 360344 282900 360476 282928
rect 360344 282888 360350 282900
rect 360470 282888 360476 282900
rect 360528 282888 360534 282940
rect 296806 282820 296812 282872
rect 296864 282820 296870 282872
rect 310882 282792 310888 282804
rect 310843 282764 310888 282792
rect 310882 282752 310888 282764
rect 310940 282752 310946 282804
rect 358722 280304 358728 280356
rect 358780 280304 358786 280356
rect 236270 280276 236276 280288
rect 236231 280248 236276 280276
rect 236270 280236 236276 280248
rect 236328 280236 236334 280288
rect 358740 280220 358768 280304
rect 244458 280208 244464 280220
rect 244419 280180 244464 280208
rect 244458 280168 244464 280180
rect 244516 280168 244522 280220
rect 265250 280168 265256 280220
rect 265308 280168 265314 280220
rect 295518 280168 295524 280220
rect 295576 280208 295582 280220
rect 295610 280208 295616 280220
rect 295576 280180 295616 280208
rect 295576 280168 295582 280180
rect 295610 280168 295616 280180
rect 295668 280168 295674 280220
rect 341150 280208 341156 280220
rect 341111 280180 341156 280208
rect 341150 280168 341156 280180
rect 341208 280168 341214 280220
rect 357437 280211 357495 280217
rect 357437 280177 357449 280211
rect 357483 280208 357495 280211
rect 357710 280208 357716 280220
rect 357483 280180 357716 280208
rect 357483 280177 357495 280180
rect 357437 280171 357495 280177
rect 357710 280168 357716 280180
rect 357768 280168 357774 280220
rect 358722 280168 358728 280220
rect 358780 280168 358786 280220
rect 389358 280208 389364 280220
rect 389319 280180 389364 280208
rect 389358 280168 389364 280180
rect 389416 280168 389422 280220
rect 470594 280208 470600 280220
rect 470555 280180 470600 280208
rect 470594 280168 470600 280180
rect 470652 280168 470658 280220
rect 235074 280100 235080 280152
rect 235132 280140 235138 280152
rect 235166 280140 235172 280152
rect 235132 280112 235172 280140
rect 235132 280100 235138 280112
rect 235166 280100 235172 280112
rect 235224 280100 235230 280152
rect 236270 280140 236276 280152
rect 236231 280112 236276 280140
rect 236270 280100 236276 280112
rect 236328 280100 236334 280152
rect 239122 280140 239128 280152
rect 239083 280112 239128 280140
rect 239122 280100 239128 280112
rect 239180 280100 239186 280152
rect 251450 280140 251456 280152
rect 251411 280112 251456 280140
rect 251450 280100 251456 280112
rect 251508 280100 251514 280152
rect 259546 280140 259552 280152
rect 259507 280112 259552 280140
rect 259546 280100 259552 280112
rect 259604 280100 259610 280152
rect 265268 280084 265296 280168
rect 273530 280100 273536 280152
rect 273588 280140 273594 280152
rect 273622 280140 273628 280152
rect 273588 280112 273628 280140
rect 273588 280100 273594 280112
rect 273622 280100 273628 280112
rect 273680 280100 273686 280152
rect 285950 280100 285956 280152
rect 286008 280140 286014 280152
rect 286134 280140 286140 280152
rect 286008 280112 286140 280140
rect 286008 280100 286014 280112
rect 286134 280100 286140 280112
rect 286192 280100 286198 280152
rect 288618 280100 288624 280152
rect 288676 280140 288682 280152
rect 288802 280140 288808 280152
rect 288676 280112 288808 280140
rect 288676 280100 288682 280112
rect 288802 280100 288808 280112
rect 288860 280100 288866 280152
rect 331398 280140 331404 280152
rect 331359 280112 331404 280140
rect 331398 280100 331404 280112
rect 331456 280100 331462 280152
rect 338850 280140 338856 280152
rect 338811 280112 338856 280140
rect 338850 280100 338856 280112
rect 338908 280100 338914 280152
rect 372706 280140 372712 280152
rect 372667 280112 372712 280140
rect 372706 280100 372712 280112
rect 372764 280100 372770 280152
rect 377122 280140 377128 280152
rect 377083 280112 377128 280140
rect 377122 280100 377128 280112
rect 377180 280100 377186 280152
rect 265250 280032 265256 280084
rect 265308 280032 265314 280084
rect 291562 278808 291568 278860
rect 291620 278848 291626 278860
rect 291746 278848 291752 278860
rect 291620 278820 291752 278848
rect 291620 278808 291626 278820
rect 291746 278808 291752 278820
rect 291804 278808 291810 278860
rect 250070 278740 250076 278792
rect 250128 278780 250134 278792
rect 250162 278780 250168 278792
rect 250128 278752 250168 278780
rect 250128 278740 250134 278752
rect 250162 278740 250168 278752
rect 250220 278740 250226 278792
rect 301038 278740 301044 278792
rect 301096 278780 301102 278792
rect 301222 278780 301228 278792
rect 301096 278752 301228 278780
rect 301096 278740 301102 278752
rect 301222 278740 301228 278752
rect 301280 278740 301286 278792
rect 302510 278740 302516 278792
rect 302568 278740 302574 278792
rect 323486 278780 323492 278792
rect 323447 278752 323492 278780
rect 323486 278740 323492 278752
rect 323544 278740 323550 278792
rect 330202 278740 330208 278792
rect 330260 278780 330266 278792
rect 330478 278780 330484 278792
rect 330260 278752 330484 278780
rect 330260 278740 330266 278752
rect 330478 278740 330484 278752
rect 330536 278740 330542 278792
rect 302528 278712 302556 278740
rect 302602 278712 302608 278724
rect 302528 278684 302608 278712
rect 302602 278672 302608 278684
rect 302660 278672 302666 278724
rect 310882 278712 310888 278724
rect 310843 278684 310888 278712
rect 310882 278672 310888 278684
rect 310940 278672 310946 278724
rect 294230 277380 294236 277432
rect 294288 277420 294294 277432
rect 294322 277420 294328 277432
rect 294288 277392 294328 277420
rect 294288 277380 294294 277392
rect 294322 277380 294328 277392
rect 294380 277380 294386 277432
rect 580166 277312 580172 277364
rect 580224 277352 580230 277364
rect 580902 277352 580908 277364
rect 580224 277324 580908 277352
rect 580224 277312 580230 277324
rect 580902 277312 580908 277324
rect 580960 277312 580966 277364
rect 337194 276060 337200 276072
rect 337155 276032 337200 276060
rect 337194 276020 337200 276032
rect 337252 276020 337258 276072
rect 302602 275952 302608 276004
rect 302660 275992 302666 276004
rect 302786 275992 302792 276004
rect 302660 275964 302792 275992
rect 302660 275952 302666 275964
rect 302786 275952 302792 275964
rect 302844 275952 302850 276004
rect 306650 275952 306656 276004
rect 306708 275992 306714 276004
rect 306926 275992 306932 276004
rect 306708 275964 306932 275992
rect 306708 275952 306714 275964
rect 306926 275952 306932 275964
rect 306984 275952 306990 276004
rect 284386 273912 284392 273964
rect 284444 273952 284450 273964
rect 284754 273952 284760 273964
rect 284444 273924 284760 273952
rect 284444 273912 284450 273924
rect 284754 273912 284760 273924
rect 284812 273912 284818 273964
rect 330110 273884 330116 273896
rect 330071 273856 330116 273884
rect 330110 273844 330116 273856
rect 330168 273844 330174 273896
rect 250162 273340 250168 273352
rect 250088 273312 250168 273340
rect 250088 273216 250116 273312
rect 250162 273300 250168 273312
rect 250220 273300 250226 273352
rect 301038 273232 301044 273284
rect 301096 273232 301102 273284
rect 357434 273232 357440 273284
rect 357492 273272 357498 273284
rect 357710 273272 357716 273284
rect 357492 273244 357716 273272
rect 357492 273232 357498 273244
rect 357710 273232 357716 273244
rect 357768 273232 357774 273284
rect 250070 273164 250076 273216
rect 250128 273164 250134 273216
rect 301056 273204 301084 273232
rect 301130 273204 301136 273216
rect 301056 273176 301136 273204
rect 301130 273164 301136 273176
rect 301188 273164 301194 273216
rect 374362 273164 374368 273216
rect 374420 273164 374426 273216
rect 375834 273164 375840 273216
rect 375892 273164 375898 273216
rect 374380 273080 374408 273164
rect 375852 273080 375880 273164
rect 259546 273068 259552 273080
rect 259507 273040 259552 273068
rect 259546 273028 259552 273040
rect 259604 273028 259610 273080
rect 374362 273028 374368 273080
rect 374420 273028 374426 273080
rect 375834 273028 375840 273080
rect 375892 273028 375898 273080
rect 299934 270620 299940 270632
rect 299768 270592 299940 270620
rect 299768 270564 299796 270592
rect 299934 270580 299940 270592
rect 299992 270580 299998 270632
rect 236270 270552 236276 270564
rect 236231 270524 236276 270552
rect 236270 270512 236276 270524
rect 236328 270512 236334 270564
rect 239125 270555 239183 270561
rect 239125 270521 239137 270555
rect 239171 270552 239183 270555
rect 239214 270552 239220 270564
rect 239171 270524 239220 270552
rect 239171 270521 239183 270524
rect 239125 270515 239183 270521
rect 239214 270512 239220 270524
rect 239272 270512 239278 270564
rect 251450 270552 251456 270564
rect 251411 270524 251456 270552
rect 251450 270512 251456 270524
rect 251508 270512 251514 270564
rect 262490 270512 262496 270564
rect 262548 270552 262554 270564
rect 262674 270552 262680 270564
rect 262548 270524 262680 270552
rect 262548 270512 262554 270524
rect 262674 270512 262680 270524
rect 262732 270512 262738 270564
rect 267734 270512 267740 270564
rect 267792 270552 267798 270564
rect 267826 270552 267832 270564
rect 267792 270524 267832 270552
rect 267792 270512 267798 270524
rect 267826 270512 267832 270524
rect 267884 270512 267890 270564
rect 299750 270512 299756 270564
rect 299808 270512 299814 270564
rect 331398 270552 331404 270564
rect 331359 270524 331404 270552
rect 331398 270512 331404 270524
rect 331456 270512 331462 270564
rect 338850 270552 338856 270564
rect 338811 270524 338856 270552
rect 338850 270512 338856 270524
rect 338908 270512 338914 270564
rect 372706 270552 372712 270564
rect 372667 270524 372712 270552
rect 372706 270512 372712 270524
rect 372764 270512 372770 270564
rect 377122 270552 377128 270564
rect 377083 270524 377128 270552
rect 377122 270512 377128 270524
rect 377180 270512 377186 270564
rect 325970 270444 325976 270496
rect 326028 270484 326034 270496
rect 326062 270484 326068 270496
rect 326028 270456 326068 270484
rect 326028 270444 326034 270456
rect 326062 270444 326068 270456
rect 326120 270444 326126 270496
rect 341242 270444 341248 270496
rect 341300 270484 341306 270496
rect 341426 270484 341432 270496
rect 341300 270456 341432 270484
rect 341300 270444 341306 270456
rect 341426 270444 341432 270456
rect 341484 270444 341490 270496
rect 389361 270487 389419 270493
rect 389361 270453 389373 270487
rect 389407 270484 389419 270487
rect 389450 270484 389456 270496
rect 389407 270456 389456 270484
rect 389407 270453 389419 270456
rect 389361 270447 389419 270453
rect 389450 270444 389456 270456
rect 389508 270444 389514 270496
rect 470594 270484 470600 270496
rect 470555 270456 470600 270484
rect 470594 270444 470600 270456
rect 470652 270444 470658 270496
rect 236270 270416 236276 270428
rect 236231 270388 236276 270416
rect 236270 270376 236276 270388
rect 236328 270376 236334 270428
rect 291746 269192 291752 269204
rect 291580 269164 291752 269192
rect 290090 269084 290096 269136
rect 290148 269124 290154 269136
rect 290182 269124 290188 269136
rect 290148 269096 290188 269124
rect 290148 269084 290154 269096
rect 290182 269084 290188 269096
rect 290240 269084 290246 269136
rect 291580 269068 291608 269164
rect 291746 269152 291752 269164
rect 291804 269152 291810 269204
rect 296806 269084 296812 269136
rect 296864 269124 296870 269136
rect 297082 269124 297088 269136
rect 296864 269096 297088 269124
rect 296864 269084 296870 269096
rect 297082 269084 297088 269096
rect 297140 269084 297146 269136
rect 324590 269084 324596 269136
rect 324648 269124 324654 269136
rect 324774 269124 324780 269136
rect 324648 269096 324780 269124
rect 324648 269084 324654 269096
rect 324774 269084 324780 269096
rect 324832 269084 324838 269136
rect 330113 269127 330171 269133
rect 330113 269093 330125 269127
rect 330159 269124 330171 269127
rect 330202 269124 330208 269136
rect 330159 269096 330208 269124
rect 330159 269093 330171 269096
rect 330113 269087 330171 269093
rect 330202 269084 330208 269096
rect 330260 269084 330266 269136
rect 358538 269084 358544 269136
rect 358596 269124 358602 269136
rect 358722 269124 358728 269136
rect 358596 269096 358728 269124
rect 358596 269084 358602 269096
rect 358722 269084 358728 269096
rect 358780 269084 358786 269136
rect 250070 269056 250076 269068
rect 250031 269028 250076 269056
rect 250070 269016 250076 269028
rect 250128 269016 250134 269068
rect 291562 269016 291568 269068
rect 291620 269016 291626 269068
rect 265250 267724 265256 267776
rect 265308 267764 265314 267776
rect 265434 267764 265440 267776
rect 265308 267736 265440 267764
rect 265308 267724 265314 267736
rect 265434 267724 265440 267736
rect 265492 267724 265498 267776
rect 294138 267724 294144 267776
rect 294196 267764 294202 267776
rect 294322 267764 294328 267776
rect 294196 267736 294328 267764
rect 294196 267724 294202 267736
rect 294322 267724 294328 267736
rect 294380 267724 294386 267776
rect 295518 267724 295524 267776
rect 295576 267764 295582 267776
rect 295794 267764 295800 267776
rect 295576 267736 295800 267764
rect 295576 267724 295582 267736
rect 295794 267724 295800 267736
rect 295852 267724 295858 267776
rect 463694 267724 463700 267776
rect 463752 267764 463758 267776
rect 463878 267764 463884 267776
rect 463752 267736 463884 267764
rect 463752 267724 463758 267736
rect 463878 267724 463884 267736
rect 463936 267724 463942 267776
rect 337010 266296 337016 266348
rect 337068 266336 337074 266348
rect 337194 266336 337200 266348
rect 337068 266308 337200 266336
rect 337068 266296 337074 266308
rect 337194 266296 337200 266308
rect 337252 266296 337258 266348
rect 327258 263684 327264 263696
rect 327184 263656 327264 263684
rect 270678 263576 270684 263628
rect 270736 263576 270742 263628
rect 270696 263492 270724 263576
rect 327184 263560 327212 263656
rect 327258 263644 327264 263656
rect 327316 263644 327322 263696
rect 360286 263576 360292 263628
rect 360344 263616 360350 263628
rect 360470 263616 360476 263628
rect 360344 263588 360476 263616
rect 360344 263576 360350 263588
rect 360470 263576 360476 263588
rect 360528 263576 360534 263628
rect 327166 263508 327172 263560
rect 327224 263508 327230 263560
rect 270678 263440 270684 263492
rect 270736 263440 270742 263492
rect 310882 263480 310888 263492
rect 310843 263452 310888 263480
rect 310882 263440 310888 263452
rect 310940 263440 310946 263492
rect 296806 262896 296812 262948
rect 296864 262936 296870 262948
rect 296990 262936 296996 262948
rect 296864 262908 296996 262936
rect 296864 262896 296870 262908
rect 296990 262896 296996 262908
rect 297048 262896 297054 262948
rect 236270 260964 236276 260976
rect 236231 260936 236276 260964
rect 236270 260924 236276 260936
rect 236328 260924 236334 260976
rect 323394 260924 323400 260976
rect 323452 260964 323458 260976
rect 323486 260964 323492 260976
rect 323452 260936 323492 260964
rect 323452 260924 323458 260936
rect 323486 260924 323492 260936
rect 323544 260924 323550 260976
rect 262582 260896 262588 260908
rect 262543 260868 262588 260896
rect 262582 260856 262588 260868
rect 262640 260856 262646 260908
rect 266630 260856 266636 260908
rect 266688 260896 266694 260908
rect 266722 260896 266728 260908
rect 266688 260868 266728 260896
rect 266688 260856 266694 260868
rect 266722 260856 266728 260868
rect 266780 260856 266786 260908
rect 288618 260856 288624 260908
rect 288676 260896 288682 260908
rect 288802 260896 288808 260908
rect 288676 260868 288808 260896
rect 288676 260856 288682 260868
rect 288802 260856 288808 260868
rect 288860 260856 288866 260908
rect 295702 260856 295708 260908
rect 295760 260896 295766 260908
rect 389358 260896 389364 260908
rect 295760 260868 295840 260896
rect 389319 260868 389364 260896
rect 295760 260856 295766 260868
rect 295812 260840 295840 260868
rect 389358 260856 389364 260868
rect 389416 260856 389422 260908
rect 470594 260896 470600 260908
rect 470555 260868 470600 260896
rect 470594 260856 470600 260868
rect 470652 260856 470658 260908
rect 235074 260788 235080 260840
rect 235132 260828 235138 260840
rect 235166 260828 235172 260840
rect 235132 260800 235172 260828
rect 235132 260788 235138 260800
rect 235166 260788 235172 260800
rect 235224 260788 235230 260840
rect 236270 260828 236276 260840
rect 236231 260800 236276 260828
rect 236270 260788 236276 260800
rect 236328 260788 236334 260840
rect 239122 260828 239128 260840
rect 239083 260800 239128 260828
rect 239122 260788 239128 260800
rect 239180 260788 239186 260840
rect 251450 260828 251456 260840
rect 251411 260800 251456 260828
rect 251450 260788 251456 260800
rect 251508 260788 251514 260840
rect 259546 260828 259552 260840
rect 259507 260800 259552 260828
rect 259546 260788 259552 260800
rect 259604 260788 259610 260840
rect 270678 260828 270684 260840
rect 270639 260800 270684 260828
rect 270678 260788 270684 260800
rect 270736 260788 270742 260840
rect 272150 260788 272156 260840
rect 272208 260788 272214 260840
rect 273530 260788 273536 260840
rect 273588 260828 273594 260840
rect 273622 260828 273628 260840
rect 273588 260800 273628 260828
rect 273588 260788 273594 260800
rect 273622 260788 273628 260800
rect 273680 260788 273686 260840
rect 295794 260788 295800 260840
rect 295852 260788 295858 260840
rect 324590 260788 324596 260840
rect 324648 260788 324654 260840
rect 338850 260828 338856 260840
rect 338811 260800 338856 260828
rect 338850 260788 338856 260800
rect 338908 260788 338914 260840
rect 341058 260828 341064 260840
rect 341019 260800 341064 260828
rect 341058 260788 341064 260800
rect 341116 260788 341122 260840
rect 372706 260828 372712 260840
rect 372667 260800 372712 260828
rect 372706 260788 372712 260800
rect 372764 260788 372770 260840
rect 377122 260828 377128 260840
rect 377083 260800 377128 260828
rect 377122 260788 377128 260800
rect 377180 260788 377186 260840
rect 463697 260831 463755 260837
rect 463697 260797 463709 260831
rect 463743 260828 463755 260831
rect 463786 260828 463792 260840
rect 463743 260800 463792 260828
rect 463743 260797 463755 260800
rect 463697 260791 463755 260797
rect 463786 260788 463792 260800
rect 463844 260788 463850 260840
rect 272168 260704 272196 260788
rect 324608 260760 324636 260788
rect 324682 260760 324688 260772
rect 324608 260732 324688 260760
rect 324682 260720 324688 260732
rect 324740 260720 324746 260772
rect 272150 260652 272156 260704
rect 272208 260652 272214 260704
rect 250073 259471 250131 259477
rect 250073 259437 250085 259471
rect 250119 259468 250131 259471
rect 250162 259468 250168 259480
rect 250119 259440 250168 259468
rect 250119 259437 250131 259440
rect 250073 259431 250131 259437
rect 250162 259428 250168 259440
rect 250220 259428 250226 259480
rect 262582 259468 262588 259480
rect 262543 259440 262588 259468
rect 262582 259428 262588 259440
rect 262640 259428 262646 259480
rect 267734 259428 267740 259480
rect 267792 259468 267798 259480
rect 267826 259468 267832 259480
rect 267792 259440 267832 259468
rect 267792 259428 267798 259440
rect 267826 259428 267832 259440
rect 267884 259428 267890 259480
rect 284570 259428 284576 259480
rect 284628 259468 284634 259480
rect 284754 259468 284760 259480
rect 284628 259440 284760 259468
rect 284628 259428 284634 259440
rect 284754 259428 284760 259440
rect 284812 259428 284818 259480
rect 330110 259428 330116 259480
rect 330168 259468 330174 259480
rect 330386 259468 330392 259480
rect 330168 259440 330392 259468
rect 330168 259428 330174 259440
rect 330386 259428 330392 259440
rect 330444 259428 330450 259480
rect 324682 259360 324688 259412
rect 324740 259400 324746 259412
rect 324774 259400 324780 259412
rect 324740 259372 324780 259400
rect 324740 259360 324746 259372
rect 324774 259360 324780 259372
rect 324832 259360 324838 259412
rect 357526 259400 357532 259412
rect 357487 259372 357532 259400
rect 357526 259360 357532 259372
rect 357584 259360 357590 259412
rect 250162 259332 250168 259344
rect 250123 259304 250168 259332
rect 250162 259292 250168 259304
rect 250220 259292 250226 259344
rect 264974 258000 264980 258052
rect 265032 258040 265038 258052
rect 265342 258040 265348 258052
rect 265032 258012 265348 258040
rect 265032 258000 265038 258012
rect 265342 258000 265348 258012
rect 265400 258000 265406 258052
rect 267918 258000 267924 258052
rect 267976 258040 267982 258052
rect 268102 258040 268108 258052
rect 267976 258012 268108 258040
rect 267976 258000 267982 258012
rect 268102 258000 268108 258012
rect 268160 258000 268166 258052
rect 301222 258000 301228 258052
rect 301280 258040 301286 258052
rect 301406 258040 301412 258052
rect 301280 258012 301412 258040
rect 301280 258000 301286 258012
rect 301406 258000 301412 258012
rect 301464 258000 301470 258052
rect 306745 258043 306803 258049
rect 306745 258009 306757 258043
rect 306791 258040 306803 258043
rect 306834 258040 306840 258052
rect 306791 258012 306840 258040
rect 306791 258009 306803 258012
rect 306745 258003 306803 258009
rect 306834 258000 306840 258012
rect 306892 258000 306898 258052
rect 330110 258000 330116 258052
rect 330168 258040 330174 258052
rect 330294 258040 330300 258052
rect 330168 258012 330300 258040
rect 330168 258000 330174 258012
rect 330294 258000 330300 258012
rect 330352 258000 330358 258052
rect 310882 256068 310888 256080
rect 310843 256040 310888 256068
rect 310882 256028 310888 256040
rect 310940 256028 310946 256080
rect 337105 254031 337163 254037
rect 337105 253997 337117 254031
rect 337151 254028 337163 254031
rect 337194 254028 337200 254040
rect 337151 254000 337200 254028
rect 337151 253997 337163 254000
rect 337105 253991 337163 253997
rect 337194 253988 337200 254000
rect 337252 253988 337258 254040
rect 374362 253852 374368 253904
rect 374420 253852 374426 253904
rect 375834 253852 375840 253904
rect 375892 253852 375898 253904
rect 374380 253768 374408 253852
rect 375852 253768 375880 253852
rect 259546 253756 259552 253768
rect 259507 253728 259552 253756
rect 259546 253716 259552 253728
rect 259604 253716 259610 253768
rect 341058 253756 341064 253768
rect 341019 253728 341064 253756
rect 341058 253716 341064 253728
rect 341116 253716 341122 253768
rect 374362 253716 374368 253768
rect 374420 253716 374426 253768
rect 375834 253716 375840 253768
rect 375892 253716 375898 253768
rect 295242 253172 295248 253224
rect 295300 253212 295306 253224
rect 295610 253212 295616 253224
rect 295300 253184 295616 253212
rect 295300 253172 295306 253184
rect 295610 253172 295616 253184
rect 295668 253172 295674 253224
rect 469858 252492 469864 252544
rect 469916 252532 469922 252544
rect 579614 252532 579620 252544
rect 469916 252504 579620 252532
rect 469916 252492 469922 252504
rect 579614 252492 579620 252504
rect 579672 252492 579678 252544
rect 2774 252016 2780 252068
rect 2832 252056 2838 252068
rect 5350 252056 5356 252068
rect 2832 252028 5356 252056
rect 2832 252016 2838 252028
rect 5350 252016 5356 252028
rect 5408 252016 5414 252068
rect 310698 251268 310704 251320
rect 310756 251308 310762 251320
rect 310885 251311 310943 251317
rect 310885 251308 310897 251311
rect 310756 251280 310897 251308
rect 310756 251268 310762 251280
rect 310885 251277 310897 251280
rect 310931 251277 310943 251311
rect 310885 251271 310943 251277
rect 236270 251240 236276 251252
rect 236231 251212 236276 251240
rect 236270 251200 236276 251212
rect 236328 251200 236334 251252
rect 239125 251243 239183 251249
rect 239125 251209 239137 251243
rect 239171 251240 239183 251243
rect 239214 251240 239220 251252
rect 239171 251212 239220 251240
rect 239171 251209 239183 251212
rect 239125 251203 239183 251209
rect 239214 251200 239220 251212
rect 239272 251200 239278 251252
rect 251450 251240 251456 251252
rect 251411 251212 251456 251240
rect 251450 251200 251456 251212
rect 251508 251200 251514 251252
rect 289998 251200 290004 251252
rect 290056 251240 290062 251252
rect 290090 251240 290096 251252
rect 290056 251212 290096 251240
rect 290056 251200 290062 251212
rect 290090 251200 290096 251212
rect 290148 251200 290154 251252
rect 327166 251200 327172 251252
rect 327224 251240 327230 251252
rect 327258 251240 327264 251252
rect 327224 251212 327264 251240
rect 327224 251200 327230 251212
rect 327258 251200 327264 251212
rect 327316 251200 327322 251252
rect 338850 251240 338856 251252
rect 338811 251212 338856 251240
rect 338850 251200 338856 251212
rect 338908 251200 338914 251252
rect 372706 251240 372712 251252
rect 372667 251212 372712 251240
rect 372706 251200 372712 251212
rect 372764 251200 372770 251252
rect 377122 251240 377128 251252
rect 377083 251212 377128 251240
rect 377122 251200 377128 251212
rect 377180 251200 377186 251252
rect 389174 251200 389180 251252
rect 389232 251240 389238 251252
rect 389358 251240 389364 251252
rect 389232 251212 389364 251240
rect 389232 251200 389238 251212
rect 389358 251200 389364 251212
rect 389416 251200 389422 251252
rect 463694 251200 463700 251252
rect 463752 251240 463758 251252
rect 463752 251212 463797 251240
rect 463752 251200 463758 251212
rect 259546 251172 259552 251184
rect 259507 251144 259552 251172
rect 259546 251132 259552 251144
rect 259604 251132 259610 251184
rect 310698 251172 310704 251184
rect 310659 251144 310704 251172
rect 310698 251132 310704 251144
rect 310756 251132 310762 251184
rect 325970 251132 325976 251184
rect 326028 251172 326034 251184
rect 326062 251172 326068 251184
rect 326028 251144 326068 251172
rect 326028 251132 326034 251144
rect 326062 251132 326068 251144
rect 326120 251132 326126 251184
rect 470594 251172 470600 251184
rect 470555 251144 470600 251172
rect 470594 251132 470600 251144
rect 470652 251132 470658 251184
rect 250165 251107 250223 251113
rect 250165 251073 250177 251107
rect 250211 251104 250223 251107
rect 250346 251104 250352 251116
rect 250211 251076 250352 251104
rect 250211 251073 250223 251076
rect 250165 251067 250223 251073
rect 250346 251064 250352 251076
rect 250404 251064 250410 251116
rect 270681 251107 270739 251113
rect 270681 251073 270693 251107
rect 270727 251104 270739 251107
rect 270770 251104 270776 251116
rect 270727 251076 270776 251104
rect 270727 251073 270739 251076
rect 270681 251067 270739 251073
rect 270770 251064 270776 251076
rect 270828 251064 270834 251116
rect 284662 249840 284668 249892
rect 284720 249880 284726 249892
rect 284754 249880 284760 249892
rect 284720 249852 284760 249880
rect 284720 249840 284726 249852
rect 284754 249840 284760 249852
rect 284812 249840 284818 249892
rect 285950 249772 285956 249824
rect 286008 249812 286014 249824
rect 286042 249812 286048 249824
rect 286008 249784 286048 249812
rect 286008 249772 286014 249784
rect 286042 249772 286048 249784
rect 286100 249772 286106 249824
rect 302694 249772 302700 249824
rect 302752 249812 302758 249824
rect 302786 249812 302792 249824
rect 302752 249784 302792 249812
rect 302752 249772 302758 249784
rect 302786 249772 302792 249784
rect 302844 249772 302850 249824
rect 323210 249772 323216 249824
rect 323268 249812 323274 249824
rect 323486 249812 323492 249824
rect 323268 249784 323492 249812
rect 323268 249772 323274 249784
rect 323486 249772 323492 249784
rect 323544 249772 323550 249824
rect 357529 249815 357587 249821
rect 357529 249781 357541 249815
rect 357575 249812 357587 249815
rect 357710 249812 357716 249824
rect 357575 249784 357716 249812
rect 357575 249781 357587 249784
rect 357529 249775 357587 249781
rect 357710 249772 357716 249784
rect 357768 249772 357774 249824
rect 358538 249772 358544 249824
rect 358596 249812 358602 249824
rect 358722 249812 358728 249824
rect 358596 249784 358728 249812
rect 358596 249772 358602 249784
rect 358722 249772 358728 249784
rect 358780 249772 358786 249824
rect 289998 249704 290004 249756
rect 290056 249744 290062 249756
rect 290182 249744 290188 249756
rect 290056 249716 290188 249744
rect 290056 249704 290062 249716
rect 290182 249704 290188 249716
rect 290240 249704 290246 249756
rect 296898 248412 296904 248464
rect 296956 248452 296962 248464
rect 296990 248452 296996 248464
rect 296956 248424 296996 248452
rect 296956 248412 296962 248424
rect 296990 248412 296996 248424
rect 297048 248412 297054 248464
rect 295518 248344 295524 248396
rect 295576 248384 295582 248396
rect 295794 248384 295800 248396
rect 295576 248356 295800 248384
rect 295576 248344 295582 248356
rect 295794 248344 295800 248356
rect 295852 248344 295858 248396
rect 306742 248384 306748 248396
rect 306703 248356 306748 248384
rect 306742 248344 306748 248356
rect 306800 248344 306806 248396
rect 337102 247160 337108 247172
rect 337063 247132 337108 247160
rect 337102 247120 337108 247132
rect 337160 247120 337166 247172
rect 337102 247024 337108 247036
rect 337063 246996 337108 247024
rect 337102 246984 337108 246996
rect 337160 246984 337166 247036
rect 285950 244984 285956 244996
rect 285911 244956 285956 244984
rect 285950 244944 285956 244956
rect 286008 244944 286014 244996
rect 272150 244440 272156 244452
rect 272111 244412 272156 244440
rect 272150 244400 272156 244412
rect 272208 244400 272214 244452
rect 360286 244264 360292 244316
rect 360344 244304 360350 244316
rect 360470 244304 360476 244316
rect 360344 244276 360476 244304
rect 360344 244264 360350 244276
rect 360470 244264 360476 244276
rect 360528 244264 360534 244316
rect 329926 244196 329932 244248
rect 329984 244236 329990 244248
rect 330202 244236 330208 244248
rect 329984 244208 330208 244236
rect 329984 244196 329990 244208
rect 330202 244196 330208 244208
rect 330260 244196 330266 244248
rect 337102 244236 337108 244248
rect 337063 244208 337108 244236
rect 337102 244196 337108 244208
rect 337160 244196 337166 244248
rect 259549 244171 259607 244177
rect 259549 244137 259561 244171
rect 259595 244168 259607 244171
rect 259638 244168 259644 244180
rect 259595 244140 259644 244168
rect 259595 244137 259607 244140
rect 259549 244131 259607 244137
rect 259638 244128 259644 244140
rect 259696 244128 259702 244180
rect 262674 241584 262680 241596
rect 262600 241556 262680 241584
rect 262600 241528 262628 241556
rect 262674 241544 262680 241556
rect 262732 241544 262738 241596
rect 270770 241584 270776 241596
rect 270696 241556 270776 241584
rect 236270 241476 236276 241528
rect 236328 241516 236334 241528
rect 236454 241516 236460 241528
rect 236328 241488 236460 241516
rect 236328 241476 236334 241488
rect 236454 241476 236460 241488
rect 236512 241476 236518 241528
rect 262582 241476 262588 241528
rect 262640 241476 262646 241528
rect 266630 241476 266636 241528
rect 266688 241516 266694 241528
rect 266722 241516 266728 241528
rect 266688 241488 266728 241516
rect 266688 241476 266694 241488
rect 266722 241476 266728 241488
rect 266780 241476 266786 241528
rect 270696 241460 270724 241556
rect 270770 241544 270776 241556
rect 270828 241544 270834 241596
rect 272150 241584 272156 241596
rect 272111 241556 272156 241584
rect 272150 241544 272156 241556
rect 272208 241544 272214 241596
rect 323486 241584 323492 241596
rect 323412 241556 323492 241584
rect 323412 241528 323440 241556
rect 323486 241544 323492 241556
rect 323544 241544 323550 241596
rect 388990 241544 388996 241596
rect 389048 241584 389054 241596
rect 389266 241584 389272 241596
rect 389048 241556 389272 241584
rect 389048 241544 389054 241556
rect 389266 241544 389272 241556
rect 389324 241544 389330 241596
rect 310701 241519 310759 241525
rect 310701 241485 310713 241519
rect 310747 241516 310759 241519
rect 310882 241516 310888 241528
rect 310747 241488 310888 241516
rect 310747 241485 310759 241488
rect 310701 241479 310759 241485
rect 310882 241476 310888 241488
rect 310940 241476 310946 241528
rect 323394 241476 323400 241528
rect 323452 241476 323458 241528
rect 470594 241516 470600 241528
rect 470555 241488 470600 241516
rect 470594 241476 470600 241488
rect 470652 241476 470658 241528
rect 270678 241408 270684 241460
rect 270736 241408 270742 241460
rect 299474 241408 299480 241460
rect 299532 241448 299538 241460
rect 331398 241448 331404 241460
rect 299532 241420 299577 241448
rect 331359 241420 331404 241448
rect 299532 241408 299538 241420
rect 331398 241408 331404 241420
rect 331456 241408 331462 241460
rect 389266 241448 389272 241460
rect 389227 241420 389272 241448
rect 389266 241408 389272 241420
rect 389324 241408 389330 241460
rect 259638 241340 259644 241392
rect 259696 241380 259702 241392
rect 259822 241380 259828 241392
rect 259696 241352 259828 241380
rect 259696 241340 259702 241352
rect 259822 241340 259828 241352
rect 259880 241340 259886 241392
rect 301314 240224 301320 240236
rect 301056 240196 301320 240224
rect 284754 240116 284760 240168
rect 284812 240156 284818 240168
rect 284938 240156 284944 240168
rect 284812 240128 284944 240156
rect 284812 240116 284818 240128
rect 284938 240116 284944 240128
rect 284996 240116 285002 240168
rect 301056 240100 301084 240196
rect 301314 240184 301320 240196
rect 301372 240184 301378 240236
rect 267734 240088 267740 240100
rect 267695 240060 267740 240088
rect 267734 240048 267740 240060
rect 267792 240048 267798 240100
rect 272150 240088 272156 240100
rect 272111 240060 272156 240088
rect 272150 240048 272156 240060
rect 272208 240048 272214 240100
rect 273530 240048 273536 240100
rect 273588 240088 273594 240100
rect 273622 240088 273628 240100
rect 273588 240060 273628 240088
rect 273588 240048 273594 240060
rect 273622 240048 273628 240060
rect 273680 240048 273686 240100
rect 294322 240048 294328 240100
rect 294380 240088 294386 240100
rect 294414 240088 294420 240100
rect 294380 240060 294420 240088
rect 294380 240048 294386 240060
rect 294414 240048 294420 240060
rect 294472 240048 294478 240100
rect 301038 240048 301044 240100
rect 301096 240048 301102 240100
rect 306742 238756 306748 238808
rect 306800 238796 306806 238808
rect 306929 238799 306987 238805
rect 306929 238796 306941 238799
rect 306800 238768 306941 238796
rect 306800 238756 306806 238768
rect 306929 238765 306941 238768
rect 306975 238765 306987 238799
rect 306929 238759 306987 238765
rect 290366 238728 290372 238740
rect 290327 238700 290372 238728
rect 290366 238688 290372 238700
rect 290424 238688 290430 238740
rect 295610 238728 295616 238740
rect 295571 238700 295616 238728
rect 295610 238688 295616 238700
rect 295668 238688 295674 238740
rect 3050 237328 3056 237380
rect 3108 237368 3114 237380
rect 15838 237368 15844 237380
rect 3108 237340 15844 237368
rect 3108 237328 3114 237340
rect 15838 237328 15844 237340
rect 15896 237328 15902 237380
rect 266722 234852 266728 234864
rect 266683 234824 266728 234852
rect 266722 234812 266728 234824
rect 266780 234812 266786 234864
rect 310882 234716 310888 234728
rect 310808 234688 310888 234716
rect 265158 234608 265164 234660
rect 265216 234608 265222 234660
rect 265176 234512 265204 234608
rect 310808 234592 310836 234688
rect 310882 234676 310888 234688
rect 310940 234676 310946 234728
rect 389269 234651 389327 234657
rect 389269 234617 389281 234651
rect 389315 234648 389327 234651
rect 389450 234648 389456 234660
rect 389315 234620 389456 234648
rect 389315 234617 389327 234620
rect 389269 234611 389327 234617
rect 389450 234608 389456 234620
rect 389508 234608 389514 234660
rect 310790 234540 310796 234592
rect 310848 234540 310854 234592
rect 374362 234540 374368 234592
rect 374420 234540 374426 234592
rect 375834 234540 375840 234592
rect 375892 234540 375898 234592
rect 265250 234512 265256 234524
rect 265176 234484 265256 234512
rect 265250 234472 265256 234484
rect 265308 234472 265314 234524
rect 272153 234515 272211 234521
rect 272153 234481 272165 234515
rect 272199 234512 272211 234515
rect 272242 234512 272248 234524
rect 272199 234484 272248 234512
rect 272199 234481 272211 234484
rect 272153 234475 272211 234481
rect 272242 234472 272248 234484
rect 272300 234472 272306 234524
rect 285950 234512 285956 234524
rect 285911 234484 285956 234512
rect 285950 234472 285956 234484
rect 286008 234472 286014 234524
rect 374380 234456 374408 234540
rect 375852 234456 375880 234540
rect 374362 234404 374368 234456
rect 374420 234404 374426 234456
rect 375834 234404 375840 234456
rect 375892 234404 375898 234456
rect 235074 231820 235080 231872
rect 235132 231860 235138 231872
rect 235166 231860 235172 231872
rect 235132 231832 235172 231860
rect 235132 231820 235138 231832
rect 235166 231820 235172 231832
rect 235224 231820 235230 231872
rect 244274 231820 244280 231872
rect 244332 231860 244338 231872
rect 244458 231860 244464 231872
rect 244332 231832 244464 231860
rect 244332 231820 244338 231832
rect 244458 231820 244464 231832
rect 244516 231820 244522 231872
rect 250070 231820 250076 231872
rect 250128 231860 250134 231872
rect 250346 231860 250352 231872
rect 250128 231832 250352 231860
rect 250128 231820 250134 231832
rect 250346 231820 250352 231832
rect 250404 231820 250410 231872
rect 251450 231820 251456 231872
rect 251508 231860 251514 231872
rect 251634 231860 251640 231872
rect 251508 231832 251640 231860
rect 251508 231820 251514 231832
rect 251634 231820 251640 231832
rect 251692 231820 251698 231872
rect 299474 231820 299480 231872
rect 299532 231860 299538 231872
rect 299532 231832 299577 231860
rect 299532 231820 299538 231832
rect 323302 231820 323308 231872
rect 323360 231860 323366 231872
rect 323486 231860 323492 231872
rect 323360 231832 323492 231860
rect 323360 231820 323366 231832
rect 323486 231820 323492 231832
rect 323544 231820 323550 231872
rect 324682 231820 324688 231872
rect 324740 231860 324746 231872
rect 324774 231860 324780 231872
rect 324740 231832 324780 231860
rect 324740 231820 324746 231832
rect 324774 231820 324780 231832
rect 324832 231820 324838 231872
rect 331398 231860 331404 231872
rect 331359 231832 331404 231860
rect 331398 231820 331404 231832
rect 331456 231820 331462 231872
rect 338666 231820 338672 231872
rect 338724 231860 338730 231872
rect 338850 231860 338856 231872
rect 338724 231832 338856 231860
rect 338724 231820 338730 231832
rect 338850 231820 338856 231832
rect 338908 231820 338914 231872
rect 341058 231820 341064 231872
rect 341116 231860 341122 231872
rect 341150 231860 341156 231872
rect 341116 231832 341156 231860
rect 341116 231820 341122 231832
rect 341150 231820 341156 231832
rect 341208 231820 341214 231872
rect 372522 231820 372528 231872
rect 372580 231860 372586 231872
rect 372706 231860 372712 231872
rect 372580 231832 372712 231860
rect 372580 231820 372586 231832
rect 372706 231820 372712 231832
rect 372764 231820 372770 231872
rect 376938 231820 376944 231872
rect 376996 231860 377002 231872
rect 377122 231860 377128 231872
rect 376996 231832 377128 231860
rect 376996 231820 377002 231832
rect 377122 231820 377128 231832
rect 377180 231820 377186 231872
rect 267737 231795 267795 231801
rect 267737 231761 267749 231795
rect 267783 231792 267795 231795
rect 267918 231792 267924 231804
rect 267783 231764 267924 231792
rect 267783 231761 267795 231764
rect 267737 231755 267795 231761
rect 267918 231752 267924 231764
rect 267976 231752 267982 231804
rect 310790 231792 310796 231804
rect 310751 231764 310796 231792
rect 310790 231752 310796 231764
rect 310848 231752 310854 231804
rect 337105 231659 337163 231665
rect 337105 231625 337117 231659
rect 337151 231656 337163 231659
rect 337194 231656 337200 231668
rect 337151 231628 337200 231656
rect 337151 231625 337163 231628
rect 337105 231619 337163 231625
rect 337194 231616 337200 231628
rect 337252 231616 337258 231668
rect 266722 230500 266728 230512
rect 266683 230472 266728 230500
rect 266722 230460 266728 230472
rect 266780 230460 266786 230512
rect 301038 230460 301044 230512
rect 301096 230500 301102 230512
rect 301222 230500 301228 230512
rect 301096 230472 301228 230500
rect 301096 230460 301102 230472
rect 301222 230460 301228 230472
rect 301280 230460 301286 230512
rect 306834 230460 306840 230512
rect 306892 230500 306898 230512
rect 306929 230503 306987 230509
rect 306929 230500 306941 230503
rect 306892 230472 306941 230500
rect 306892 230460 306898 230472
rect 306929 230469 306941 230472
rect 306975 230469 306987 230503
rect 306929 230463 306987 230469
rect 327166 230460 327172 230512
rect 327224 230500 327230 230512
rect 327350 230500 327356 230512
rect 327224 230472 327356 230500
rect 327224 230460 327230 230472
rect 327350 230460 327356 230472
rect 327408 230460 327414 230512
rect 358538 230460 358544 230512
rect 358596 230500 358602 230512
rect 358722 230500 358728 230512
rect 358596 230472 358728 230500
rect 358596 230460 358602 230472
rect 358722 230460 358728 230472
rect 358780 230460 358786 230512
rect 290366 230432 290372 230444
rect 290327 230404 290372 230432
rect 290366 230392 290372 230404
rect 290424 230392 290430 230444
rect 295610 229140 295616 229152
rect 295571 229112 295616 229140
rect 295610 229100 295616 229112
rect 295668 229100 295674 229152
rect 270678 224992 270684 225004
rect 270639 224964 270684 224992
rect 270678 224952 270684 224964
rect 270736 224952 270742 225004
rect 341061 224995 341119 225001
rect 341061 224961 341073 224995
rect 341107 224992 341119 224995
rect 341150 224992 341156 225004
rect 341107 224964 341156 224992
rect 341107 224961 341119 224964
rect 341061 224955 341119 224961
rect 341150 224952 341156 224964
rect 341208 224952 341214 225004
rect 360286 224952 360292 225004
rect 360344 224992 360350 225004
rect 360470 224992 360476 225004
rect 360344 224964 360476 224992
rect 360344 224952 360350 224964
rect 360470 224952 360476 224964
rect 360528 224952 360534 225004
rect 301222 222272 301228 222284
rect 301056 222244 301228 222272
rect 236270 222164 236276 222216
rect 236328 222204 236334 222216
rect 236454 222204 236460 222216
rect 236328 222176 236460 222204
rect 236328 222164 236334 222176
rect 236454 222164 236460 222176
rect 236512 222164 236518 222216
rect 259638 222164 259644 222216
rect 259696 222204 259702 222216
rect 259822 222204 259828 222216
rect 259696 222176 259828 222204
rect 259696 222164 259702 222176
rect 259822 222164 259828 222176
rect 259880 222164 259886 222216
rect 262674 222164 262680 222216
rect 262732 222204 262738 222216
rect 262766 222204 262772 222216
rect 262732 222176 262772 222204
rect 262732 222164 262738 222176
rect 262766 222164 262772 222176
rect 262824 222164 262830 222216
rect 265158 222164 265164 222216
rect 265216 222204 265222 222216
rect 265342 222204 265348 222216
rect 265216 222176 265348 222204
rect 265216 222164 265222 222176
rect 265342 222164 265348 222176
rect 265400 222164 265406 222216
rect 284754 222164 284760 222216
rect 284812 222164 284818 222216
rect 295518 222164 295524 222216
rect 295576 222204 295582 222216
rect 295610 222204 295616 222216
rect 295576 222176 295616 222204
rect 295576 222164 295582 222176
rect 295610 222164 295616 222176
rect 295668 222164 295674 222216
rect 284772 222080 284800 222164
rect 301056 222148 301084 222244
rect 301222 222232 301228 222244
rect 301280 222232 301286 222284
rect 302510 222164 302516 222216
rect 302568 222204 302574 222216
rect 302694 222204 302700 222216
rect 302568 222176 302700 222204
rect 302568 222164 302574 222176
rect 302694 222164 302700 222176
rect 302752 222164 302758 222216
rect 310793 222207 310851 222213
rect 310793 222173 310805 222207
rect 310839 222204 310851 222207
rect 310882 222204 310888 222216
rect 310839 222176 310888 222204
rect 310839 222173 310851 222176
rect 310793 222167 310851 222173
rect 310882 222164 310888 222176
rect 310940 222164 310946 222216
rect 324682 222164 324688 222216
rect 324740 222204 324746 222216
rect 324774 222204 324780 222216
rect 324740 222176 324780 222204
rect 324740 222164 324746 222176
rect 324774 222164 324780 222176
rect 324832 222164 324838 222216
rect 341058 222204 341064 222216
rect 341019 222176 341064 222204
rect 341058 222164 341064 222176
rect 341116 222164 341122 222216
rect 389266 222164 389272 222216
rect 389324 222204 389330 222216
rect 389542 222204 389548 222216
rect 389324 222176 389548 222204
rect 389324 222164 389330 222176
rect 389542 222164 389548 222176
rect 389600 222164 389606 222216
rect 463786 222164 463792 222216
rect 463844 222204 463850 222216
rect 464062 222204 464068 222216
rect 463844 222176 464068 222204
rect 463844 222164 463850 222176
rect 464062 222164 464068 222176
rect 464120 222164 464126 222216
rect 470410 222164 470416 222216
rect 470468 222204 470474 222216
rect 470594 222204 470600 222216
rect 470468 222176 470600 222204
rect 470468 222164 470474 222176
rect 470594 222164 470600 222176
rect 470652 222164 470658 222216
rect 299474 222096 299480 222148
rect 299532 222136 299538 222148
rect 299532 222108 299577 222136
rect 299532 222096 299538 222108
rect 301038 222096 301044 222148
rect 301096 222096 301102 222148
rect 259638 222028 259644 222080
rect 259696 222068 259702 222080
rect 259822 222068 259828 222080
rect 259696 222040 259828 222068
rect 259696 222028 259702 222040
rect 259822 222028 259828 222040
rect 259880 222028 259886 222080
rect 284754 222028 284760 222080
rect 284812 222028 284818 222080
rect 270678 220844 270684 220856
rect 270639 220816 270684 220844
rect 270678 220804 270684 220816
rect 270736 220804 270742 220856
rect 288894 220804 288900 220856
rect 288952 220844 288958 220856
rect 289078 220844 289084 220856
rect 288952 220816 289084 220844
rect 288952 220804 288958 220816
rect 289078 220804 289084 220816
rect 289136 220804 289142 220856
rect 290182 220804 290188 220856
rect 290240 220844 290246 220856
rect 290366 220844 290372 220856
rect 290240 220816 290372 220844
rect 290240 220804 290246 220816
rect 290366 220804 290372 220816
rect 290424 220804 290430 220856
rect 291654 220804 291660 220856
rect 291712 220844 291718 220856
rect 291930 220844 291936 220856
rect 291712 220816 291936 220844
rect 291712 220804 291718 220816
rect 291930 220804 291936 220816
rect 291988 220804 291994 220856
rect 294322 220804 294328 220856
rect 294380 220844 294386 220856
rect 294414 220844 294420 220856
rect 294380 220816 294420 220844
rect 294380 220804 294386 220816
rect 294414 220804 294420 220816
rect 294472 220804 294478 220856
rect 337105 220847 337163 220853
rect 337105 220813 337117 220847
rect 337151 220844 337163 220847
rect 337286 220844 337292 220856
rect 337151 220816 337292 220844
rect 337151 220813 337163 220816
rect 337105 220807 337163 220813
rect 337286 220804 337292 220816
rect 337344 220804 337350 220856
rect 290182 219416 290188 219428
rect 290143 219388 290188 219416
rect 290182 219376 290188 219388
rect 290240 219376 290246 219428
rect 291654 219416 291660 219428
rect 291615 219388 291660 219416
rect 291654 219376 291660 219388
rect 291712 219376 291718 219428
rect 317506 219376 317512 219428
rect 317564 219416 317570 219428
rect 317690 219416 317696 219428
rect 317564 219388 317696 219416
rect 317564 219376 317570 219388
rect 317690 219376 317696 219388
rect 317748 219376 317754 219428
rect 310882 215404 310888 215416
rect 310808 215376 310888 215404
rect 310808 215280 310836 215376
rect 310882 215364 310888 215376
rect 310940 215364 310946 215416
rect 389542 215404 389548 215416
rect 389468 215376 389548 215404
rect 389468 215280 389496 215376
rect 389542 215364 389548 215376
rect 389600 215364 389606 215416
rect 464062 215404 464068 215416
rect 463988 215376 464068 215404
rect 463988 215280 464016 215376
rect 464062 215364 464068 215376
rect 464120 215364 464126 215416
rect 273438 215228 273444 215280
rect 273496 215268 273502 215280
rect 273622 215268 273628 215280
rect 273496 215240 273628 215268
rect 273496 215228 273502 215240
rect 273622 215228 273628 215240
rect 273680 215228 273686 215280
rect 310790 215228 310796 215280
rect 310848 215228 310854 215280
rect 374362 215228 374368 215280
rect 374420 215228 374426 215280
rect 375834 215228 375840 215280
rect 375892 215228 375898 215280
rect 389450 215228 389456 215280
rect 389508 215228 389514 215280
rect 463970 215228 463976 215280
rect 464028 215228 464034 215280
rect 374380 215144 374408 215228
rect 375852 215144 375880 215228
rect 374362 215092 374368 215144
rect 374420 215092 374426 215144
rect 375834 215092 375840 215144
rect 375892 215092 375898 215144
rect 337286 212616 337292 212628
rect 337212 212588 337292 212616
rect 235074 212508 235080 212560
rect 235132 212548 235138 212560
rect 235166 212548 235172 212560
rect 235132 212520 235172 212548
rect 235132 212508 235138 212520
rect 235166 212508 235172 212520
rect 235224 212508 235230 212560
rect 244274 212508 244280 212560
rect 244332 212548 244338 212560
rect 244458 212548 244464 212560
rect 244332 212520 244464 212548
rect 244332 212508 244338 212520
rect 244458 212508 244464 212520
rect 244516 212508 244522 212560
rect 250070 212508 250076 212560
rect 250128 212548 250134 212560
rect 250346 212548 250352 212560
rect 250128 212520 250352 212548
rect 250128 212508 250134 212520
rect 250346 212508 250352 212520
rect 250404 212508 250410 212560
rect 251450 212508 251456 212560
rect 251508 212548 251514 212560
rect 251634 212548 251640 212560
rect 251508 212520 251640 212548
rect 251508 212508 251514 212520
rect 251634 212508 251640 212520
rect 251692 212508 251698 212560
rect 265158 212508 265164 212560
rect 265216 212548 265222 212560
rect 265250 212548 265256 212560
rect 265216 212520 265256 212548
rect 265216 212508 265222 212520
rect 265250 212508 265256 212520
rect 265308 212508 265314 212560
rect 266630 212508 266636 212560
rect 266688 212548 266694 212560
rect 266814 212548 266820 212560
rect 266688 212520 266820 212548
rect 266688 212508 266694 212520
rect 266814 212508 266820 212520
rect 266872 212508 266878 212560
rect 267826 212508 267832 212560
rect 267884 212548 267890 212560
rect 267918 212548 267924 212560
rect 267884 212520 267924 212548
rect 267884 212508 267890 212520
rect 267918 212508 267924 212520
rect 267976 212508 267982 212560
rect 284754 212508 284760 212560
rect 284812 212508 284818 212560
rect 299474 212508 299480 212560
rect 299532 212548 299538 212560
rect 299532 212520 299577 212548
rect 299532 212508 299538 212520
rect 323302 212508 323308 212560
rect 323360 212548 323366 212560
rect 323486 212548 323492 212560
rect 323360 212520 323492 212548
rect 323360 212508 323366 212520
rect 323486 212508 323492 212520
rect 323544 212508 323550 212560
rect 324682 212508 324688 212560
rect 324740 212548 324746 212560
rect 324774 212548 324780 212560
rect 324740 212520 324780 212548
rect 324740 212508 324746 212520
rect 324774 212508 324780 212520
rect 324832 212508 324838 212560
rect 331398 212508 331404 212560
rect 331456 212548 331462 212560
rect 331582 212548 331588 212560
rect 331456 212520 331588 212548
rect 331456 212508 331462 212520
rect 331582 212508 331588 212520
rect 331640 212508 331646 212560
rect 284772 212480 284800 212508
rect 337212 212492 337240 212588
rect 337286 212576 337292 212588
rect 337344 212576 337350 212628
rect 338666 212508 338672 212560
rect 338724 212548 338730 212560
rect 338850 212548 338856 212560
rect 338724 212520 338856 212548
rect 338724 212508 338730 212520
rect 338850 212508 338856 212520
rect 338908 212508 338914 212560
rect 372522 212508 372528 212560
rect 372580 212548 372586 212560
rect 372706 212548 372712 212560
rect 372580 212520 372712 212548
rect 372580 212508 372586 212520
rect 372706 212508 372712 212520
rect 372764 212508 372770 212560
rect 376938 212508 376944 212560
rect 376996 212548 377002 212560
rect 377122 212548 377128 212560
rect 376996 212520 377128 212548
rect 376996 212508 377002 212520
rect 377122 212508 377128 212520
rect 377180 212508 377186 212560
rect 284938 212480 284944 212492
rect 284772 212452 284944 212480
rect 284938 212440 284944 212452
rect 284996 212440 285002 212492
rect 290182 212480 290188 212492
rect 290143 212452 290188 212480
rect 290182 212440 290188 212452
rect 290240 212440 290246 212492
rect 291654 212480 291660 212492
rect 291615 212452 291660 212480
rect 291654 212440 291660 212452
rect 291712 212440 291718 212492
rect 310790 212480 310796 212492
rect 310751 212452 310796 212480
rect 310790 212440 310796 212452
rect 310848 212440 310854 212492
rect 337194 212440 337200 212492
rect 337252 212440 337258 212492
rect 299842 211148 299848 211200
rect 299900 211188 299906 211200
rect 299934 211188 299940 211200
rect 299900 211160 299940 211188
rect 299900 211148 299906 211160
rect 299934 211148 299940 211160
rect 299992 211148 299998 211200
rect 250070 211080 250076 211132
rect 250128 211120 250134 211132
rect 250254 211120 250260 211132
rect 250128 211092 250260 211120
rect 250128 211080 250134 211092
rect 250254 211080 250260 211092
rect 250312 211080 250318 211132
rect 267826 211080 267832 211132
rect 267884 211120 267890 211132
rect 267918 211120 267924 211132
rect 267884 211092 267924 211120
rect 267884 211080 267890 211092
rect 267918 211080 267924 211092
rect 267976 211080 267982 211132
rect 294230 211080 294236 211132
rect 294288 211120 294294 211132
rect 294322 211120 294328 211132
rect 294288 211092 294328 211120
rect 294288 211080 294294 211092
rect 294322 211080 294328 211092
rect 294380 211080 294386 211132
rect 306650 211080 306656 211132
rect 306708 211120 306714 211132
rect 306834 211120 306840 211132
rect 306708 211092 306840 211120
rect 306708 211080 306714 211092
rect 306834 211080 306840 211092
rect 306892 211080 306898 211132
rect 337194 211080 337200 211132
rect 337252 211120 337258 211132
rect 337378 211120 337384 211132
rect 337252 211092 337384 211120
rect 337252 211080 337258 211092
rect 337378 211080 337384 211092
rect 337436 211080 337442 211132
rect 317506 209788 317512 209840
rect 317564 209828 317570 209840
rect 317690 209828 317696 209840
rect 317564 209800 317696 209828
rect 317564 209788 317570 209800
rect 317690 209788 317696 209800
rect 317748 209788 317754 209840
rect 306650 209720 306656 209772
rect 306708 209760 306714 209772
rect 306926 209760 306932 209772
rect 306708 209732 306932 209760
rect 306708 209720 306714 209732
rect 306926 209720 306932 209732
rect 306984 209720 306990 209772
rect 341242 209720 341248 209772
rect 341300 209760 341306 209772
rect 341334 209760 341340 209772
rect 341300 209732 341340 209760
rect 341300 209720 341306 209732
rect 341334 209720 341340 209732
rect 341392 209720 341398 209772
rect 262582 207884 262588 207936
rect 262640 207924 262646 207936
rect 262766 207924 262772 207936
rect 262640 207896 262772 207924
rect 262640 207884 262646 207896
rect 262766 207884 262772 207896
rect 262824 207884 262830 207936
rect 302602 207788 302608 207800
rect 302563 207760 302608 207788
rect 302602 207748 302608 207760
rect 302660 207748 302666 207800
rect 266630 205640 266636 205692
rect 266688 205640 266694 205692
rect 270678 205680 270684 205692
rect 270639 205652 270684 205680
rect 270678 205640 270684 205652
rect 270736 205640 270742 205692
rect 323302 205640 323308 205692
rect 323360 205640 323366 205692
rect 360286 205640 360292 205692
rect 360344 205680 360350 205692
rect 360470 205680 360476 205692
rect 360344 205652 360476 205680
rect 360344 205640 360350 205652
rect 360470 205640 360476 205652
rect 360528 205640 360534 205692
rect 266648 205612 266676 205640
rect 266722 205612 266728 205624
rect 266648 205584 266728 205612
rect 266722 205572 266728 205584
rect 266780 205572 266786 205624
rect 323320 205544 323348 205640
rect 323394 205544 323400 205556
rect 323320 205516 323400 205544
rect 323394 205504 323400 205516
rect 323452 205504 323458 205556
rect 236270 202852 236276 202904
rect 236328 202892 236334 202904
rect 236454 202892 236460 202904
rect 236328 202864 236460 202892
rect 236328 202852 236334 202864
rect 236454 202852 236460 202864
rect 236512 202852 236518 202904
rect 270678 202892 270684 202904
rect 270639 202864 270684 202892
rect 270678 202852 270684 202864
rect 270736 202852 270742 202904
rect 285950 202852 285956 202904
rect 286008 202892 286014 202904
rect 286134 202892 286140 202904
rect 286008 202864 286140 202892
rect 286008 202852 286014 202864
rect 286134 202852 286140 202864
rect 286192 202852 286198 202904
rect 295518 202852 295524 202904
rect 295576 202892 295582 202904
rect 295610 202892 295616 202904
rect 295576 202864 295616 202892
rect 295576 202852 295582 202864
rect 295610 202852 295616 202864
rect 295668 202852 295674 202904
rect 296806 202852 296812 202904
rect 296864 202892 296870 202904
rect 296898 202892 296904 202904
rect 296864 202864 296904 202892
rect 296864 202852 296870 202864
rect 296898 202852 296904 202864
rect 296956 202852 296962 202904
rect 302602 202892 302608 202904
rect 302563 202864 302608 202892
rect 302602 202852 302608 202864
rect 302660 202852 302666 202904
rect 310793 202895 310851 202901
rect 310793 202861 310805 202895
rect 310839 202892 310851 202895
rect 310882 202892 310888 202904
rect 310839 202864 310888 202892
rect 310839 202861 310851 202864
rect 310793 202855 310851 202861
rect 310882 202852 310888 202864
rect 310940 202852 310946 202904
rect 324590 202852 324596 202904
rect 324648 202892 324654 202904
rect 324682 202892 324688 202904
rect 324648 202864 324688 202892
rect 324648 202852 324654 202864
rect 324682 202852 324688 202864
rect 324740 202852 324746 202904
rect 329926 202852 329932 202904
rect 329984 202892 329990 202904
rect 330110 202892 330116 202904
rect 329984 202864 330116 202892
rect 329984 202852 329990 202864
rect 330110 202852 330116 202864
rect 330168 202852 330174 202904
rect 389266 202852 389272 202904
rect 389324 202892 389330 202904
rect 389542 202892 389548 202904
rect 389324 202864 389548 202892
rect 389324 202852 389330 202864
rect 389542 202852 389548 202864
rect 389600 202852 389606 202904
rect 463786 202852 463792 202904
rect 463844 202892 463850 202904
rect 464062 202892 464068 202904
rect 463844 202864 464068 202892
rect 463844 202852 463850 202864
rect 464062 202852 464068 202864
rect 464120 202852 464126 202904
rect 470410 202852 470416 202904
rect 470468 202892 470474 202904
rect 470594 202892 470600 202904
rect 470468 202864 470600 202892
rect 470468 202852 470474 202864
rect 470594 202852 470600 202864
rect 470652 202852 470658 202904
rect 273530 202784 273536 202836
rect 273588 202824 273594 202836
rect 273622 202824 273628 202836
rect 273588 202796 273628 202824
rect 273588 202784 273594 202796
rect 273622 202784 273628 202796
rect 273680 202784 273686 202836
rect 250070 201424 250076 201476
rect 250128 201464 250134 201476
rect 250346 201464 250352 201476
rect 250128 201436 250352 201464
rect 250128 201424 250134 201436
rect 250346 201424 250352 201436
rect 250404 201424 250410 201476
rect 301038 201424 301044 201476
rect 301096 201424 301102 201476
rect 301056 201396 301084 201424
rect 301130 201396 301136 201408
rect 301056 201368 301136 201396
rect 301130 201356 301136 201368
rect 301188 201356 301194 201408
rect 250070 200104 250076 200116
rect 250031 200076 250076 200104
rect 250070 200064 250076 200076
rect 250128 200064 250134 200116
rect 289906 200064 289912 200116
rect 289964 200104 289970 200116
rect 290182 200104 290188 200116
rect 289964 200076 290188 200104
rect 289964 200064 289970 200076
rect 290182 200064 290188 200076
rect 290240 200064 290246 200116
rect 291378 200064 291384 200116
rect 291436 200104 291442 200116
rect 291654 200104 291660 200116
rect 291436 200076 291660 200104
rect 291436 200064 291442 200076
rect 291654 200064 291660 200076
rect 291712 200064 291718 200116
rect 299750 200064 299756 200116
rect 299808 200104 299814 200116
rect 299842 200104 299848 200116
rect 299808 200076 299848 200104
rect 299808 200064 299814 200076
rect 299842 200064 299848 200076
rect 299900 200064 299906 200116
rect 306742 200064 306748 200116
rect 306800 200104 306806 200116
rect 306834 200104 306840 200116
rect 306800 200076 306840 200104
rect 306800 200064 306806 200076
rect 306834 200064 306840 200076
rect 306892 200064 306898 200116
rect 317506 200064 317512 200116
rect 317564 200104 317570 200116
rect 317690 200104 317696 200116
rect 317564 200076 317696 200104
rect 317564 200064 317570 200076
rect 317690 200064 317696 200076
rect 317748 200064 317754 200116
rect 341242 198704 341248 198756
rect 341300 198744 341306 198756
rect 341334 198744 341340 198756
rect 341300 198716 341340 198744
rect 341300 198704 341306 198716
rect 341334 198704 341340 198716
rect 341392 198704 341398 198756
rect 266722 198132 266728 198144
rect 266648 198104 266728 198132
rect 266648 198076 266676 198104
rect 266722 198092 266728 198104
rect 266780 198092 266786 198144
rect 266630 198024 266636 198076
rect 266688 198024 266694 198076
rect 285766 198024 285772 198076
rect 285824 198064 285830 198076
rect 285950 198064 285956 198076
rect 285824 198036 285956 198064
rect 285824 198024 285830 198036
rect 285950 198024 285956 198036
rect 286008 198024 286014 198076
rect 294230 198024 294236 198076
rect 294288 198064 294294 198076
rect 294414 198064 294420 198076
rect 294288 198036 294420 198064
rect 294288 198024 294294 198036
rect 294414 198024 294420 198036
rect 294472 198024 294478 198076
rect 329926 198024 329932 198076
rect 329984 198064 329990 198076
rect 330110 198064 330116 198076
rect 329984 198036 330116 198064
rect 329984 198024 329990 198036
rect 330110 198024 330116 198036
rect 330168 198024 330174 198076
rect 310882 196092 310888 196104
rect 310808 196064 310888 196092
rect 310808 195968 310836 196064
rect 310882 196052 310888 196064
rect 310940 196052 310946 196104
rect 389542 196092 389548 196104
rect 389468 196064 389548 196092
rect 389468 195968 389496 196064
rect 389542 196052 389548 196064
rect 389600 196052 389606 196104
rect 464062 196092 464068 196104
rect 463988 196064 464068 196092
rect 463988 195968 464016 196064
rect 464062 196052 464068 196064
rect 464120 196052 464126 196104
rect 310790 195916 310796 195968
rect 310848 195916 310854 195968
rect 357526 195916 357532 195968
rect 357584 195956 357590 195968
rect 357710 195956 357716 195968
rect 357584 195928 357716 195956
rect 357584 195916 357590 195928
rect 357710 195916 357716 195928
rect 357768 195916 357774 195968
rect 374362 195916 374368 195968
rect 374420 195916 374426 195968
rect 375834 195916 375840 195968
rect 375892 195916 375898 195968
rect 389450 195916 389456 195968
rect 389508 195916 389514 195968
rect 463970 195916 463976 195968
rect 464028 195916 464034 195968
rect 374380 195832 374408 195916
rect 375852 195832 375880 195916
rect 374362 195780 374368 195832
rect 374420 195780 374426 195832
rect 375834 195780 375840 195832
rect 375892 195780 375898 195832
rect 288710 193332 288716 193384
rect 288768 193332 288774 193384
rect 337102 193332 337108 193384
rect 337160 193332 337166 193384
rect 288728 193248 288756 193332
rect 337120 193248 337148 193332
rect 230842 193196 230848 193248
rect 230900 193236 230906 193248
rect 231026 193236 231032 193248
rect 230900 193208 231032 193236
rect 230900 193196 230906 193208
rect 231026 193196 231032 193208
rect 231084 193196 231090 193248
rect 235074 193196 235080 193248
rect 235132 193236 235138 193248
rect 235166 193236 235172 193248
rect 235132 193208 235172 193236
rect 235132 193196 235138 193208
rect 235166 193196 235172 193208
rect 235224 193196 235230 193248
rect 239122 193196 239128 193248
rect 239180 193236 239186 193248
rect 239214 193236 239220 193248
rect 239180 193208 239220 193236
rect 239180 193196 239186 193208
rect 239214 193196 239220 193208
rect 239272 193196 239278 193248
rect 244274 193196 244280 193248
rect 244332 193236 244338 193248
rect 244458 193236 244464 193248
rect 244332 193208 244464 193236
rect 244332 193196 244338 193208
rect 244458 193196 244464 193208
rect 244516 193196 244522 193248
rect 251450 193196 251456 193248
rect 251508 193236 251514 193248
rect 251634 193236 251640 193248
rect 251508 193208 251640 193236
rect 251508 193196 251514 193208
rect 251634 193196 251640 193208
rect 251692 193196 251698 193248
rect 259730 193196 259736 193248
rect 259788 193236 259794 193248
rect 259914 193236 259920 193248
rect 259788 193208 259920 193236
rect 259788 193196 259794 193208
rect 259914 193196 259920 193208
rect 259972 193196 259978 193248
rect 265250 193196 265256 193248
rect 265308 193236 265314 193248
rect 265342 193236 265348 193248
rect 265308 193208 265348 193236
rect 265308 193196 265314 193208
rect 265342 193196 265348 193208
rect 265400 193196 265406 193248
rect 267826 193196 267832 193248
rect 267884 193236 267890 193248
rect 267918 193236 267924 193248
rect 267884 193208 267924 193236
rect 267884 193196 267890 193208
rect 267918 193196 267924 193208
rect 267976 193196 267982 193248
rect 288710 193196 288716 193248
rect 288768 193196 288774 193248
rect 323302 193196 323308 193248
rect 323360 193236 323366 193248
rect 323486 193236 323492 193248
rect 323360 193208 323492 193236
rect 323360 193196 323366 193208
rect 323486 193196 323492 193208
rect 323544 193196 323550 193248
rect 324590 193196 324596 193248
rect 324648 193236 324654 193248
rect 324682 193236 324688 193248
rect 324648 193208 324688 193236
rect 324648 193196 324654 193208
rect 324682 193196 324688 193208
rect 324740 193196 324746 193248
rect 331398 193196 331404 193248
rect 331456 193236 331462 193248
rect 331582 193236 331588 193248
rect 331456 193208 331588 193236
rect 331456 193196 331462 193208
rect 331582 193196 331588 193208
rect 331640 193196 331646 193248
rect 337102 193196 337108 193248
rect 337160 193196 337166 193248
rect 338666 193196 338672 193248
rect 338724 193236 338730 193248
rect 338850 193236 338856 193248
rect 338724 193208 338856 193236
rect 338724 193196 338730 193208
rect 338850 193196 338856 193208
rect 338908 193196 338914 193248
rect 372522 193196 372528 193248
rect 372580 193236 372586 193248
rect 372706 193236 372712 193248
rect 372580 193208 372712 193236
rect 372580 193196 372586 193208
rect 372706 193196 372712 193208
rect 372764 193196 372770 193248
rect 376938 193196 376944 193248
rect 376996 193236 377002 193248
rect 377122 193236 377128 193248
rect 376996 193208 377128 193236
rect 376996 193196 377002 193208
rect 377122 193196 377128 193208
rect 377180 193196 377186 193248
rect 367002 193168 367008 193180
rect 366963 193140 367008 193168
rect 367002 193128 367008 193140
rect 367060 193128 367066 193180
rect 324682 191768 324688 191820
rect 324740 191808 324746 191820
rect 324866 191808 324872 191820
rect 324740 191780 324872 191808
rect 324740 191768 324746 191780
rect 324866 191768 324872 191780
rect 324924 191768 324930 191820
rect 358538 191768 358544 191820
rect 358596 191808 358602 191820
rect 358814 191808 358820 191820
rect 358596 191780 358820 191808
rect 358596 191768 358602 191780
rect 358814 191768 358820 191780
rect 358872 191768 358878 191820
rect 317506 190476 317512 190528
rect 317564 190516 317570 190528
rect 317690 190516 317696 190528
rect 317564 190488 317696 190516
rect 317564 190476 317570 190488
rect 317690 190476 317696 190488
rect 317748 190476 317754 190528
rect 264974 190408 264980 190460
rect 265032 190448 265038 190460
rect 265250 190448 265256 190460
rect 265032 190420 265256 190448
rect 265032 190408 265038 190420
rect 265250 190408 265256 190420
rect 265308 190408 265314 190460
rect 299842 190448 299848 190460
rect 299803 190420 299848 190448
rect 299842 190408 299848 190420
rect 299900 190408 299906 190460
rect 302513 190451 302571 190457
rect 302513 190417 302525 190451
rect 302559 190448 302571 190451
rect 302786 190448 302792 190460
rect 302559 190420 302792 190448
rect 302559 190417 302571 190420
rect 302513 190411 302571 190417
rect 302786 190408 302792 190420
rect 302844 190408 302850 190460
rect 306834 190448 306840 190460
rect 306795 190420 306840 190448
rect 306834 190408 306840 190420
rect 306892 190408 306898 190460
rect 288710 189020 288716 189032
rect 288671 188992 288716 189020
rect 288710 188980 288716 188992
rect 288768 188980 288774 189032
rect 341242 188980 341248 189032
rect 341300 189020 341306 189032
rect 341426 189020 341432 189032
rect 341300 188992 341432 189020
rect 341300 188980 341306 188992
rect 341426 188980 341432 188992
rect 341484 188980 341490 189032
rect 339770 188408 339776 188420
rect 339731 188380 339776 188408
rect 339770 188368 339776 188380
rect 339828 188368 339834 188420
rect 330110 186940 330116 186992
rect 330168 186980 330174 186992
rect 330294 186980 330300 186992
rect 330168 186952 330300 186980
rect 330168 186940 330174 186952
rect 330294 186940 330300 186952
rect 330352 186940 330358 186992
rect 296898 186436 296904 186448
rect 296824 186408 296904 186436
rect 266630 186328 266636 186380
rect 266688 186328 266694 186380
rect 267734 186368 267740 186380
rect 267695 186340 267740 186368
rect 267734 186328 267740 186340
rect 267792 186328 267798 186380
rect 270678 186368 270684 186380
rect 270639 186340 270684 186368
rect 270678 186328 270684 186340
rect 270736 186328 270742 186380
rect 295610 186368 295616 186380
rect 295536 186340 295616 186368
rect 250070 186300 250076 186312
rect 250031 186272 250076 186300
rect 250070 186260 250076 186272
rect 250128 186260 250134 186312
rect 266648 186232 266676 186328
rect 295536 186312 295564 186340
rect 295610 186328 295616 186340
rect 295668 186328 295674 186380
rect 296824 186312 296852 186408
rect 296898 186396 296904 186408
rect 296956 186396 296962 186448
rect 327258 186436 327264 186448
rect 327184 186408 327264 186436
rect 327184 186312 327212 186408
rect 327258 186396 327264 186408
rect 327316 186396 327322 186448
rect 295518 186260 295524 186312
rect 295576 186260 295582 186312
rect 296806 186260 296812 186312
rect 296864 186260 296870 186312
rect 327166 186260 327172 186312
rect 327224 186260 327230 186312
rect 266722 186232 266728 186244
rect 266648 186204 266728 186232
rect 266722 186192 266728 186204
rect 266780 186192 266786 186244
rect 236270 183540 236276 183592
rect 236328 183580 236334 183592
rect 236454 183580 236460 183592
rect 236328 183552 236460 183580
rect 236328 183540 236334 183552
rect 236454 183540 236460 183552
rect 236512 183540 236518 183592
rect 267734 183580 267740 183592
rect 267695 183552 267740 183580
rect 267734 183540 267740 183552
rect 267792 183540 267798 183592
rect 270678 183580 270684 183592
rect 270639 183552 270684 183580
rect 270678 183540 270684 183552
rect 270736 183540 270742 183592
rect 284754 183540 284760 183592
rect 284812 183540 284818 183592
rect 294230 183540 294236 183592
rect 294288 183580 294294 183592
rect 294414 183580 294420 183592
rect 294288 183552 294420 183580
rect 294288 183540 294294 183552
rect 294414 183540 294420 183552
rect 294472 183540 294478 183592
rect 310882 183540 310888 183592
rect 310940 183580 310946 183592
rect 311066 183580 311072 183592
rect 310940 183552 311072 183580
rect 310940 183540 310946 183552
rect 311066 183540 311072 183552
rect 311124 183540 311130 183592
rect 339773 183583 339831 183589
rect 339773 183549 339785 183583
rect 339819 183580 339831 183583
rect 339862 183580 339868 183592
rect 339819 183552 339868 183580
rect 339819 183549 339831 183552
rect 339773 183543 339831 183549
rect 339862 183540 339868 183552
rect 339920 183540 339926 183592
rect 367002 183580 367008 183592
rect 366963 183552 367008 183580
rect 367002 183540 367008 183552
rect 367060 183540 367066 183592
rect 389266 183540 389272 183592
rect 389324 183580 389330 183592
rect 389542 183580 389548 183592
rect 389324 183552 389548 183580
rect 389324 183540 389330 183552
rect 389542 183540 389548 183552
rect 389600 183540 389606 183592
rect 463786 183540 463792 183592
rect 463844 183580 463850 183592
rect 464062 183580 464068 183592
rect 463844 183552 464068 183580
rect 463844 183540 463850 183552
rect 464062 183540 464068 183552
rect 464120 183540 464126 183592
rect 470410 183540 470416 183592
rect 470468 183580 470474 183592
rect 470594 183580 470600 183592
rect 470468 183552 470600 183580
rect 470468 183540 470474 183552
rect 470594 183540 470600 183552
rect 470652 183540 470658 183592
rect 273530 183472 273536 183524
rect 273588 183512 273594 183524
rect 273622 183512 273628 183524
rect 273588 183484 273628 183512
rect 273588 183472 273594 183484
rect 273622 183472 273628 183484
rect 273680 183472 273686 183524
rect 284772 183456 284800 183540
rect 284754 183404 284760 183456
rect 284812 183404 284818 183456
rect 232314 182152 232320 182164
rect 232275 182124 232320 182152
rect 232314 182112 232320 182124
rect 232372 182112 232378 182164
rect 301038 182112 301044 182164
rect 301096 182152 301102 182164
rect 301222 182152 301228 182164
rect 301096 182124 301228 182152
rect 301096 182112 301102 182124
rect 301222 182112 301228 182124
rect 301280 182112 301286 182164
rect 324498 182112 324504 182164
rect 324556 182152 324562 182164
rect 324556 182124 324728 182152
rect 324556 182112 324562 182124
rect 324700 182096 324728 182124
rect 326062 182112 326068 182164
rect 326120 182152 326126 182164
rect 326246 182152 326252 182164
rect 326120 182124 326252 182152
rect 326120 182112 326126 182124
rect 326246 182112 326252 182124
rect 326304 182112 326310 182164
rect 324682 182044 324688 182096
rect 324740 182044 324746 182096
rect 358722 182016 358728 182028
rect 358683 181988 358728 182016
rect 358722 181976 358728 181988
rect 358780 181976 358786 182028
rect 299842 180860 299848 180872
rect 299803 180832 299848 180860
rect 299842 180820 299848 180832
rect 299900 180820 299906 180872
rect 302510 180860 302516 180872
rect 302471 180832 302516 180860
rect 302510 180820 302516 180832
rect 302568 180820 302574 180872
rect 306834 180860 306840 180872
rect 306795 180832 306840 180860
rect 306834 180820 306840 180832
rect 306892 180820 306898 180872
rect 265158 180752 265164 180804
rect 265216 180792 265222 180804
rect 265250 180792 265256 180804
rect 265216 180764 265256 180792
rect 265216 180752 265222 180764
rect 265250 180752 265256 180764
rect 265308 180752 265314 180804
rect 272242 180752 272248 180804
rect 272300 180792 272306 180804
rect 272426 180792 272432 180804
rect 272300 180764 272432 180792
rect 272300 180752 272306 180764
rect 272426 180752 272432 180764
rect 272484 180752 272490 180804
rect 284754 180792 284760 180804
rect 284715 180764 284760 180792
rect 284754 180752 284760 180764
rect 284812 180752 284818 180804
rect 317506 180752 317512 180804
rect 317564 180792 317570 180804
rect 317690 180792 317696 180804
rect 317564 180764 317696 180792
rect 317564 180752 317570 180764
rect 317690 180752 317696 180764
rect 317748 180752 317754 180804
rect 259638 179568 259644 179580
rect 259599 179540 259644 179568
rect 259638 179528 259644 179540
rect 259696 179528 259702 179580
rect 288713 179435 288771 179441
rect 288713 179401 288725 179435
rect 288759 179432 288771 179435
rect 288894 179432 288900 179444
rect 288759 179404 288900 179432
rect 288759 179401 288771 179404
rect 288713 179395 288771 179401
rect 288894 179392 288900 179404
rect 288952 179392 288958 179444
rect 265250 179364 265256 179376
rect 265211 179336 265256 179364
rect 265250 179324 265256 179336
rect 265308 179324 265314 179376
rect 341242 179364 341248 179376
rect 341203 179336 341248 179364
rect 341242 179324 341248 179336
rect 341300 179324 341306 179376
rect 294230 178712 294236 178764
rect 294288 178752 294294 178764
rect 294414 178752 294420 178764
rect 294288 178724 294420 178752
rect 294288 178712 294294 178724
rect 294414 178712 294420 178724
rect 294472 178712 294478 178764
rect 295518 178712 295524 178764
rect 295576 178752 295582 178764
rect 295702 178752 295708 178764
rect 295576 178724 295708 178752
rect 295576 178712 295582 178724
rect 295702 178712 295708 178724
rect 295760 178712 295766 178764
rect 296806 178712 296812 178764
rect 296864 178752 296870 178764
rect 296990 178752 296996 178764
rect 296864 178724 296996 178752
rect 296864 178712 296870 178724
rect 296990 178712 296996 178724
rect 297048 178712 297054 178764
rect 250070 177284 250076 177336
rect 250128 177324 250134 177336
rect 250346 177324 250352 177336
rect 250128 177296 250352 177324
rect 250128 177284 250134 177296
rect 250346 177284 250352 177296
rect 250404 177284 250410 177336
rect 310882 176780 310888 176792
rect 310808 176752 310888 176780
rect 310808 176656 310836 176752
rect 310882 176740 310888 176752
rect 310940 176740 310946 176792
rect 389542 176780 389548 176792
rect 389468 176752 389548 176780
rect 389468 176656 389496 176752
rect 389542 176740 389548 176752
rect 389600 176740 389606 176792
rect 463878 176672 463884 176724
rect 463936 176712 463942 176724
rect 464062 176712 464068 176724
rect 463936 176684 464068 176712
rect 463936 176672 463942 176684
rect 464062 176672 464068 176684
rect 464120 176672 464126 176724
rect 310790 176604 310796 176656
rect 310848 176604 310854 176656
rect 338850 176604 338856 176656
rect 338908 176604 338914 176656
rect 374362 176604 374368 176656
rect 374420 176604 374426 176656
rect 375834 176604 375840 176656
rect 375892 176604 375898 176656
rect 389450 176604 389456 176656
rect 389508 176604 389514 176656
rect 338868 176520 338896 176604
rect 374380 176520 374408 176604
rect 375852 176520 375880 176604
rect 338850 176468 338856 176520
rect 338908 176468 338914 176520
rect 374362 176468 374368 176520
rect 374420 176468 374426 176520
rect 375834 176468 375840 176520
rect 375892 176468 375898 176520
rect 366910 174060 366916 174072
rect 366871 174032 366916 174060
rect 366910 174020 366916 174032
rect 366968 174020 366974 174072
rect 259641 173995 259699 174001
rect 259641 173961 259653 173995
rect 259687 173992 259699 173995
rect 259730 173992 259736 174004
rect 259687 173964 259736 173992
rect 259687 173961 259699 173964
rect 259641 173955 259699 173961
rect 259730 173952 259736 173964
rect 259788 173952 259794 174004
rect 366818 173952 366824 174004
rect 366876 173992 366882 174004
rect 367002 173992 367008 174004
rect 366876 173964 367008 173992
rect 366876 173952 366882 173964
rect 367002 173952 367008 173964
rect 367060 173952 367066 174004
rect 230842 173884 230848 173936
rect 230900 173924 230906 173936
rect 231026 173924 231032 173936
rect 230900 173896 231032 173924
rect 230900 173884 230906 173896
rect 231026 173884 231032 173896
rect 231084 173884 231090 173936
rect 235074 173884 235080 173936
rect 235132 173924 235138 173936
rect 235166 173924 235172 173936
rect 235132 173896 235172 173924
rect 235132 173884 235138 173896
rect 235166 173884 235172 173896
rect 235224 173884 235230 173936
rect 236362 173884 236368 173936
rect 236420 173924 236426 173936
rect 236454 173924 236460 173936
rect 236420 173896 236460 173924
rect 236420 173884 236426 173896
rect 236454 173884 236460 173896
rect 236512 173884 236518 173936
rect 239122 173884 239128 173936
rect 239180 173924 239186 173936
rect 239214 173924 239220 173936
rect 239180 173896 239220 173924
rect 239180 173884 239186 173896
rect 239214 173884 239220 173896
rect 239272 173884 239278 173936
rect 251450 173884 251456 173936
rect 251508 173924 251514 173936
rect 251634 173924 251640 173936
rect 251508 173896 251640 173924
rect 251508 173884 251514 173896
rect 251634 173884 251640 173896
rect 251692 173884 251698 173936
rect 266630 173884 266636 173936
rect 266688 173924 266694 173936
rect 266814 173924 266820 173936
rect 266688 173896 266820 173924
rect 266688 173884 266694 173896
rect 266814 173884 266820 173896
rect 266872 173884 266878 173936
rect 323302 173884 323308 173936
rect 323360 173924 323366 173936
rect 323486 173924 323492 173936
rect 323360 173896 323492 173924
rect 323360 173884 323366 173896
rect 323486 173884 323492 173896
rect 323544 173884 323550 173936
rect 327166 173884 327172 173936
rect 327224 173924 327230 173936
rect 327258 173924 327264 173936
rect 327224 173896 327264 173924
rect 327224 173884 327230 173896
rect 327258 173884 327264 173896
rect 327316 173884 327322 173936
rect 331398 173884 331404 173936
rect 331456 173924 331462 173936
rect 331582 173924 331588 173936
rect 331456 173896 331588 173924
rect 331456 173884 331462 173896
rect 331582 173884 331588 173896
rect 331640 173884 331646 173936
rect 337102 173884 337108 173936
rect 337160 173924 337166 173936
rect 337378 173924 337384 173936
rect 337160 173896 337384 173924
rect 337160 173884 337166 173896
rect 337378 173884 337384 173896
rect 337436 173884 337442 173936
rect 339678 173884 339684 173936
rect 339736 173924 339742 173936
rect 339862 173924 339868 173936
rect 339736 173896 339868 173924
rect 339736 173884 339742 173896
rect 339862 173884 339868 173896
rect 339920 173884 339926 173936
rect 357618 173884 357624 173936
rect 357676 173924 357682 173936
rect 357894 173924 357900 173936
rect 357676 173896 357900 173924
rect 357676 173884 357682 173896
rect 357894 173884 357900 173896
rect 357952 173884 357958 173936
rect 360470 173884 360476 173936
rect 360528 173924 360534 173936
rect 360562 173924 360568 173936
rect 360528 173896 360568 173924
rect 360528 173884 360534 173896
rect 360562 173884 360568 173896
rect 360620 173884 360626 173936
rect 366910 173924 366916 173936
rect 366871 173896 366916 173924
rect 366910 173884 366916 173896
rect 366968 173884 366974 173936
rect 372522 173884 372528 173936
rect 372580 173924 372586 173936
rect 372798 173924 372804 173936
rect 372580 173896 372804 173924
rect 372580 173884 372586 173896
rect 372798 173884 372804 173896
rect 372856 173884 372862 173936
rect 376938 173884 376944 173936
rect 376996 173924 377002 173936
rect 377122 173924 377128 173936
rect 376996 173896 377128 173924
rect 376996 173884 377002 173896
rect 377122 173884 377128 173896
rect 377180 173884 377186 173936
rect 358725 173859 358783 173865
rect 358725 173825 358737 173859
rect 358771 173856 358783 173859
rect 358814 173856 358820 173868
rect 358771 173828 358820 173856
rect 358771 173825 358783 173828
rect 358725 173819 358783 173825
rect 358814 173816 358820 173828
rect 358872 173816 358878 173868
rect 232314 172564 232320 172576
rect 232275 172536 232320 172564
rect 232314 172524 232320 172536
rect 232372 172524 232378 172576
rect 232222 172496 232228 172508
rect 232183 172468 232228 172496
rect 232222 172456 232228 172468
rect 232280 172456 232286 172508
rect 270494 172456 270500 172508
rect 270552 172496 270558 172508
rect 270770 172496 270776 172508
rect 270552 172468 270776 172496
rect 270552 172456 270558 172468
rect 270770 172456 270776 172468
rect 270828 172456 270834 172508
rect 301038 172456 301044 172508
rect 301096 172496 301102 172508
rect 301130 172496 301136 172508
rect 301096 172468 301136 172496
rect 301096 172456 301102 172468
rect 301130 172456 301136 172468
rect 301188 172456 301194 172508
rect 330110 172456 330116 172508
rect 330168 172496 330174 172508
rect 330294 172496 330300 172508
rect 330168 172468 330300 172496
rect 330168 172456 330174 172468
rect 330294 172456 330300 172468
rect 330352 172456 330358 172508
rect 337102 172496 337108 172508
rect 337063 172468 337108 172496
rect 337102 172456 337108 172468
rect 337160 172456 337166 172508
rect 284757 171139 284815 171145
rect 284757 171105 284769 171139
rect 284803 171136 284815 171139
rect 284938 171136 284944 171148
rect 284803 171108 284944 171136
rect 284803 171105 284815 171108
rect 284757 171099 284815 171105
rect 284938 171096 284944 171108
rect 284996 171096 285002 171148
rect 267826 171068 267832 171080
rect 267787 171040 267832 171068
rect 267826 171028 267832 171040
rect 267884 171028 267890 171080
rect 294414 171068 294420 171080
rect 294375 171040 294420 171068
rect 294414 171028 294420 171040
rect 294472 171028 294478 171080
rect 306834 171028 306840 171080
rect 306892 171068 306898 171080
rect 307018 171068 307024 171080
rect 306892 171040 307024 171068
rect 306892 171028 306898 171040
rect 307018 171028 307024 171040
rect 307076 171028 307082 171080
rect 341242 169776 341248 169788
rect 341203 169748 341248 169776
rect 341242 169736 341248 169748
rect 341300 169736 341306 169788
rect 259730 169056 259736 169108
rect 259788 169096 259794 169108
rect 259914 169096 259920 169108
rect 259788 169068 259920 169096
rect 259788 169056 259794 169068
rect 259914 169056 259920 169068
rect 259972 169056 259978 169108
rect 310790 167016 310796 167068
rect 310848 167016 310854 167068
rect 310808 166920 310836 167016
rect 310882 166920 310888 166932
rect 310808 166892 310888 166920
rect 310882 166880 310888 166892
rect 310940 166880 310946 166932
rect 2774 165452 2780 165504
rect 2832 165492 2838 165504
rect 5258 165492 5264 165504
rect 2832 165464 5264 165492
rect 2832 165452 2838 165464
rect 5258 165452 5264 165464
rect 5316 165452 5322 165504
rect 358722 164228 358728 164280
rect 358780 164268 358786 164280
rect 358814 164268 358820 164280
rect 358780 164240 358820 164268
rect 358780 164228 358786 164240
rect 358814 164228 358820 164240
rect 358872 164228 358878 164280
rect 232222 164200 232228 164212
rect 232183 164172 232228 164200
rect 232222 164160 232228 164172
rect 232280 164160 232286 164212
rect 244274 164160 244280 164212
rect 244332 164200 244338 164212
rect 244458 164200 244464 164212
rect 244332 164172 244464 164200
rect 244332 164160 244338 164172
rect 244458 164160 244464 164172
rect 244516 164160 244522 164212
rect 251450 164160 251456 164212
rect 251508 164200 251514 164212
rect 251634 164200 251640 164212
rect 251508 164172 251640 164200
rect 251508 164160 251514 164172
rect 251634 164160 251640 164172
rect 251692 164160 251698 164212
rect 259638 164160 259644 164212
rect 259696 164200 259702 164212
rect 259822 164200 259828 164212
rect 259696 164172 259828 164200
rect 259696 164160 259702 164172
rect 259822 164160 259828 164172
rect 259880 164160 259886 164212
rect 295518 164160 295524 164212
rect 295576 164200 295582 164212
rect 295702 164200 295708 164212
rect 295576 164172 295708 164200
rect 295576 164160 295582 164172
rect 295702 164160 295708 164172
rect 295760 164160 295766 164212
rect 337102 164200 337108 164212
rect 337063 164172 337108 164200
rect 337102 164160 337108 164172
rect 337160 164160 337166 164212
rect 372798 164200 372804 164212
rect 372759 164172 372804 164200
rect 372798 164160 372804 164172
rect 372856 164160 372862 164212
rect 376938 164160 376944 164212
rect 376996 164200 377002 164212
rect 377122 164200 377128 164212
rect 376996 164172 377128 164200
rect 376996 164160 377002 164172
rect 377122 164160 377128 164172
rect 377180 164160 377186 164212
rect 463786 164160 463792 164212
rect 463844 164200 463850 164212
rect 464062 164200 464068 164212
rect 463844 164172 464068 164200
rect 463844 164160 463850 164172
rect 464062 164160 464068 164172
rect 464120 164160 464126 164212
rect 284754 162868 284760 162920
rect 284812 162908 284818 162920
rect 284938 162908 284944 162920
rect 284812 162880 284944 162908
rect 284812 162868 284818 162880
rect 284938 162868 284944 162880
rect 284996 162868 285002 162920
rect 285766 162800 285772 162852
rect 285824 162840 285830 162852
rect 285950 162840 285956 162852
rect 285824 162812 285956 162840
rect 285824 162800 285830 162812
rect 285950 162800 285956 162812
rect 286008 162800 286014 162852
rect 325878 162800 325884 162852
rect 325936 162840 325942 162852
rect 326154 162840 326160 162852
rect 325936 162812 326160 162840
rect 325936 162800 325942 162812
rect 326154 162800 326160 162812
rect 326212 162800 326218 162852
rect 329926 162800 329932 162852
rect 329984 162840 329990 162852
rect 330110 162840 330116 162852
rect 329984 162812 330116 162840
rect 329984 162800 329990 162812
rect 330110 162800 330116 162812
rect 330168 162800 330174 162852
rect 357526 162800 357532 162852
rect 357584 162840 357590 162852
rect 357802 162840 357808 162852
rect 357584 162812 357808 162840
rect 357584 162800 357590 162812
rect 357802 162800 357808 162812
rect 357860 162800 357866 162852
rect 358722 162840 358728 162852
rect 358683 162812 358728 162840
rect 358722 162800 358728 162812
rect 358780 162800 358786 162852
rect 267826 162772 267832 162784
rect 267787 162744 267832 162772
rect 267826 162732 267832 162744
rect 267884 162732 267890 162784
rect 288894 161548 288900 161560
rect 288820 161520 288900 161548
rect 262582 161440 262588 161492
rect 262640 161480 262646 161492
rect 262674 161480 262680 161492
rect 262640 161452 262680 161480
rect 262640 161440 262646 161452
rect 262674 161440 262680 161452
rect 262732 161440 262738 161492
rect 265253 161483 265311 161489
rect 265253 161449 265265 161483
rect 265299 161480 265311 161483
rect 265342 161480 265348 161492
rect 265299 161452 265348 161480
rect 265299 161449 265311 161452
rect 265253 161443 265311 161449
rect 265342 161440 265348 161452
rect 265400 161440 265406 161492
rect 288820 161424 288848 161520
rect 288894 161508 288900 161520
rect 288952 161508 288958 161560
rect 289998 161508 290004 161560
rect 290056 161508 290062 161560
rect 290016 161480 290044 161508
rect 290090 161480 290096 161492
rect 290016 161452 290096 161480
rect 290090 161440 290096 161452
rect 290148 161440 290154 161492
rect 294414 161480 294420 161492
rect 294375 161452 294420 161480
rect 294414 161440 294420 161452
rect 294472 161440 294478 161492
rect 296990 161440 296996 161492
rect 297048 161480 297054 161492
rect 297082 161480 297088 161492
rect 297048 161452 297088 161480
rect 297048 161440 297054 161452
rect 297082 161440 297088 161452
rect 297140 161440 297146 161492
rect 302510 161440 302516 161492
rect 302568 161480 302574 161492
rect 302602 161480 302608 161492
rect 302568 161452 302608 161480
rect 302568 161440 302574 161452
rect 302602 161440 302608 161452
rect 302660 161440 302666 161492
rect 267826 161412 267832 161424
rect 267787 161384 267832 161412
rect 267826 161372 267832 161384
rect 267884 161372 267890 161424
rect 288802 161372 288808 161424
rect 288860 161372 288866 161424
rect 306834 161412 306840 161424
rect 306795 161384 306840 161412
rect 306834 161372 306840 161384
rect 306892 161372 306898 161424
rect 291378 161304 291384 161356
rect 291436 161344 291442 161356
rect 291562 161344 291568 161356
rect 291436 161316 291568 161344
rect 291436 161304 291442 161316
rect 291562 161304 291568 161316
rect 291620 161304 291626 161356
rect 288710 160012 288716 160064
rect 288768 160052 288774 160064
rect 288802 160052 288808 160064
rect 288768 160024 288808 160052
rect 288768 160012 288774 160024
rect 288802 160012 288808 160024
rect 288860 160012 288866 160064
rect 291473 160055 291531 160061
rect 291473 160021 291485 160055
rect 291519 160052 291531 160055
rect 291562 160052 291568 160064
rect 291519 160024 291568 160052
rect 291519 160021 291531 160024
rect 291473 160015 291531 160021
rect 291562 160012 291568 160024
rect 291620 160012 291626 160064
rect 294414 160052 294420 160064
rect 294375 160024 294420 160052
rect 294414 160012 294420 160024
rect 294472 160012 294478 160064
rect 341242 160052 341248 160064
rect 341203 160024 341248 160052
rect 341242 160012 341248 160024
rect 341300 160012 341306 160064
rect 372798 159304 372804 159316
rect 372759 159276 372804 159304
rect 372798 159264 372804 159276
rect 372856 159264 372862 159316
rect 417878 157496 417884 157548
rect 417936 157536 417942 157548
rect 418154 157536 418160 157548
rect 417936 157508 418160 157536
rect 417936 157496 417942 157508
rect 418154 157496 418160 157508
rect 418212 157496 418218 157548
rect 437198 157496 437204 157548
rect 437256 157536 437262 157548
rect 437474 157536 437480 157548
rect 437256 157508 437480 157536
rect 437256 157496 437262 157508
rect 437474 157496 437480 157508
rect 437532 157496 437538 157548
rect 456518 157496 456524 157548
rect 456576 157536 456582 157548
rect 456886 157536 456892 157548
rect 456576 157508 456892 157536
rect 456576 157496 456582 157508
rect 456886 157496 456892 157508
rect 456944 157496 456950 157548
rect 306282 157428 306288 157480
rect 306340 157468 306346 157480
rect 314562 157468 314568 157480
rect 306340 157440 314568 157468
rect 306340 157428 306346 157440
rect 314562 157428 314568 157440
rect 314620 157428 314626 157480
rect 230750 157360 230756 157412
rect 230808 157360 230814 157412
rect 282638 157360 282644 157412
rect 282696 157400 282702 157412
rect 288894 157400 288900 157412
rect 282696 157372 288900 157400
rect 282696 157360 282702 157372
rect 288894 157360 288900 157372
rect 288952 157360 288958 157412
rect 327166 157360 327172 157412
rect 327224 157360 327230 157412
rect 230768 157332 230796 157360
rect 230842 157332 230848 157344
rect 230768 157304 230848 157332
rect 230842 157292 230848 157304
rect 230900 157292 230906 157344
rect 327184 157264 327212 157360
rect 374362 157292 374368 157344
rect 374420 157292 374426 157344
rect 375834 157292 375840 157344
rect 375892 157292 375898 157344
rect 327258 157264 327264 157276
rect 327184 157236 327264 157264
rect 327258 157224 327264 157236
rect 327316 157224 327322 157276
rect 374380 157208 374408 157292
rect 375852 157208 375880 157292
rect 374362 157156 374368 157208
rect 374420 157156 374426 157208
rect 375834 157156 375840 157208
rect 375892 157156 375898 157208
rect 339586 154640 339592 154692
rect 339644 154640 339650 154692
rect 247218 154572 247224 154624
rect 247276 154612 247282 154624
rect 247310 154612 247316 154624
rect 247276 154584 247316 154612
rect 247276 154572 247282 154584
rect 247310 154572 247316 154584
rect 247368 154572 247374 154624
rect 339604 154556 339632 154640
rect 302510 154504 302516 154556
rect 302568 154544 302574 154556
rect 302602 154544 302608 154556
rect 302568 154516 302608 154544
rect 302568 154504 302574 154516
rect 302602 154504 302608 154516
rect 302660 154504 302666 154556
rect 337194 154544 337200 154556
rect 337155 154516 337200 154544
rect 337194 154504 337200 154516
rect 337252 154504 337258 154556
rect 339586 154504 339592 154556
rect 339644 154504 339650 154556
rect 358722 154544 358728 154556
rect 358683 154516 358728 154544
rect 358722 154504 358728 154516
rect 358780 154504 358786 154556
rect 367002 154544 367008 154556
rect 366963 154516 367008 154544
rect 367002 154504 367008 154516
rect 367060 154504 367066 154556
rect 389450 154504 389456 154556
rect 389508 154544 389514 154556
rect 389634 154544 389640 154556
rect 389508 154516 389640 154544
rect 389508 154504 389514 154516
rect 389634 154504 389640 154516
rect 389692 154504 389698 154556
rect 470410 154504 470416 154556
rect 470468 154544 470474 154556
rect 470594 154544 470600 154556
rect 470468 154516 470600 154544
rect 470468 154504 470474 154516
rect 470594 154504 470600 154516
rect 470652 154504 470658 154556
rect 259641 154207 259699 154213
rect 259641 154173 259653 154207
rect 259687 154204 259699 154207
rect 259822 154204 259828 154216
rect 259687 154176 259828 154204
rect 259687 154173 259699 154176
rect 259641 154167 259699 154173
rect 259822 154164 259828 154176
rect 259880 154164 259886 154216
rect 272150 153212 272156 153264
rect 272208 153252 272214 153264
rect 272242 153252 272248 153264
rect 272208 153224 272248 153252
rect 272208 153212 272214 153224
rect 272242 153212 272248 153224
rect 272300 153212 272306 153264
rect 285950 153144 285956 153196
rect 286008 153184 286014 153196
rect 286042 153184 286048 153196
rect 286008 153156 286048 153184
rect 286008 153144 286014 153156
rect 286042 153144 286048 153156
rect 286100 153144 286106 153196
rect 302418 153144 302424 153196
rect 302476 153184 302482 153196
rect 302510 153184 302516 153196
rect 302476 153156 302516 153184
rect 302476 153144 302482 153156
rect 302510 153144 302516 153156
rect 302568 153144 302574 153196
rect 310790 153184 310796 153196
rect 310751 153156 310796 153184
rect 310790 153144 310796 153156
rect 310848 153144 310854 153196
rect 375834 153184 375840 153196
rect 375795 153156 375840 153184
rect 375834 153144 375840 153156
rect 375892 153144 375898 153196
rect 264974 153076 264980 153128
rect 265032 153116 265038 153128
rect 265342 153116 265348 153128
rect 265032 153088 265348 153116
rect 265032 153076 265038 153088
rect 265342 153076 265348 153088
rect 265400 153076 265406 153128
rect 337197 152371 337255 152377
rect 337197 152337 337209 152371
rect 337243 152368 337255 152371
rect 337286 152368 337292 152380
rect 337243 152340 337292 152368
rect 337243 152337 337255 152340
rect 337197 152331 337255 152337
rect 337286 152328 337292 152340
rect 337344 152328 337350 152380
rect 267826 151824 267832 151836
rect 267787 151796 267832 151824
rect 267826 151784 267832 151796
rect 267884 151784 267890 151836
rect 296898 151784 296904 151836
rect 296956 151824 296962 151836
rect 297082 151824 297088 151836
rect 296956 151796 297088 151824
rect 296956 151784 296962 151796
rect 297082 151784 297088 151796
rect 297140 151784 297146 151836
rect 306837 151827 306895 151833
rect 306837 151793 306849 151827
rect 306883 151824 306895 151827
rect 306926 151824 306932 151836
rect 306883 151796 306932 151824
rect 306883 151793 306895 151796
rect 306837 151787 306895 151793
rect 306926 151784 306932 151796
rect 306984 151784 306990 151836
rect 3326 151716 3332 151768
rect 3384 151756 3390 151768
rect 17218 151756 17224 151768
rect 3384 151728 17224 151756
rect 3384 151716 3390 151728
rect 17218 151716 17224 151728
rect 17276 151716 17282 151768
rect 264974 151756 264980 151768
rect 264935 151728 264980 151756
rect 264974 151716 264980 151728
rect 265032 151716 265038 151768
rect 339773 151759 339831 151765
rect 339773 151725 339785 151759
rect 339819 151756 339831 151759
rect 339862 151756 339868 151768
rect 339819 151728 339868 151756
rect 339819 151725 339831 151728
rect 339773 151719 339831 151725
rect 339862 151716 339868 151728
rect 339920 151716 339926 151768
rect 294417 150467 294475 150473
rect 294417 150433 294429 150467
rect 294463 150464 294475 150467
rect 294506 150464 294512 150476
rect 294463 150436 294512 150464
rect 294463 150433 294475 150436
rect 294417 150427 294475 150433
rect 294506 150424 294512 150436
rect 294564 150424 294570 150476
rect 294233 150331 294291 150337
rect 294233 150297 294245 150331
rect 294279 150328 294291 150331
rect 294506 150328 294512 150340
rect 294279 150300 294512 150328
rect 294279 150297 294291 150300
rect 294233 150291 294291 150297
rect 294506 150288 294512 150300
rect 294564 150288 294570 150340
rect 291470 149104 291476 149116
rect 291431 149076 291476 149104
rect 291470 149064 291476 149076
rect 291528 149064 291534 149116
rect 338850 147636 338856 147688
rect 338908 147636 338914 147688
rect 310790 147608 310796 147620
rect 310751 147580 310796 147608
rect 310790 147568 310796 147580
rect 310848 147568 310854 147620
rect 338868 147608 338896 147636
rect 338942 147608 338948 147620
rect 338868 147580 338948 147608
rect 338942 147568 338948 147580
rect 339000 147568 339006 147620
rect 259638 145024 259644 145036
rect 259599 144996 259644 145024
rect 259638 144984 259644 144996
rect 259696 144984 259702 145036
rect 357526 144916 357532 144968
rect 357584 144956 357590 144968
rect 357802 144956 357808 144968
rect 357584 144928 357808 144956
rect 357584 144916 357590 144928
rect 357802 144916 357808 144928
rect 357860 144916 357866 144968
rect 358722 144916 358728 144968
rect 358780 144956 358786 144968
rect 358814 144956 358820 144968
rect 358780 144928 358820 144956
rect 358780 144916 358786 144928
rect 358814 144916 358820 144928
rect 358872 144916 358878 144968
rect 367002 144956 367008 144968
rect 366963 144928 367008 144956
rect 367002 144916 367008 144928
rect 367060 144916 367066 144968
rect 235994 144848 236000 144900
rect 236052 144888 236058 144900
rect 236270 144888 236276 144900
rect 236052 144860 236276 144888
rect 236052 144848 236058 144860
rect 236270 144848 236276 144860
rect 236328 144848 236334 144900
rect 244274 144848 244280 144900
rect 244332 144888 244338 144900
rect 244458 144888 244464 144900
rect 244332 144860 244464 144888
rect 244332 144848 244338 144860
rect 244458 144848 244464 144860
rect 244516 144848 244522 144900
rect 247126 144848 247132 144900
rect 247184 144888 247190 144900
rect 247218 144888 247224 144900
rect 247184 144860 247224 144888
rect 247184 144848 247190 144860
rect 247218 144848 247224 144860
rect 247276 144848 247282 144900
rect 270678 144888 270684 144900
rect 270639 144860 270684 144888
rect 270678 144848 270684 144860
rect 270736 144848 270742 144900
rect 272150 144848 272156 144900
rect 272208 144888 272214 144900
rect 272242 144888 272248 144900
rect 272208 144860 272248 144888
rect 272208 144848 272214 144860
rect 272242 144848 272248 144860
rect 272300 144848 272306 144900
rect 323302 144848 323308 144900
rect 323360 144888 323366 144900
rect 323394 144888 323400 144900
rect 323360 144860 323400 144888
rect 323360 144848 323366 144860
rect 323394 144848 323400 144860
rect 323452 144848 323458 144900
rect 324590 144848 324596 144900
rect 324648 144888 324654 144900
rect 324774 144888 324780 144900
rect 324648 144860 324780 144888
rect 324648 144848 324654 144860
rect 324774 144848 324780 144860
rect 324832 144848 324838 144900
rect 325878 144848 325884 144900
rect 325936 144848 325942 144900
rect 327166 144848 327172 144900
rect 327224 144888 327230 144900
rect 327350 144888 327356 144900
rect 327224 144860 327356 144888
rect 327224 144848 327230 144860
rect 327350 144848 327356 144860
rect 327408 144848 327414 144900
rect 376938 144848 376944 144900
rect 376996 144888 377002 144900
rect 377122 144888 377128 144900
rect 376996 144860 377128 144888
rect 376996 144848 377002 144860
rect 377122 144848 377128 144860
rect 377180 144848 377186 144900
rect 325896 144820 325924 144848
rect 325970 144820 325976 144832
rect 325896 144792 325976 144820
rect 325970 144780 325976 144792
rect 326028 144780 326034 144832
rect 265066 143556 265072 143608
rect 265124 143556 265130 143608
rect 375834 143596 375840 143608
rect 375795 143568 375840 143596
rect 375834 143556 375840 143568
rect 375892 143556 375898 143608
rect 250254 143528 250260 143540
rect 250215 143500 250260 143528
rect 250254 143488 250260 143500
rect 250312 143488 250318 143540
rect 262582 143488 262588 143540
rect 262640 143528 262646 143540
rect 262858 143528 262864 143540
rect 262640 143500 262864 143528
rect 262640 143488 262646 143500
rect 262858 143488 262864 143500
rect 262916 143488 262922 143540
rect 265084 143472 265112 143556
rect 323302 143488 323308 143540
rect 323360 143528 323366 143540
rect 323486 143528 323492 143540
rect 323360 143500 323492 143528
rect 323360 143488 323366 143500
rect 323486 143488 323492 143500
rect 323544 143488 323550 143540
rect 325970 143528 325976 143540
rect 325931 143500 325976 143528
rect 325970 143488 325976 143500
rect 326028 143488 326034 143540
rect 330110 143528 330116 143540
rect 330071 143500 330116 143528
rect 330110 143488 330116 143500
rect 330168 143488 330174 143540
rect 357250 143488 357256 143540
rect 357308 143528 357314 143540
rect 357526 143528 357532 143540
rect 357308 143500 357532 143528
rect 357308 143488 357314 143500
rect 357526 143488 357532 143500
rect 357584 143488 357590 143540
rect 358722 143528 358728 143540
rect 358683 143500 358728 143528
rect 358722 143488 358728 143500
rect 358780 143488 358786 143540
rect 360286 143528 360292 143540
rect 360247 143500 360292 143528
rect 360286 143488 360292 143500
rect 360344 143488 360350 143540
rect 265066 143420 265072 143472
rect 265124 143420 265130 143472
rect 341242 143392 341248 143404
rect 341203 143364 341248 143392
rect 341242 143352 341248 143364
rect 341300 143352 341306 143404
rect 264977 142171 265035 142177
rect 264977 142137 264989 142171
rect 265023 142168 265035 142171
rect 265250 142168 265256 142180
rect 265023 142140 265256 142168
rect 265023 142137 265035 142140
rect 264977 142131 265035 142137
rect 265250 142128 265256 142140
rect 265308 142128 265314 142180
rect 288618 142128 288624 142180
rect 288676 142168 288682 142180
rect 288802 142168 288808 142180
rect 288676 142140 288808 142168
rect 288676 142128 288682 142140
rect 288802 142128 288808 142140
rect 288860 142128 288866 142180
rect 290090 142128 290096 142180
rect 290148 142168 290154 142180
rect 290182 142168 290188 142180
rect 290148 142140 290188 142168
rect 290148 142128 290154 142140
rect 290182 142128 290188 142140
rect 290240 142128 290246 142180
rect 317506 142128 317512 142180
rect 317564 142168 317570 142180
rect 317690 142168 317696 142180
rect 317564 142140 317696 142168
rect 317564 142128 317570 142140
rect 317690 142128 317696 142140
rect 317748 142128 317754 142180
rect 339770 142168 339776 142180
rect 339731 142140 339776 142168
rect 339770 142128 339776 142140
rect 339828 142128 339834 142180
rect 296806 142100 296812 142112
rect 296767 142072 296812 142100
rect 296806 142060 296812 142072
rect 296864 142060 296870 142112
rect 301133 142103 301191 142109
rect 301133 142069 301145 142103
rect 301179 142100 301191 142103
rect 301222 142100 301228 142112
rect 301179 142072 301228 142100
rect 301179 142069 301191 142072
rect 301133 142063 301191 142069
rect 301222 142060 301228 142072
rect 301280 142060 301286 142112
rect 294230 140808 294236 140820
rect 294191 140780 294236 140808
rect 294230 140768 294236 140780
rect 294288 140768 294294 140820
rect 270678 139992 270684 140004
rect 270639 139964 270684 139992
rect 270678 139952 270684 139964
rect 270736 139952 270742 140004
rect 291470 139380 291476 139392
rect 291431 139352 291476 139380
rect 291470 139340 291476 139352
rect 291528 139340 291534 139392
rect 310793 138703 310851 138709
rect 310793 138669 310805 138703
rect 310839 138700 310851 138703
rect 310882 138700 310888 138712
rect 310839 138672 310888 138700
rect 310839 138669 310851 138672
rect 310793 138663 310851 138669
rect 310882 138660 310888 138672
rect 310940 138660 310946 138712
rect 330113 138703 330171 138709
rect 330113 138669 330125 138703
rect 330159 138700 330171 138703
rect 330202 138700 330208 138712
rect 330159 138672 330208 138700
rect 330159 138669 330171 138672
rect 330113 138663 330171 138669
rect 330202 138660 330208 138672
rect 330260 138660 330266 138712
rect 372709 138159 372767 138165
rect 372709 138125 372721 138159
rect 372755 138156 372767 138159
rect 372798 138156 372804 138168
rect 372755 138128 372804 138156
rect 372755 138125 372767 138128
rect 372709 138119 372767 138125
rect 372798 138116 372804 138128
rect 372856 138116 372862 138168
rect 239122 137980 239128 138032
rect 239180 137980 239186 138032
rect 338758 137980 338764 138032
rect 338816 138020 338822 138032
rect 338942 138020 338948 138032
rect 338816 137992 338948 138020
rect 338816 137980 338822 137992
rect 338942 137980 338948 137992
rect 339000 137980 339006 138032
rect 389358 137980 389364 138032
rect 389416 137980 389422 138032
rect 239140 137952 239168 137980
rect 239214 137952 239220 137964
rect 239140 137924 239220 137952
rect 239214 137912 239220 137924
rect 239272 137912 239278 137964
rect 317506 137912 317512 137964
rect 317564 137952 317570 137964
rect 317782 137952 317788 137964
rect 317564 137924 317788 137952
rect 317564 137912 317570 137924
rect 317782 137912 317788 137924
rect 317840 137912 317846 137964
rect 360289 137955 360347 137961
rect 360289 137921 360301 137955
rect 360335 137952 360347 137955
rect 360378 137952 360384 137964
rect 360335 137924 360384 137952
rect 360335 137921 360347 137924
rect 360289 137915 360347 137921
rect 360378 137912 360384 137924
rect 360436 137912 360442 137964
rect 389376 137952 389404 137980
rect 389450 137952 389456 137964
rect 389376 137924 389456 137952
rect 389450 137912 389456 137924
rect 389508 137912 389514 137964
rect 299750 137368 299756 137420
rect 299808 137408 299814 137420
rect 299934 137408 299940 137420
rect 299808 137380 299940 137408
rect 299808 137368 299814 137380
rect 299934 137368 299940 137380
rect 299992 137368 299998 137420
rect 306742 137368 306748 137420
rect 306800 137408 306806 137420
rect 306926 137408 306932 137420
rect 306800 137380 306932 137408
rect 306800 137368 306806 137380
rect 306926 137368 306932 137380
rect 306984 137368 306990 137420
rect 2774 136348 2780 136400
rect 2832 136388 2838 136400
rect 5166 136388 5172 136400
rect 2832 136360 5172 136388
rect 2832 136348 2838 136360
rect 5166 136348 5172 136360
rect 5224 136348 5230 136400
rect 372706 135300 372712 135312
rect 372667 135272 372712 135300
rect 372706 135260 372712 135272
rect 372764 135260 372770 135312
rect 302510 135192 302516 135244
rect 302568 135232 302574 135244
rect 302602 135232 302608 135244
rect 302568 135204 302608 135232
rect 302568 135192 302574 135204
rect 302602 135192 302608 135204
rect 302660 135192 302666 135244
rect 327169 135235 327227 135241
rect 327169 135201 327181 135235
rect 327215 135232 327227 135235
rect 327258 135232 327264 135244
rect 327215 135204 327264 135232
rect 327215 135201 327227 135204
rect 327169 135195 327227 135201
rect 327258 135192 327264 135204
rect 327316 135192 327322 135244
rect 358722 135232 358728 135244
rect 358683 135204 358728 135232
rect 358722 135192 358728 135204
rect 358780 135192 358786 135244
rect 470410 135192 470416 135244
rect 470468 135232 470474 135244
rect 470594 135232 470600 135244
rect 470468 135204 470600 135232
rect 470468 135192 470474 135204
rect 470594 135192 470600 135204
rect 470652 135192 470658 135244
rect 250257 133943 250315 133949
rect 250257 133909 250269 133943
rect 250303 133940 250315 133943
rect 250346 133940 250352 133952
rect 250303 133912 250352 133940
rect 250303 133909 250315 133912
rect 250257 133903 250315 133909
rect 250346 133900 250352 133912
rect 250404 133900 250410 133952
rect 302510 133872 302516 133884
rect 302471 133844 302516 133872
rect 302510 133832 302516 133844
rect 302568 133832 302574 133884
rect 306742 133872 306748 133884
rect 306703 133844 306748 133872
rect 306742 133832 306748 133844
rect 306800 133832 306806 133884
rect 337102 133872 337108 133884
rect 337063 133844 337108 133872
rect 337102 133832 337108 133844
rect 337160 133832 337166 133884
rect 375834 133872 375840 133884
rect 375795 133844 375840 133872
rect 375834 133832 375840 133844
rect 375892 133832 375898 133884
rect 389450 133872 389456 133884
rect 389411 133844 389456 133872
rect 389450 133832 389456 133844
rect 389508 133832 389514 133884
rect 289998 132472 290004 132524
rect 290056 132512 290062 132524
rect 290090 132512 290096 132524
rect 290056 132484 290096 132512
rect 290056 132472 290062 132484
rect 290090 132472 290096 132484
rect 290148 132472 290154 132524
rect 295518 132472 295524 132524
rect 295576 132512 295582 132524
rect 295610 132512 295616 132524
rect 295576 132484 295616 132512
rect 295576 132472 295582 132484
rect 295610 132472 295616 132484
rect 295668 132472 295674 132524
rect 296809 132515 296867 132521
rect 296809 132481 296821 132515
rect 296855 132512 296867 132515
rect 296898 132512 296904 132524
rect 296855 132484 296904 132512
rect 296855 132481 296867 132484
rect 296809 132475 296867 132481
rect 296898 132472 296904 132484
rect 296956 132472 296962 132524
rect 301130 132512 301136 132524
rect 301091 132484 301136 132512
rect 301130 132472 301136 132484
rect 301188 132472 301194 132524
rect 325970 132512 325976 132524
rect 325931 132484 325976 132512
rect 325970 132472 325976 132484
rect 326028 132472 326034 132524
rect 284662 132444 284668 132456
rect 284623 132416 284668 132444
rect 284662 132404 284668 132416
rect 284720 132404 284726 132456
rect 270494 130364 270500 130416
rect 270552 130404 270558 130416
rect 270678 130404 270684 130416
rect 270552 130376 270684 130404
rect 270552 130364 270558 130376
rect 270678 130364 270684 130376
rect 270736 130364 270742 130416
rect 272150 130364 272156 130416
rect 272208 130404 272214 130416
rect 272334 130404 272340 130416
rect 272208 130376 272340 130404
rect 272208 130364 272214 130376
rect 272334 130364 272340 130376
rect 272392 130364 272398 130416
rect 463878 130364 463884 130416
rect 463936 130404 463942 130416
rect 464062 130404 464068 130416
rect 463936 130376 464068 130404
rect 463936 130364 463942 130376
rect 464062 130364 464068 130376
rect 464120 130364 464126 130416
rect 327166 129724 327172 129736
rect 327127 129696 327172 129724
rect 327166 129684 327172 129696
rect 327224 129684 327230 129736
rect 259730 128324 259736 128376
rect 259788 128324 259794 128376
rect 259748 128296 259776 128324
rect 259822 128296 259828 128308
rect 259748 128268 259828 128296
rect 259822 128256 259828 128268
rect 259880 128256 259886 128308
rect 310790 128296 310796 128308
rect 310751 128268 310796 128296
rect 310790 128256 310796 128268
rect 310848 128256 310854 128308
rect 284662 126936 284668 126948
rect 284623 126908 284668 126936
rect 284662 126896 284668 126908
rect 284720 126896 284726 126948
rect 358722 125604 358728 125656
rect 358780 125644 358786 125656
rect 358814 125644 358820 125656
rect 358780 125616 358820 125644
rect 358780 125604 358786 125616
rect 358814 125604 358820 125616
rect 358872 125604 358878 125656
rect 251450 125576 251456 125588
rect 251411 125548 251456 125576
rect 251450 125536 251456 125548
rect 251508 125536 251514 125588
rect 265158 125536 265164 125588
rect 265216 125576 265222 125588
rect 265342 125576 265348 125588
rect 265216 125548 265348 125576
rect 265216 125536 265222 125548
rect 265342 125536 265348 125548
rect 265400 125536 265406 125588
rect 266538 125536 266544 125588
rect 266596 125576 266602 125588
rect 266722 125576 266728 125588
rect 266596 125548 266728 125576
rect 266596 125536 266602 125548
rect 266722 125536 266728 125548
rect 266780 125536 266786 125588
rect 267734 125536 267740 125588
rect 267792 125576 267798 125588
rect 267918 125576 267924 125588
rect 267792 125548 267924 125576
rect 267792 125536 267798 125548
rect 267918 125536 267924 125548
rect 267976 125536 267982 125588
rect 270678 125576 270684 125588
rect 270639 125548 270684 125576
rect 270678 125536 270684 125548
rect 270736 125536 270742 125588
rect 272150 125576 272156 125588
rect 272111 125548 272156 125576
rect 272150 125536 272156 125548
rect 272208 125536 272214 125588
rect 323210 125536 323216 125588
rect 323268 125576 323274 125588
rect 323394 125576 323400 125588
rect 323268 125548 323400 125576
rect 323268 125536 323274 125548
rect 323394 125536 323400 125548
rect 323452 125536 323458 125588
rect 324590 125536 324596 125588
rect 324648 125576 324654 125588
rect 324774 125576 324780 125588
rect 324648 125548 324780 125576
rect 324648 125536 324654 125548
rect 324774 125536 324780 125548
rect 324832 125536 324838 125588
rect 327166 125536 327172 125588
rect 327224 125576 327230 125588
rect 327350 125576 327356 125588
rect 327224 125548 327356 125576
rect 327224 125536 327230 125548
rect 327350 125536 327356 125548
rect 327408 125536 327414 125588
rect 367002 125576 367008 125588
rect 366963 125548 367008 125576
rect 367002 125536 367008 125548
rect 367060 125536 367066 125588
rect 372706 125576 372712 125588
rect 372667 125548 372712 125576
rect 372706 125536 372712 125548
rect 372764 125536 372770 125588
rect 259730 125468 259736 125520
rect 259788 125508 259794 125520
rect 259822 125508 259828 125520
rect 259788 125480 259828 125508
rect 259788 125468 259794 125480
rect 259822 125468 259828 125480
rect 259880 125468 259886 125520
rect 310793 125511 310851 125517
rect 310793 125477 310805 125511
rect 310839 125508 310851 125511
rect 310882 125508 310888 125520
rect 310839 125480 310888 125508
rect 310839 125477 310851 125480
rect 310793 125471 310851 125477
rect 310882 125468 310888 125480
rect 310940 125468 310946 125520
rect 302513 124219 302571 124225
rect 302513 124185 302525 124219
rect 302559 124216 302571 124219
rect 302602 124216 302608 124228
rect 302559 124188 302608 124216
rect 302559 124185 302571 124188
rect 302513 124179 302571 124185
rect 302602 124176 302608 124188
rect 302660 124176 302666 124228
rect 306745 124219 306803 124225
rect 306745 124185 306757 124219
rect 306791 124216 306803 124219
rect 306834 124216 306840 124228
rect 306791 124188 306840 124216
rect 306791 124185 306803 124188
rect 306745 124179 306803 124185
rect 306834 124176 306840 124188
rect 306892 124176 306898 124228
rect 330110 124176 330116 124228
rect 330168 124216 330174 124228
rect 330294 124216 330300 124228
rect 330168 124188 330300 124216
rect 330168 124176 330174 124188
rect 330294 124176 330300 124188
rect 330352 124176 330358 124228
rect 337105 124219 337163 124225
rect 337105 124185 337117 124219
rect 337151 124216 337163 124219
rect 337194 124216 337200 124228
rect 337151 124188 337200 124216
rect 337151 124185 337163 124188
rect 337105 124179 337163 124185
rect 337194 124176 337200 124188
rect 337252 124176 337258 124228
rect 375834 124216 375840 124228
rect 375795 124188 375840 124216
rect 375834 124176 375840 124188
rect 375892 124176 375898 124228
rect 300946 124108 300952 124160
rect 301004 124108 301010 124160
rect 358722 124148 358728 124160
rect 358683 124120 358728 124148
rect 358722 124108 358728 124120
rect 358780 124108 358786 124160
rect 300964 124024 300992 124108
rect 300946 123972 300952 124024
rect 301004 123972 301010 124024
rect 288802 122856 288808 122868
rect 288763 122828 288808 122856
rect 288802 122816 288808 122828
rect 288860 122816 288866 122868
rect 389174 122816 389180 122868
rect 389232 122856 389238 122868
rect 389453 122859 389511 122865
rect 389453 122856 389465 122859
rect 389232 122828 389465 122856
rect 389232 122816 389238 122828
rect 389453 122825 389465 122828
rect 389499 122825 389511 122859
rect 389453 122819 389511 122825
rect 235077 122791 235135 122797
rect 235077 122757 235089 122791
rect 235123 122788 235135 122791
rect 235166 122788 235172 122800
rect 235123 122760 235172 122788
rect 235123 122757 235135 122760
rect 235077 122751 235135 122757
rect 235166 122748 235172 122760
rect 235224 122748 235230 122800
rect 239125 122791 239183 122797
rect 239125 122757 239137 122791
rect 239171 122788 239183 122791
rect 239214 122788 239220 122800
rect 239171 122760 239220 122788
rect 239171 122757 239183 122760
rect 239125 122751 239183 122757
rect 239214 122748 239220 122760
rect 239272 122748 239278 122800
rect 284662 122748 284668 122800
rect 284720 122788 284726 122800
rect 284846 122788 284852 122800
rect 284720 122760 284852 122788
rect 284720 122748 284726 122760
rect 284846 122748 284852 122760
rect 284904 122748 284910 122800
rect 289998 122788 290004 122800
rect 289959 122760 290004 122788
rect 289998 122748 290004 122760
rect 290056 122748 290062 122800
rect 301130 122788 301136 122800
rect 301091 122760 301136 122788
rect 301130 122748 301136 122760
rect 301188 122748 301194 122800
rect 306653 122791 306711 122797
rect 306653 122757 306665 122791
rect 306699 122788 306711 122791
rect 306834 122788 306840 122800
rect 306699 122760 306840 122788
rect 306699 122757 306711 122760
rect 306653 122751 306711 122757
rect 306834 122748 306840 122760
rect 306892 122748 306898 122800
rect 330110 122788 330116 122800
rect 330071 122760 330116 122788
rect 330110 122748 330116 122760
rect 330168 122748 330174 122800
rect 337194 122788 337200 122800
rect 337155 122760 337200 122788
rect 337194 122748 337200 122760
rect 337252 122748 337258 122800
rect 296898 122720 296904 122732
rect 296859 122692 296904 122720
rect 296898 122680 296904 122692
rect 296956 122680 296962 122732
rect 2774 122340 2780 122392
rect 2832 122380 2838 122392
rect 5074 122380 5080 122392
rect 2832 122352 5080 122380
rect 2832 122340 2838 122352
rect 5074 122340 5080 122352
rect 5132 122340 5138 122392
rect 288802 121456 288808 121508
rect 288860 121496 288866 121508
rect 291473 121499 291531 121505
rect 288860 121468 288905 121496
rect 288860 121456 288866 121468
rect 291473 121465 291485 121499
rect 291519 121496 291531 121499
rect 291654 121496 291660 121508
rect 291519 121468 291660 121496
rect 291519 121465 291531 121468
rect 291473 121459 291531 121465
rect 291654 121456 291660 121468
rect 291712 121456 291718 121508
rect 295794 121388 295800 121440
rect 295852 121428 295858 121440
rect 295852 121400 295897 121428
rect 295852 121388 295858 121400
rect 244458 120708 244464 120760
rect 244516 120748 244522 120760
rect 244642 120748 244648 120760
rect 244516 120720 244648 120748
rect 244516 120708 244522 120720
rect 244642 120708 244648 120720
rect 244700 120708 244706 120760
rect 267826 120640 267832 120692
rect 267884 120680 267890 120692
rect 267918 120680 267924 120692
rect 267884 120652 267924 120680
rect 267884 120640 267890 120652
rect 267918 120640 267924 120652
rect 267976 120640 267982 120692
rect 270678 120680 270684 120692
rect 270639 120652 270684 120680
rect 270678 120640 270684 120652
rect 270736 120640 270742 120692
rect 272150 120680 272156 120692
rect 272111 120652 272156 120680
rect 272150 120640 272156 120652
rect 272208 120640 272214 120692
rect 273530 118736 273536 118788
rect 273588 118736 273594 118788
rect 357526 118776 357532 118788
rect 357452 118748 357532 118776
rect 273548 118652 273576 118736
rect 357452 118652 357480 118748
rect 357526 118736 357532 118748
rect 357584 118736 357590 118788
rect 360378 118668 360384 118720
rect 360436 118668 360442 118720
rect 377122 118668 377128 118720
rect 377180 118668 377186 118720
rect 463878 118668 463884 118720
rect 463936 118668 463942 118720
rect 273530 118600 273536 118652
rect 273588 118600 273594 118652
rect 357434 118600 357440 118652
rect 357492 118600 357498 118652
rect 360396 118640 360424 118668
rect 360470 118640 360476 118652
rect 360396 118612 360476 118640
rect 360470 118600 360476 118612
rect 360528 118600 360534 118652
rect 377140 118584 377168 118668
rect 463896 118640 463924 118668
rect 463970 118640 463976 118652
rect 463896 118612 463976 118640
rect 463970 118600 463976 118612
rect 464028 118600 464034 118652
rect 377122 118532 377128 118584
rect 377180 118532 377186 118584
rect 239122 118028 239128 118040
rect 239083 118000 239128 118028
rect 239122 117988 239128 118000
rect 239180 117988 239186 118040
rect 325881 118031 325939 118037
rect 325881 117997 325893 118031
rect 325927 118028 325939 118031
rect 325970 118028 325976 118040
rect 325927 118000 325976 118028
rect 325927 117997 325939 118000
rect 325881 117991 325939 117997
rect 325970 117988 325976 118000
rect 326028 117988 326034 118040
rect 337194 118028 337200 118040
rect 337155 118000 337200 118028
rect 337194 117988 337200 118000
rect 337252 117988 337258 118040
rect 310790 116056 310796 116068
rect 310751 116028 310796 116056
rect 310790 116016 310796 116028
rect 310848 116016 310854 116068
rect 367002 116056 367008 116068
rect 366963 116028 367008 116056
rect 367002 116016 367008 116028
rect 367060 116016 367066 116068
rect 251450 115988 251456 116000
rect 251411 115960 251456 115988
rect 251450 115948 251456 115960
rect 251508 115948 251514 116000
rect 372706 115988 372712 116000
rect 372667 115960 372712 115988
rect 372706 115948 372712 115960
rect 372764 115948 372770 116000
rect 310790 115920 310796 115932
rect 310751 115892 310796 115920
rect 310790 115880 310796 115892
rect 310848 115880 310854 115932
rect 367002 115920 367008 115932
rect 366963 115892 367008 115920
rect 367002 115880 367008 115892
rect 367060 115880 367066 115932
rect 377033 115923 377091 115929
rect 377033 115889 377045 115923
rect 377079 115920 377091 115923
rect 377122 115920 377128 115932
rect 377079 115892 377128 115920
rect 377079 115889 377091 115892
rect 377033 115883 377091 115889
rect 377122 115880 377128 115892
rect 377180 115880 377186 115932
rect 358722 114560 358728 114572
rect 358683 114532 358728 114560
rect 358722 114520 358728 114532
rect 358780 114520 358786 114572
rect 267826 114492 267832 114504
rect 267787 114464 267832 114492
rect 267826 114452 267832 114464
rect 267884 114452 267890 114504
rect 374362 114492 374368 114504
rect 374323 114464 374368 114492
rect 374362 114452 374368 114464
rect 374420 114452 374426 114504
rect 375834 114492 375840 114504
rect 375795 114464 375840 114492
rect 375834 114452 375840 114464
rect 375892 114452 375898 114504
rect 301130 114424 301136 114436
rect 301091 114396 301136 114424
rect 301130 114384 301136 114396
rect 301188 114384 301194 114436
rect 235074 113200 235080 113212
rect 235035 113172 235080 113200
rect 235074 113160 235080 113172
rect 235132 113160 235138 113212
rect 289998 113200 290004 113212
rect 289959 113172 290004 113200
rect 289998 113160 290004 113172
rect 290056 113160 290062 113212
rect 296898 113200 296904 113212
rect 296859 113172 296904 113200
rect 296898 113160 296904 113172
rect 296956 113160 296962 113212
rect 302418 113160 302424 113212
rect 302476 113200 302482 113212
rect 302602 113200 302608 113212
rect 302476 113172 302608 113200
rect 302476 113160 302482 113172
rect 302602 113160 302608 113172
rect 302660 113160 302666 113212
rect 306650 113200 306656 113212
rect 306611 113172 306656 113200
rect 306650 113160 306656 113172
rect 306708 113160 306714 113212
rect 330110 113200 330116 113212
rect 330071 113172 330116 113200
rect 330110 113160 330116 113172
rect 330168 113160 330174 113212
rect 327169 113135 327227 113141
rect 327169 113101 327181 113135
rect 327215 113132 327227 113135
rect 327258 113132 327264 113144
rect 327215 113104 327264 113132
rect 327215 113101 327227 113104
rect 327169 113095 327227 113101
rect 327258 113092 327264 113104
rect 327316 113092 327322 113144
rect 295518 111800 295524 111852
rect 295576 111840 295582 111852
rect 295797 111843 295855 111849
rect 295797 111840 295809 111843
rect 295576 111812 295809 111840
rect 295576 111800 295582 111812
rect 295797 111809 295809 111812
rect 295843 111809 295855 111843
rect 295797 111803 295855 111809
rect 456518 110644 456524 110696
rect 456576 110684 456582 110696
rect 458818 110684 458824 110696
rect 456576 110656 458824 110684
rect 456576 110644 456582 110656
rect 458818 110644 458824 110656
rect 458876 110644 458882 110696
rect 307662 110576 307668 110628
rect 307720 110616 307726 110628
rect 315942 110616 315948 110628
rect 307720 110588 315948 110616
rect 307720 110576 307726 110588
rect 315942 110576 315948 110588
rect 316000 110576 316006 110628
rect 417878 110576 417884 110628
rect 417936 110616 417942 110628
rect 418154 110616 418160 110628
rect 417936 110588 418160 110616
rect 417936 110576 417942 110588
rect 418154 110576 418160 110588
rect 418212 110576 418218 110628
rect 437198 110576 437204 110628
rect 437256 110616 437262 110628
rect 437474 110616 437480 110628
rect 437256 110588 437480 110616
rect 437256 110576 437262 110588
rect 437474 110576 437480 110588
rect 437532 110576 437538 110628
rect 270402 110440 270408 110492
rect 270460 110480 270466 110492
rect 278682 110480 278688 110492
rect 270460 110452 278688 110480
rect 270460 110440 270466 110452
rect 278682 110440 278688 110452
rect 278740 110440 278746 110492
rect 272150 109012 272156 109064
rect 272208 109012 272214 109064
rect 463786 109012 463792 109064
rect 463844 109052 463850 109064
rect 463970 109052 463976 109064
rect 463844 109024 463976 109052
rect 463844 109012 463850 109024
rect 463970 109012 463976 109024
rect 464028 109012 464034 109064
rect 272168 108928 272196 109012
rect 278774 108944 278780 108996
rect 278832 108984 278838 108996
rect 279050 108984 279056 108996
rect 278832 108956 279056 108984
rect 278832 108944 278838 108956
rect 279050 108944 279056 108956
rect 279108 108944 279114 108996
rect 310790 108984 310796 108996
rect 310751 108956 310796 108984
rect 310790 108944 310796 108956
rect 310848 108944 310854 108996
rect 272150 108876 272156 108928
rect 272208 108876 272214 108928
rect 265158 106292 265164 106344
rect 265216 106332 265222 106344
rect 265250 106332 265256 106344
rect 265216 106304 265256 106332
rect 265216 106292 265222 106304
rect 265250 106292 265256 106304
rect 265308 106292 265314 106344
rect 367002 106332 367008 106344
rect 366963 106304 367008 106332
rect 367002 106292 367008 106304
rect 367060 106292 367066 106344
rect 377030 106332 377036 106344
rect 376991 106304 377036 106332
rect 377030 106292 377036 106304
rect 377088 106292 377094 106344
rect 251450 106264 251456 106276
rect 251411 106236 251456 106264
rect 251450 106224 251456 106236
rect 251508 106224 251514 106276
rect 259546 106224 259552 106276
rect 259604 106264 259610 106276
rect 259822 106264 259828 106276
rect 259604 106236 259828 106264
rect 259604 106224 259610 106236
rect 259822 106224 259828 106236
rect 259880 106224 259886 106276
rect 266633 106267 266691 106273
rect 266633 106233 266645 106267
rect 266679 106264 266691 106267
rect 266722 106264 266728 106276
rect 266679 106236 266728 106264
rect 266679 106233 266691 106236
rect 266633 106227 266691 106233
rect 266722 106224 266728 106236
rect 266780 106224 266786 106276
rect 270678 106224 270684 106276
rect 270736 106224 270742 106276
rect 272150 106224 272156 106276
rect 272208 106264 272214 106276
rect 272242 106264 272248 106276
rect 272208 106236 272248 106264
rect 272208 106224 272214 106236
rect 272242 106224 272248 106236
rect 272300 106224 272306 106276
rect 317690 106224 317696 106276
rect 317748 106264 317754 106276
rect 317874 106264 317880 106276
rect 317748 106236 317880 106264
rect 317748 106224 317754 106236
rect 317874 106224 317880 106236
rect 317932 106224 317938 106276
rect 357526 106224 357532 106276
rect 357584 106264 357590 106276
rect 357618 106264 357624 106276
rect 357584 106236 357624 106264
rect 357584 106224 357590 106236
rect 357618 106224 357624 106236
rect 357676 106224 357682 106276
rect 377122 106264 377128 106276
rect 377083 106236 377128 106264
rect 377122 106224 377128 106236
rect 377180 106224 377186 106276
rect 267826 106196 267832 106208
rect 267787 106168 267832 106196
rect 267826 106156 267832 106168
rect 267884 106156 267890 106208
rect 270696 106140 270724 106224
rect 270678 106088 270684 106140
rect 270736 106088 270742 106140
rect 374362 104972 374368 104984
rect 374323 104944 374368 104972
rect 374362 104932 374368 104944
rect 374420 104932 374426 104984
rect 375834 104972 375840 104984
rect 375795 104944 375840 104972
rect 375834 104932 375840 104944
rect 375892 104932 375898 104984
rect 288710 104864 288716 104916
rect 288768 104904 288774 104916
rect 288894 104904 288900 104916
rect 288768 104876 288900 104904
rect 288768 104864 288774 104876
rect 288894 104864 288900 104876
rect 288952 104864 288958 104916
rect 291562 104864 291568 104916
rect 291620 104904 291626 104916
rect 291654 104904 291660 104916
rect 291620 104876 291660 104904
rect 291620 104864 291626 104876
rect 291654 104864 291660 104876
rect 291712 104864 291718 104916
rect 296806 104864 296812 104916
rect 296864 104904 296870 104916
rect 296898 104904 296904 104916
rect 296864 104876 296904 104904
rect 296864 104864 296870 104876
rect 296898 104864 296904 104876
rect 296956 104864 296962 104916
rect 302418 104864 302424 104916
rect 302476 104904 302482 104916
rect 302510 104904 302516 104916
rect 302476 104876 302516 104904
rect 302476 104864 302482 104876
rect 302510 104864 302516 104876
rect 302568 104864 302574 104916
rect 306650 104864 306656 104916
rect 306708 104904 306714 104916
rect 306834 104904 306840 104916
rect 306708 104876 306840 104904
rect 306708 104864 306714 104876
rect 306834 104864 306840 104876
rect 306892 104864 306898 104916
rect 325878 104904 325884 104916
rect 325839 104876 325884 104904
rect 325878 104864 325884 104876
rect 325936 104864 325942 104916
rect 230842 104836 230848 104848
rect 230803 104808 230848 104836
rect 230842 104796 230848 104808
rect 230900 104796 230906 104848
rect 265158 104836 265164 104848
rect 265119 104808 265164 104836
rect 265158 104796 265164 104808
rect 265216 104796 265222 104848
rect 267826 104836 267832 104848
rect 267787 104808 267832 104836
rect 267826 104796 267832 104808
rect 267884 104796 267890 104848
rect 272242 104836 272248 104848
rect 272203 104808 272248 104836
rect 272242 104796 272248 104808
rect 272300 104796 272306 104848
rect 273530 104836 273536 104848
rect 273491 104808 273536 104836
rect 273530 104796 273536 104808
rect 273588 104796 273594 104848
rect 301130 104796 301136 104848
rect 301188 104836 301194 104848
rect 301314 104836 301320 104848
rect 301188 104808 301320 104836
rect 301188 104796 301194 104808
rect 301314 104796 301320 104808
rect 301372 104796 301378 104848
rect 357618 104836 357624 104848
rect 357579 104808 357624 104836
rect 357618 104796 357624 104808
rect 357676 104796 357682 104848
rect 358722 104836 358728 104848
rect 358683 104808 358728 104836
rect 358722 104796 358728 104808
rect 358780 104796 358786 104848
rect 374362 104836 374368 104848
rect 374323 104808 374368 104836
rect 374362 104796 374368 104808
rect 374420 104796 374426 104848
rect 375834 104836 375840 104848
rect 375795 104808 375840 104836
rect 375834 104796 375840 104808
rect 375892 104796 375898 104848
rect 327166 103544 327172 103556
rect 327127 103516 327172 103544
rect 327166 103504 327172 103516
rect 327224 103504 327230 103556
rect 285950 103476 285956 103488
rect 285911 103448 285956 103476
rect 285950 103436 285956 103448
rect 286008 103436 286014 103488
rect 288710 103436 288716 103488
rect 288768 103436 288774 103488
rect 337102 103436 337108 103488
rect 337160 103476 337166 103488
rect 337197 103479 337255 103485
rect 337197 103476 337209 103479
rect 337160 103448 337209 103476
rect 337160 103436 337166 103448
rect 337197 103445 337209 103448
rect 337243 103445 337255 103479
rect 337197 103439 337255 103445
rect 341061 103479 341119 103485
rect 341061 103445 341073 103479
rect 341107 103476 341119 103479
rect 341150 103476 341156 103488
rect 341107 103448 341156 103476
rect 341107 103445 341119 103448
rect 341061 103439 341119 103445
rect 341150 103436 341156 103448
rect 341208 103436 341214 103488
rect 288728 103408 288756 103436
rect 288802 103408 288808 103420
rect 288728 103380 288808 103408
rect 288802 103368 288808 103380
rect 288860 103368 288866 103420
rect 295518 101980 295524 101992
rect 295479 101952 295524 101980
rect 295518 101940 295524 101952
rect 295576 101940 295582 101992
rect 235074 101396 235080 101448
rect 235132 101436 235138 101448
rect 235258 101436 235264 101448
rect 235132 101408 235264 101436
rect 235132 101396 235138 101408
rect 235258 101396 235264 101408
rect 235316 101396 235322 101448
rect 232222 100036 232228 100088
rect 232280 100076 232286 100088
rect 232317 100079 232375 100085
rect 232317 100076 232329 100079
rect 232280 100048 232329 100076
rect 232280 100036 232286 100048
rect 232317 100045 232329 100048
rect 232363 100045 232375 100079
rect 232317 100039 232375 100045
rect 270678 100036 270684 100088
rect 270736 100076 270742 100088
rect 270862 100076 270868 100088
rect 270736 100048 270868 100076
rect 270736 100036 270742 100048
rect 270862 100036 270868 100048
rect 270920 100036 270926 100088
rect 294230 100036 294236 100088
rect 294288 100076 294294 100088
rect 294414 100076 294420 100088
rect 294288 100048 294420 100076
rect 294288 100036 294294 100048
rect 294414 100036 294420 100048
rect 294472 100036 294478 100088
rect 323394 99424 323400 99476
rect 323452 99424 323458 99476
rect 239122 99356 239128 99408
rect 239180 99356 239186 99408
rect 244366 99356 244372 99408
rect 244424 99396 244430 99408
rect 244424 99368 244504 99396
rect 244424 99356 244430 99368
rect 239140 99272 239168 99356
rect 244476 99340 244504 99368
rect 278866 99356 278872 99408
rect 278924 99396 278930 99408
rect 279050 99396 279056 99408
rect 278924 99368 279056 99396
rect 278924 99356 278930 99368
rect 279050 99356 279056 99368
rect 279108 99356 279114 99408
rect 323412 99340 323440 99424
rect 244458 99288 244464 99340
rect 244516 99288 244522 99340
rect 323394 99288 323400 99340
rect 323452 99288 323458 99340
rect 374362 99328 374368 99340
rect 374323 99300 374368 99328
rect 374362 99288 374368 99300
rect 374420 99288 374426 99340
rect 377122 99328 377128 99340
rect 377083 99300 377128 99328
rect 377122 99288 377128 99300
rect 377180 99288 377186 99340
rect 239122 99220 239128 99272
rect 239180 99220 239186 99272
rect 389361 99195 389419 99201
rect 389361 99161 389373 99195
rect 389407 99192 389419 99195
rect 389450 99192 389456 99204
rect 389407 99164 389456 99192
rect 389407 99161 389419 99164
rect 389361 99155 389419 99161
rect 389450 99152 389456 99164
rect 389508 99152 389514 99204
rect 306834 98676 306840 98728
rect 306892 98716 306898 98728
rect 307018 98716 307024 98728
rect 306892 98688 307024 98716
rect 306892 98676 306898 98688
rect 307018 98676 307024 98688
rect 307076 98676 307082 98728
rect 330202 98716 330208 98728
rect 330163 98688 330208 98716
rect 330202 98676 330208 98688
rect 330260 98676 330266 98728
rect 310882 96812 310888 96824
rect 310808 96784 310888 96812
rect 310808 96688 310836 96784
rect 310882 96772 310888 96784
rect 310940 96772 310946 96824
rect 250070 96636 250076 96688
rect 250128 96676 250134 96688
rect 250162 96676 250168 96688
rect 250128 96648 250168 96676
rect 250128 96636 250134 96648
rect 250162 96636 250168 96648
rect 250220 96636 250226 96688
rect 251450 96676 251456 96688
rect 251411 96648 251456 96676
rect 251450 96636 251456 96648
rect 251508 96636 251514 96688
rect 266630 96676 266636 96688
rect 266591 96648 266636 96676
rect 266630 96636 266636 96648
rect 266688 96636 266694 96688
rect 302510 96636 302516 96688
rect 302568 96636 302574 96688
rect 310790 96636 310796 96688
rect 310848 96636 310854 96688
rect 236270 96608 236276 96620
rect 236231 96580 236276 96608
rect 236270 96568 236276 96580
rect 236328 96568 236334 96620
rect 247126 96608 247132 96620
rect 247087 96580 247132 96608
rect 247126 96568 247132 96580
rect 247184 96568 247190 96620
rect 265158 96608 265164 96620
rect 265119 96580 265164 96608
rect 265158 96568 265164 96580
rect 265216 96568 265222 96620
rect 272245 96543 272303 96549
rect 272245 96509 272257 96543
rect 272291 96540 272303 96543
rect 272334 96540 272340 96552
rect 272291 96512 272340 96540
rect 272291 96509 272303 96512
rect 272245 96503 272303 96509
rect 272334 96500 272340 96512
rect 272392 96500 272398 96552
rect 302528 96540 302556 96636
rect 317782 96608 317788 96620
rect 317743 96580 317788 96608
rect 317782 96568 317788 96580
rect 317840 96568 317846 96620
rect 360286 96568 360292 96620
rect 360344 96608 360350 96620
rect 360378 96608 360384 96620
rect 360344 96580 360384 96608
rect 360344 96568 360350 96580
rect 360378 96568 360384 96580
rect 360436 96568 360442 96620
rect 367002 96608 367008 96620
rect 366963 96580 367008 96608
rect 367002 96568 367008 96580
rect 367060 96568 367066 96620
rect 302602 96540 302608 96552
rect 302528 96512 302608 96540
rect 302602 96500 302608 96512
rect 302660 96500 302666 96552
rect 325970 95276 325976 95328
rect 326028 95316 326034 95328
rect 326028 95288 326108 95316
rect 326028 95276 326034 95288
rect 326080 95260 326108 95288
rect 230842 95248 230848 95260
rect 230803 95220 230848 95248
rect 230842 95208 230848 95220
rect 230900 95208 230906 95260
rect 267829 95251 267887 95257
rect 267829 95217 267841 95251
rect 267875 95248 267887 95251
rect 267918 95248 267924 95260
rect 267875 95220 267924 95248
rect 267875 95217 267887 95220
rect 267829 95211 267887 95217
rect 267918 95208 267924 95220
rect 267976 95208 267982 95260
rect 273533 95251 273591 95257
rect 273533 95217 273545 95251
rect 273579 95248 273591 95251
rect 273622 95248 273628 95260
rect 273579 95220 273628 95248
rect 273579 95217 273591 95220
rect 273533 95211 273591 95217
rect 273622 95208 273628 95220
rect 273680 95208 273686 95260
rect 296806 95208 296812 95260
rect 296864 95208 296870 95260
rect 326062 95208 326068 95260
rect 326120 95208 326126 95260
rect 357618 95248 357624 95260
rect 357579 95220 357624 95248
rect 357618 95208 357624 95220
rect 357676 95208 357682 95260
rect 358725 95251 358783 95257
rect 358725 95217 358737 95251
rect 358771 95248 358783 95251
rect 358814 95248 358820 95260
rect 358771 95220 358820 95248
rect 358771 95217 358783 95220
rect 358725 95211 358783 95217
rect 358814 95208 358820 95220
rect 358872 95208 358878 95260
rect 375834 95248 375840 95260
rect 375795 95220 375840 95248
rect 375834 95208 375840 95220
rect 375892 95208 375898 95260
rect 289998 95140 290004 95192
rect 290056 95180 290062 95192
rect 290090 95180 290096 95192
rect 290056 95152 290096 95180
rect 290056 95140 290062 95152
rect 290090 95140 290096 95152
rect 290148 95140 290154 95192
rect 296824 95112 296852 95208
rect 324590 95140 324596 95192
rect 324648 95180 324654 95192
rect 324774 95180 324780 95192
rect 324648 95152 324780 95180
rect 324648 95140 324654 95152
rect 324774 95140 324780 95152
rect 324832 95140 324838 95192
rect 339678 95140 339684 95192
rect 339736 95180 339742 95192
rect 339773 95183 339831 95189
rect 339773 95180 339785 95183
rect 339736 95152 339785 95180
rect 339736 95140 339742 95152
rect 339773 95149 339785 95152
rect 339819 95149 339831 95183
rect 339773 95143 339831 95149
rect 296990 95112 296996 95124
rect 296824 95084 296996 95112
rect 296990 95072 296996 95084
rect 297048 95072 297054 95124
rect 291654 93916 291660 93968
rect 291712 93916 291718 93968
rect 285953 93891 286011 93897
rect 285953 93857 285965 93891
rect 285999 93888 286011 93891
rect 286134 93888 286140 93900
rect 285999 93860 286140 93888
rect 285999 93857 286011 93860
rect 285953 93851 286011 93857
rect 286134 93848 286140 93860
rect 286192 93848 286198 93900
rect 291672 93888 291700 93916
rect 291746 93888 291752 93900
rect 291672 93860 291752 93888
rect 291746 93848 291752 93860
rect 291804 93848 291810 93900
rect 337194 93848 337200 93900
rect 337252 93888 337258 93900
rect 337252 93860 337297 93888
rect 337252 93848 337258 93860
rect 463694 93848 463700 93900
rect 463752 93888 463758 93900
rect 463878 93888 463884 93900
rect 463752 93860 463884 93888
rect 463752 93848 463758 93860
rect 463878 93848 463884 93860
rect 463936 93848 463942 93900
rect 301130 93820 301136 93832
rect 301091 93792 301136 93820
rect 301130 93780 301136 93792
rect 301188 93780 301194 93832
rect 306742 93820 306748 93832
rect 306703 93792 306748 93820
rect 306742 93780 306748 93792
rect 306800 93780 306806 93832
rect 295521 92531 295579 92537
rect 295521 92497 295533 92531
rect 295567 92528 295579 92531
rect 295702 92528 295708 92540
rect 295567 92500 295708 92528
rect 295567 92497 295579 92500
rect 295521 92491 295579 92497
rect 295702 92488 295708 92500
rect 295760 92488 295766 92540
rect 267918 92420 267924 92472
rect 267976 92460 267982 92472
rect 268102 92460 268108 92472
rect 267976 92432 268108 92460
rect 267976 92420 267982 92432
rect 268102 92420 268108 92432
rect 268160 92420 268166 92472
rect 327258 90380 327264 90432
rect 327316 90420 327322 90432
rect 327442 90420 327448 90432
rect 327316 90392 327448 90420
rect 327316 90380 327322 90392
rect 327442 90380 327448 90392
rect 327500 90380 327506 90432
rect 337010 90380 337016 90432
rect 337068 90420 337074 90432
rect 337194 90420 337200 90432
rect 337068 90392 337200 90420
rect 337068 90380 337074 90392
rect 337194 90380 337200 90392
rect 337252 90380 337258 90432
rect 284754 90216 284760 90228
rect 284715 90188 284760 90216
rect 284754 90176 284760 90188
rect 284812 90176 284818 90228
rect 247126 89672 247132 89684
rect 247087 89644 247132 89672
rect 247126 89632 247132 89644
rect 247184 89632 247190 89684
rect 317782 89672 317788 89684
rect 317743 89644 317788 89672
rect 317782 89632 317788 89644
rect 317840 89632 317846 89684
rect 389358 87904 389364 87916
rect 389319 87876 389364 87904
rect 389358 87864 389364 87876
rect 389416 87864 389422 87916
rect 336918 87184 336924 87236
rect 336976 87184 336982 87236
rect 395890 87184 395896 87236
rect 395948 87184 395954 87236
rect 395982 87184 395988 87236
rect 396040 87184 396046 87236
rect 251174 87048 251180 87100
rect 251232 87088 251238 87100
rect 260650 87088 260656 87100
rect 251232 87060 260656 87088
rect 251232 87048 251238 87060
rect 260650 87048 260656 87060
rect 260708 87048 260714 87100
rect 336936 87032 336964 87184
rect 376754 87048 376760 87100
rect 376812 87088 376818 87100
rect 386230 87088 386236 87100
rect 376812 87060 386236 87088
rect 376812 87048 376818 87060
rect 386230 87048 386236 87060
rect 386288 87048 386294 87100
rect 386414 87048 386420 87100
rect 386472 87088 386478 87100
rect 395798 87088 395804 87100
rect 386472 87060 395804 87088
rect 386472 87048 386478 87060
rect 395798 87048 395804 87060
rect 395856 87048 395862 87100
rect 395908 87032 395936 87184
rect 396000 87032 396028 87184
rect 437198 87116 437204 87168
rect 437256 87156 437262 87168
rect 437474 87156 437480 87168
rect 437256 87128 437480 87156
rect 437256 87116 437262 87128
rect 437474 87116 437480 87128
rect 437532 87116 437538 87168
rect 456518 87116 456524 87168
rect 456576 87156 456582 87168
rect 456978 87156 456984 87168
rect 456576 87128 456984 87156
rect 456576 87116 456582 87128
rect 456978 87116 456984 87128
rect 457036 87116 457042 87168
rect 494606 87116 494612 87168
rect 494664 87156 494670 87168
rect 502242 87156 502248 87168
rect 494664 87128 502248 87156
rect 494664 87116 494670 87128
rect 502242 87116 502248 87128
rect 502300 87116 502306 87168
rect 417878 87048 417884 87100
rect 417936 87088 417942 87100
rect 418154 87088 418160 87100
rect 417936 87060 418160 87088
rect 417936 87048 417942 87060
rect 418154 87048 418160 87060
rect 418212 87048 418218 87100
rect 232314 87020 232320 87032
rect 232275 86992 232320 87020
rect 232314 86980 232320 86992
rect 232372 86980 232378 87032
rect 236270 87020 236276 87032
rect 236231 86992 236276 87020
rect 236270 86980 236276 86992
rect 236328 86980 236334 87032
rect 295702 86980 295708 87032
rect 295760 86980 295766 87032
rect 326062 87020 326068 87032
rect 325988 86992 326068 87020
rect 251450 86952 251456 86964
rect 251411 86924 251456 86952
rect 251450 86912 251456 86924
rect 251508 86912 251514 86964
rect 295720 86896 295748 86980
rect 325988 86964 326016 86992
rect 326062 86980 326068 86992
rect 326120 86980 326126 87032
rect 336918 86980 336924 87032
rect 336976 86980 336982 87032
rect 367002 87020 367008 87032
rect 366963 86992 367008 87020
rect 367002 86980 367008 86992
rect 367060 86980 367066 87032
rect 395890 86980 395896 87032
rect 395948 86980 395954 87032
rect 395982 86980 395988 87032
rect 396040 86980 396046 87032
rect 325970 86912 325976 86964
rect 326028 86912 326034 86964
rect 330202 86952 330208 86964
rect 330163 86924 330208 86952
rect 330202 86912 330208 86924
rect 330260 86912 330266 86964
rect 331306 86912 331312 86964
rect 331364 86912 331370 86964
rect 331398 86912 331404 86964
rect 331456 86912 331462 86964
rect 360197 86955 360255 86961
rect 360197 86921 360209 86955
rect 360243 86952 360255 86955
rect 360378 86952 360384 86964
rect 360243 86924 360384 86952
rect 360243 86921 360255 86924
rect 360197 86915 360255 86921
rect 360378 86912 360384 86924
rect 360436 86912 360442 86964
rect 295702 86844 295708 86896
rect 295760 86844 295766 86896
rect 301133 86887 301191 86893
rect 301133 86853 301145 86887
rect 301179 86884 301191 86887
rect 301222 86884 301228 86896
rect 301179 86856 301228 86884
rect 301179 86853 301191 86856
rect 301133 86847 301191 86853
rect 301222 86844 301228 86856
rect 301280 86844 301286 86896
rect 317690 86844 317696 86896
rect 317748 86884 317754 86896
rect 317874 86884 317880 86896
rect 317748 86856 317880 86884
rect 317748 86844 317754 86856
rect 317874 86844 317880 86856
rect 317932 86844 317938 86896
rect 331324 86828 331352 86912
rect 331416 86828 331444 86912
rect 331306 86776 331312 86828
rect 331364 86776 331370 86828
rect 331398 86776 331404 86828
rect 331456 86776 331462 86828
rect 286134 85660 286140 85672
rect 286060 85632 286140 85660
rect 286060 85604 286088 85632
rect 286134 85620 286140 85632
rect 286192 85620 286198 85672
rect 284754 85592 284760 85604
rect 284715 85564 284760 85592
rect 284754 85552 284760 85564
rect 284812 85552 284818 85604
rect 286042 85552 286048 85604
rect 286100 85552 286106 85604
rect 291565 85595 291623 85601
rect 291565 85561 291577 85595
rect 291611 85592 291623 85595
rect 291654 85592 291660 85604
rect 291611 85564 291660 85592
rect 291611 85561 291623 85564
rect 291565 85555 291623 85561
rect 291654 85552 291660 85564
rect 291712 85552 291718 85604
rect 294230 85552 294236 85604
rect 294288 85592 294294 85604
rect 294414 85592 294420 85604
rect 294288 85564 294420 85592
rect 294288 85552 294294 85564
rect 294414 85552 294420 85564
rect 294472 85552 294478 85604
rect 358538 85552 358544 85604
rect 358596 85592 358602 85604
rect 358630 85592 358636 85604
rect 358596 85564 358636 85592
rect 358596 85552 358602 85564
rect 358630 85552 358636 85564
rect 358688 85552 358694 85604
rect 232314 85524 232320 85536
rect 232275 85496 232320 85524
rect 232314 85484 232320 85496
rect 232372 85484 232378 85536
rect 236270 85524 236276 85536
rect 236231 85496 236276 85524
rect 236270 85484 236276 85496
rect 236328 85484 236334 85536
rect 324593 85527 324651 85533
rect 324593 85493 324605 85527
rect 324639 85524 324651 85527
rect 324682 85524 324688 85536
rect 324639 85496 324688 85524
rect 324639 85493 324651 85496
rect 324593 85487 324651 85493
rect 324682 85484 324688 85496
rect 324740 85484 324746 85536
rect 357526 85524 357532 85536
rect 357487 85496 357532 85524
rect 357526 85484 357532 85496
rect 357584 85484 357590 85536
rect 291562 84232 291568 84244
rect 291523 84204 291568 84232
rect 291562 84192 291568 84204
rect 291620 84192 291626 84244
rect 306745 84235 306803 84241
rect 306745 84201 306757 84235
rect 306791 84232 306803 84235
rect 306834 84232 306840 84244
rect 306791 84204 306840 84232
rect 306791 84201 306803 84204
rect 306745 84195 306803 84201
rect 306834 84192 306840 84204
rect 306892 84192 306898 84244
rect 270770 84164 270776 84176
rect 270731 84136 270776 84164
rect 270770 84124 270776 84136
rect 270828 84124 270834 84176
rect 284754 84164 284760 84176
rect 284715 84136 284760 84164
rect 284754 84124 284760 84136
rect 284812 84124 284818 84176
rect 337010 84124 337016 84176
rect 337068 84124 337074 84176
rect 337028 84096 337056 84124
rect 337197 84099 337255 84105
rect 337197 84096 337209 84099
rect 337028 84068 337209 84096
rect 337197 84065 337209 84068
rect 337243 84065 337255 84099
rect 337197 84059 337255 84065
rect 265250 82804 265256 82816
rect 265211 82776 265256 82804
rect 265250 82764 265256 82776
rect 265308 82764 265314 82816
rect 267826 82764 267832 82816
rect 267884 82804 267890 82816
rect 268010 82804 268016 82816
rect 267884 82776 268016 82804
rect 267884 82764 267890 82776
rect 268010 82764 268016 82776
rect 268068 82764 268074 82816
rect 301222 82804 301228 82816
rect 301183 82776 301228 82804
rect 301222 82764 301228 82776
rect 301280 82764 301286 82816
rect 302602 82804 302608 82816
rect 302563 82776 302608 82804
rect 302602 82764 302608 82776
rect 302660 82764 302666 82816
rect 249794 80724 249800 80776
rect 249852 80764 249858 80776
rect 250070 80764 250076 80776
rect 249852 80736 250076 80764
rect 249852 80724 249858 80736
rect 250070 80724 250076 80736
rect 250128 80724 250134 80776
rect 247218 80220 247224 80232
rect 247179 80192 247224 80220
rect 247218 80180 247224 80192
rect 247276 80180 247282 80232
rect 234982 80044 234988 80096
rect 235040 80084 235046 80096
rect 235166 80084 235172 80096
rect 235040 80056 235172 80084
rect 235040 80044 235046 80056
rect 235166 80044 235172 80056
rect 235224 80044 235230 80096
rect 303890 80044 303896 80096
rect 303948 80044 303954 80096
rect 338850 80044 338856 80096
rect 338908 80044 338914 80096
rect 389358 80044 389364 80096
rect 389416 80044 389422 80096
rect 463786 80044 463792 80096
rect 463844 80044 463850 80096
rect 303908 79960 303936 80044
rect 338868 79960 338896 80044
rect 303890 79908 303896 79960
rect 303948 79908 303954 79960
rect 338850 79908 338856 79960
rect 338908 79908 338914 79960
rect 372430 79908 372436 79960
rect 372488 79948 372494 79960
rect 372798 79948 372804 79960
rect 372488 79920 372804 79948
rect 372488 79908 372494 79920
rect 372798 79908 372804 79920
rect 372856 79908 372862 79960
rect 389376 79948 389404 80044
rect 463804 79960 463832 80044
rect 389450 79948 389456 79960
rect 389376 79920 389456 79948
rect 389450 79908 389456 79920
rect 389508 79908 389514 79960
rect 463786 79908 463792 79960
rect 463844 79908 463850 79960
rect 2774 79840 2780 79892
rect 2832 79880 2838 79892
rect 4982 79880 4988 79892
rect 2832 79852 4988 79880
rect 2832 79840 2838 79852
rect 4982 79840 4988 79852
rect 5040 79840 5046 79892
rect 285953 78523 286011 78529
rect 285953 78489 285965 78523
rect 285999 78520 286011 78523
rect 286042 78520 286048 78532
rect 285999 78492 286048 78520
rect 285999 78489 286011 78492
rect 285953 78483 286011 78489
rect 286042 78480 286048 78492
rect 286100 78480 286106 78532
rect 367002 77392 367008 77444
rect 367060 77392 367066 77444
rect 336826 77324 336832 77376
rect 336884 77324 336890 77376
rect 336918 77324 336924 77376
rect 336976 77324 336982 77376
rect 247218 77296 247224 77308
rect 247179 77268 247224 77296
rect 247218 77256 247224 77268
rect 247276 77256 247282 77308
rect 251450 77296 251456 77308
rect 251411 77268 251456 77296
rect 251450 77256 251456 77268
rect 251508 77256 251514 77308
rect 266630 77256 266636 77308
rect 266688 77296 266694 77308
rect 266722 77296 266728 77308
rect 266688 77268 266728 77296
rect 266688 77256 266694 77268
rect 266722 77256 266728 77268
rect 266780 77256 266786 77308
rect 299750 77256 299756 77308
rect 299808 77296 299814 77308
rect 299842 77296 299848 77308
rect 299808 77268 299848 77296
rect 299808 77256 299814 77268
rect 299842 77256 299848 77268
rect 299900 77256 299906 77308
rect 323394 77296 323400 77308
rect 323355 77268 323400 77296
rect 323394 77256 323400 77268
rect 323452 77256 323458 77308
rect 336844 77240 336872 77324
rect 336936 77240 336964 77324
rect 367020 77308 367048 77392
rect 339770 77296 339776 77308
rect 339731 77268 339776 77296
rect 339770 77256 339776 77268
rect 339828 77256 339834 77308
rect 341058 77296 341064 77308
rect 341019 77268 341064 77296
rect 341058 77256 341064 77268
rect 341116 77256 341122 77308
rect 360194 77296 360200 77308
rect 360155 77268 360200 77296
rect 360194 77256 360200 77268
rect 360252 77256 360258 77308
rect 367002 77256 367008 77308
rect 367060 77256 367066 77308
rect 272242 77188 272248 77240
rect 272300 77228 272306 77240
rect 272334 77228 272340 77240
rect 272300 77200 272340 77228
rect 272300 77188 272306 77200
rect 272334 77188 272340 77200
rect 272392 77188 272398 77240
rect 303890 77188 303896 77240
rect 303948 77228 303954 77240
rect 303982 77228 303988 77240
rect 303948 77200 303988 77228
rect 303948 77188 303954 77200
rect 303982 77188 303988 77200
rect 304040 77188 304046 77240
rect 336826 77188 336832 77240
rect 336884 77188 336890 77240
rect 336918 77188 336924 77240
rect 336976 77188 336982 77240
rect 389361 77231 389419 77237
rect 389361 77197 389373 77231
rect 389407 77228 389419 77231
rect 389450 77228 389456 77240
rect 389407 77200 389456 77228
rect 389407 77197 389419 77200
rect 389361 77191 389419 77197
rect 389450 77188 389456 77200
rect 389508 77188 389514 77240
rect 341058 77160 341064 77172
rect 341019 77132 341064 77160
rect 341058 77120 341064 77132
rect 341116 77120 341122 77172
rect 309042 76236 309048 76288
rect 309100 76276 309106 76288
rect 317322 76276 317328 76288
rect 309100 76248 317328 76276
rect 309100 76236 309106 76248
rect 317322 76236 317328 76248
rect 317380 76236 317386 76288
rect 417878 76100 417884 76152
rect 417936 76140 417942 76152
rect 420362 76140 420368 76152
rect 417936 76112 420368 76140
rect 417936 76100 417942 76112
rect 420362 76100 420368 76112
rect 420420 76100 420426 76152
rect 253842 76032 253848 76084
rect 253900 76072 253906 76084
rect 259270 76072 259276 76084
rect 253900 76044 259276 76072
rect 253900 76032 253906 76044
rect 259270 76032 259276 76044
rect 259328 76032 259334 76084
rect 437198 76032 437204 76084
rect 437256 76072 437262 76084
rect 437474 76072 437480 76084
rect 437256 76044 437480 76072
rect 437256 76032 437262 76044
rect 437474 76032 437480 76044
rect 437532 76032 437538 76084
rect 456518 76032 456524 76084
rect 456576 76072 456582 76084
rect 456794 76072 456800 76084
rect 456576 76044 456800 76072
rect 456576 76032 456582 76044
rect 456794 76032 456800 76044
rect 456852 76032 456858 76084
rect 232314 75936 232320 75948
rect 232275 75908 232320 75936
rect 232314 75896 232320 75908
rect 232372 75896 232378 75948
rect 236270 75936 236276 75948
rect 236231 75908 236276 75936
rect 236270 75896 236276 75908
rect 236328 75896 236334 75948
rect 288710 75896 288716 75948
rect 288768 75936 288774 75948
rect 288802 75936 288808 75948
rect 288768 75908 288808 75936
rect 288768 75896 288774 75908
rect 288802 75896 288808 75908
rect 288860 75896 288866 75948
rect 289906 75896 289912 75948
rect 289964 75936 289970 75948
rect 290090 75936 290096 75948
rect 289964 75908 290096 75936
rect 289964 75896 289970 75908
rect 290090 75896 290096 75908
rect 290148 75896 290154 75948
rect 291378 75896 291384 75948
rect 291436 75936 291442 75948
rect 291562 75936 291568 75948
rect 291436 75908 291568 75936
rect 291436 75896 291442 75908
rect 291562 75896 291568 75908
rect 291620 75896 291626 75948
rect 295518 75896 295524 75948
rect 295576 75936 295582 75948
rect 295702 75936 295708 75948
rect 295576 75908 295708 75936
rect 295576 75896 295582 75908
rect 295702 75896 295708 75908
rect 295760 75896 295766 75948
rect 296806 75896 296812 75948
rect 296864 75936 296870 75948
rect 296990 75936 296996 75948
rect 296864 75908 296996 75936
rect 296864 75896 296870 75908
rect 296990 75896 296996 75908
rect 297048 75896 297054 75948
rect 323394 75936 323400 75948
rect 323355 75908 323400 75936
rect 323394 75896 323400 75908
rect 323452 75896 323458 75948
rect 324590 75936 324596 75948
rect 324551 75908 324596 75936
rect 324590 75896 324596 75908
rect 324648 75896 324654 75948
rect 357529 75939 357587 75945
rect 357529 75905 357541 75939
rect 357575 75936 357587 75939
rect 357618 75936 357624 75948
rect 357575 75908 357624 75936
rect 357575 75905 357587 75908
rect 357529 75899 357587 75905
rect 357618 75896 357624 75908
rect 357676 75896 357682 75948
rect 358538 75896 358544 75948
rect 358596 75936 358602 75948
rect 358722 75936 358728 75948
rect 358596 75908 358728 75936
rect 358596 75896 358602 75908
rect 358722 75896 358728 75908
rect 358780 75896 358786 75948
rect 250070 75868 250076 75880
rect 250031 75840 250076 75868
rect 250070 75828 250076 75840
rect 250128 75828 250134 75880
rect 272153 75871 272211 75877
rect 272153 75837 272165 75871
rect 272199 75868 272211 75871
rect 272242 75868 272248 75880
rect 272199 75840 272248 75868
rect 272199 75837 272211 75840
rect 272153 75831 272211 75837
rect 272242 75828 272248 75840
rect 272300 75828 272306 75880
rect 372709 75871 372767 75877
rect 372709 75837 372721 75871
rect 372755 75868 372767 75871
rect 372798 75868 372804 75880
rect 372755 75840 372804 75868
rect 372755 75837 372767 75840
rect 372709 75831 372767 75837
rect 372798 75828 372804 75840
rect 372856 75828 372862 75880
rect 284757 75803 284815 75809
rect 284757 75769 284769 75803
rect 284803 75800 284815 75803
rect 284846 75800 284852 75812
rect 284803 75772 284852 75800
rect 284803 75769 284815 75772
rect 284757 75763 284815 75769
rect 284846 75760 284852 75772
rect 284904 75760 284910 75812
rect 270770 74576 270776 74588
rect 270731 74548 270776 74576
rect 270770 74536 270776 74548
rect 270828 74536 270834 74588
rect 306742 74536 306748 74588
rect 306800 74576 306806 74588
rect 306834 74576 306840 74588
rect 306800 74548 306840 74576
rect 306800 74536 306806 74548
rect 306834 74536 306840 74548
rect 306892 74536 306898 74588
rect 266722 74508 266728 74520
rect 266683 74480 266728 74508
rect 266722 74468 266728 74480
rect 266780 74468 266786 74520
rect 288710 74468 288716 74520
rect 288768 74508 288774 74520
rect 288986 74508 288992 74520
rect 288768 74480 288992 74508
rect 288768 74468 288774 74480
rect 288986 74468 288992 74480
rect 289044 74468 289050 74520
rect 265250 73216 265256 73228
rect 265211 73188 265256 73216
rect 265250 73176 265256 73188
rect 265308 73176 265314 73228
rect 301222 73216 301228 73228
rect 301183 73188 301228 73216
rect 301222 73176 301228 73188
rect 301280 73176 301286 73228
rect 302605 73219 302663 73225
rect 302605 73185 302617 73219
rect 302651 73216 302663 73219
rect 302694 73216 302700 73228
rect 302651 73188 302700 73216
rect 302651 73185 302663 73188
rect 302605 73179 302663 73185
rect 302694 73176 302700 73188
rect 302752 73176 302758 73228
rect 324590 72428 324596 72480
rect 324648 72468 324654 72480
rect 324774 72468 324780 72480
rect 324648 72440 324780 72468
rect 324648 72428 324654 72440
rect 324774 72428 324780 72440
rect 324832 72428 324838 72480
rect 267826 71748 267832 71800
rect 267884 71788 267890 71800
rect 268010 71788 268016 71800
rect 267884 71760 268016 71788
rect 267884 71748 267890 71760
rect 268010 71748 268016 71760
rect 268068 71748 268074 71800
rect 239122 70456 239128 70508
rect 239180 70456 239186 70508
rect 244458 70496 244464 70508
rect 244419 70468 244464 70496
rect 244458 70456 244464 70468
rect 244516 70456 244522 70508
rect 273533 70499 273591 70505
rect 273533 70465 273545 70499
rect 273579 70496 273591 70499
rect 273622 70496 273628 70508
rect 273579 70468 273628 70496
rect 273579 70465 273591 70468
rect 273533 70459 273591 70465
rect 273622 70456 273628 70468
rect 273680 70456 273686 70508
rect 325970 70496 325976 70508
rect 325896 70468 325976 70496
rect 239140 70372 239168 70456
rect 325896 70372 325924 70468
rect 325970 70456 325976 70468
rect 326028 70456 326034 70508
rect 239122 70320 239128 70372
rect 239180 70320 239186 70372
rect 325878 70320 325884 70372
rect 325936 70320 325942 70372
rect 341061 70295 341119 70301
rect 341061 70261 341073 70295
rect 341107 70292 341119 70295
rect 341150 70292 341156 70304
rect 341107 70264 341156 70292
rect 341107 70261 341119 70264
rect 341061 70255 341119 70261
rect 341150 70252 341156 70264
rect 341208 70252 341214 70304
rect 301041 69683 301099 69689
rect 301041 69649 301053 69683
rect 301087 69680 301099 69683
rect 301222 69680 301228 69692
rect 301087 69652 301228 69680
rect 301087 69649 301099 69652
rect 301041 69643 301099 69649
rect 301222 69640 301228 69652
rect 301280 69640 301286 69692
rect 236270 67600 236276 67652
rect 236328 67600 236334 67652
rect 273530 67640 273536 67652
rect 273491 67612 273536 67640
rect 273530 67600 273536 67612
rect 273588 67600 273594 67652
rect 323302 67600 323308 67652
rect 323360 67640 323366 67652
rect 323394 67640 323400 67652
rect 323360 67612 323400 67640
rect 323360 67600 323366 67612
rect 323394 67600 323400 67612
rect 323452 67600 323458 67652
rect 330110 67600 330116 67652
rect 330168 67640 330174 67652
rect 330294 67640 330300 67652
rect 330168 67612 330300 67640
rect 330168 67600 330174 67612
rect 330294 67600 330300 67612
rect 330352 67600 330358 67652
rect 389358 67640 389364 67652
rect 389319 67612 389364 67640
rect 389358 67600 389364 67612
rect 389416 67600 389422 67652
rect 236288 67572 236316 67600
rect 236362 67572 236368 67584
rect 236288 67544 236368 67572
rect 236362 67532 236368 67544
rect 236420 67532 236426 67584
rect 247126 67532 247132 67584
rect 247184 67572 247190 67584
rect 247218 67572 247224 67584
rect 247184 67544 247224 67572
rect 247184 67532 247190 67544
rect 247218 67532 247224 67544
rect 247276 67532 247282 67584
rect 244458 66280 244464 66292
rect 244419 66252 244464 66280
rect 244458 66240 244464 66252
rect 244516 66240 244522 66292
rect 250070 66280 250076 66292
rect 250031 66252 250076 66280
rect 250070 66240 250076 66252
rect 250128 66240 250134 66292
rect 259638 66240 259644 66292
rect 259696 66280 259702 66292
rect 259730 66280 259736 66292
rect 259696 66252 259736 66280
rect 259696 66240 259702 66252
rect 259730 66240 259736 66252
rect 259788 66240 259794 66292
rect 272150 66280 272156 66292
rect 272111 66252 272156 66280
rect 272150 66240 272156 66252
rect 272208 66240 272214 66292
rect 285950 66280 285956 66292
rect 285911 66252 285956 66280
rect 285950 66240 285956 66252
rect 286008 66240 286014 66292
rect 337194 66280 337200 66292
rect 337155 66252 337200 66280
rect 337194 66240 337200 66252
rect 337252 66240 337258 66292
rect 372706 66280 372712 66292
rect 372667 66252 372712 66280
rect 372706 66240 372712 66252
rect 372764 66240 372770 66292
rect 232314 66212 232320 66224
rect 232275 66184 232320 66212
rect 232314 66172 232320 66184
rect 232372 66172 232378 66224
rect 270678 66212 270684 66224
rect 270639 66184 270684 66212
rect 270678 66172 270684 66184
rect 270736 66172 270742 66224
rect 296806 66212 296812 66224
rect 296767 66184 296812 66212
rect 296806 66172 296812 66184
rect 296864 66172 296870 66224
rect 310790 66212 310796 66224
rect 310751 66184 310796 66212
rect 310790 66172 310796 66184
rect 310848 66172 310854 66224
rect 323302 66212 323308 66224
rect 323263 66184 323308 66212
rect 323302 66172 323308 66184
rect 323360 66172 323366 66224
rect 324685 66215 324743 66221
rect 324685 66181 324697 66215
rect 324731 66212 324743 66215
rect 324774 66212 324780 66224
rect 324731 66184 324780 66212
rect 324731 66181 324743 66184
rect 324685 66175 324743 66181
rect 324774 66172 324780 66184
rect 324832 66172 324838 66224
rect 329929 66215 329987 66221
rect 329929 66181 329941 66215
rect 329975 66212 329987 66215
rect 330110 66212 330116 66224
rect 329975 66184 330116 66212
rect 329975 66181 329987 66184
rect 329929 66175 329987 66181
rect 330110 66172 330116 66184
rect 330168 66172 330174 66224
rect 266725 64923 266783 64929
rect 266725 64889 266737 64923
rect 266771 64920 266783 64923
rect 266906 64920 266912 64932
rect 266771 64892 266912 64920
rect 266771 64889 266783 64892
rect 266725 64883 266783 64889
rect 266906 64880 266912 64892
rect 266964 64880 266970 64932
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 24118 64852 24124 64864
rect 3384 64824 24124 64852
rect 3384 64812 3390 64824
rect 24118 64812 24124 64824
rect 24176 64812 24182 64864
rect 294230 64852 294236 64864
rect 294191 64824 294236 64852
rect 294230 64812 294236 64824
rect 294288 64812 294294 64864
rect 273162 63656 273168 63708
rect 273220 63696 273226 63708
rect 278682 63696 278688 63708
rect 273220 63668 278688 63696
rect 273220 63656 273226 63668
rect 278682 63656 278688 63668
rect 278740 63656 278746 63708
rect 417878 63656 417884 63708
rect 417936 63696 417942 63708
rect 418154 63696 418160 63708
rect 417936 63668 418160 63696
rect 417936 63656 417942 63668
rect 418154 63656 418160 63668
rect 418212 63656 418218 63708
rect 437198 63656 437204 63708
rect 437256 63696 437262 63708
rect 437474 63696 437480 63708
rect 437256 63668 437480 63696
rect 437256 63656 437262 63668
rect 437474 63656 437480 63668
rect 437532 63656 437538 63708
rect 456518 63656 456524 63708
rect 456576 63696 456582 63708
rect 456886 63696 456892 63708
rect 456576 63668 456892 63696
rect 456576 63656 456582 63668
rect 456886 63656 456892 63668
rect 456944 63656 456950 63708
rect 265253 63495 265311 63501
rect 265253 63461 265265 63495
rect 265299 63492 265311 63495
rect 265342 63492 265348 63504
rect 265299 63464 265348 63492
rect 265299 63461 265311 63464
rect 265253 63455 265311 63461
rect 265342 63452 265348 63464
rect 265400 63452 265406 63504
rect 230753 61455 230811 61461
rect 230753 61421 230765 61455
rect 230799 61452 230811 61455
rect 230842 61452 230848 61464
rect 230799 61424 230848 61452
rect 230799 61421 230811 61424
rect 230753 61415 230811 61421
rect 230842 61412 230848 61424
rect 230900 61412 230906 61464
rect 236273 61455 236331 61461
rect 236273 61421 236285 61455
rect 236319 61452 236331 61455
rect 236362 61452 236368 61464
rect 236319 61424 236368 61452
rect 236319 61421 236331 61424
rect 236273 61415 236331 61421
rect 236362 61412 236368 61424
rect 236420 61412 236426 61464
rect 272150 60732 272156 60784
rect 272208 60732 272214 60784
rect 272168 60648 272196 60732
rect 273438 60664 273444 60716
rect 273496 60704 273502 60716
rect 273622 60704 273628 60716
rect 273496 60676 273628 60704
rect 273496 60664 273502 60676
rect 273622 60664 273628 60676
rect 273680 60664 273686 60716
rect 310790 60704 310796 60716
rect 310751 60676 310796 60704
rect 310790 60664 310796 60676
rect 310848 60664 310854 60716
rect 341150 60664 341156 60716
rect 341208 60704 341214 60716
rect 341334 60704 341340 60716
rect 341208 60676 341340 60704
rect 341208 60664 341214 60676
rect 341334 60664 341340 60676
rect 341392 60664 341398 60716
rect 360286 60664 360292 60716
rect 360344 60704 360350 60716
rect 360470 60704 360476 60716
rect 360344 60676 360476 60704
rect 360344 60664 360350 60676
rect 360470 60664 360476 60676
rect 360528 60664 360534 60716
rect 272150 60596 272156 60648
rect 272208 60596 272214 60648
rect 262674 60364 262680 60376
rect 262635 60336 262680 60364
rect 262674 60324 262680 60336
rect 262732 60324 262738 60376
rect 302513 59551 302571 59557
rect 302513 59517 302525 59551
rect 302559 59548 302571 59551
rect 302694 59548 302700 59560
rect 302559 59520 302700 59548
rect 302559 59517 302571 59520
rect 302513 59511 302571 59517
rect 302694 59508 302700 59520
rect 302752 59508 302758 59560
rect 325878 58012 325884 58064
rect 325936 58012 325942 58064
rect 284754 57944 284760 57996
rect 284812 57984 284818 57996
rect 284846 57984 284852 57996
rect 284812 57956 284852 57984
rect 284812 57944 284818 57956
rect 284846 57944 284852 57956
rect 284904 57944 284910 57996
rect 285950 57944 285956 57996
rect 286008 57984 286014 57996
rect 286042 57984 286048 57996
rect 286008 57956 286048 57984
rect 286008 57944 286014 57956
rect 286042 57944 286048 57956
rect 286100 57944 286106 57996
rect 325896 57928 325924 58012
rect 327166 57944 327172 57996
rect 327224 57944 327230 57996
rect 325878 57876 325884 57928
rect 325936 57876 325942 57928
rect 327184 57848 327212 57944
rect 341334 57916 341340 57928
rect 341295 57888 341340 57916
rect 341334 57876 341340 57888
rect 341392 57876 341398 57928
rect 360378 57876 360384 57928
rect 360436 57916 360442 57928
rect 360470 57916 360476 57928
rect 360436 57888 360476 57916
rect 360436 57876 360442 57888
rect 360470 57876 360476 57888
rect 360528 57876 360534 57928
rect 367002 57916 367008 57928
rect 366963 57888 367008 57916
rect 367002 57876 367008 57888
rect 367060 57876 367066 57928
rect 389174 57916 389180 57928
rect 389135 57888 389180 57916
rect 389174 57876 389180 57888
rect 389232 57876 389238 57928
rect 470594 57916 470600 57928
rect 470555 57888 470600 57916
rect 470594 57876 470600 57888
rect 470652 57876 470658 57928
rect 327258 57848 327264 57860
rect 327184 57820 327264 57848
rect 327258 57808 327264 57820
rect 327316 57808 327322 57860
rect 295518 57032 295524 57044
rect 295479 57004 295524 57032
rect 295518 56992 295524 57004
rect 295576 56992 295582 57044
rect 232314 56624 232320 56636
rect 232275 56596 232320 56624
rect 232314 56584 232320 56596
rect 232372 56584 232378 56636
rect 259638 56624 259644 56636
rect 259564 56596 259644 56624
rect 259564 56568 259592 56596
rect 259638 56584 259644 56596
rect 259696 56584 259702 56636
rect 324682 56624 324688 56636
rect 324643 56596 324688 56624
rect 324682 56584 324688 56596
rect 324740 56584 324746 56636
rect 329926 56624 329932 56636
rect 329887 56596 329932 56624
rect 329926 56584 329932 56596
rect 329984 56584 329990 56636
rect 358722 56584 358728 56636
rect 358780 56624 358786 56636
rect 358814 56624 358820 56636
rect 358780 56596 358820 56624
rect 358780 56584 358786 56596
rect 358814 56584 358820 56596
rect 358872 56584 358878 56636
rect 250070 56556 250076 56568
rect 250031 56528 250076 56556
rect 250070 56516 250076 56528
rect 250128 56516 250134 56568
rect 259546 56516 259552 56568
rect 259604 56516 259610 56568
rect 285953 56559 286011 56565
rect 285953 56525 285965 56559
rect 285999 56556 286011 56559
rect 286042 56556 286048 56568
rect 285999 56528 286048 56556
rect 285999 56525 286011 56528
rect 285953 56519 286011 56525
rect 286042 56516 286048 56528
rect 286100 56516 286106 56568
rect 310790 56516 310796 56568
rect 310848 56556 310854 56568
rect 310882 56556 310888 56568
rect 310848 56528 310888 56556
rect 310848 56516 310854 56528
rect 310882 56516 310888 56528
rect 310940 56516 310946 56568
rect 339678 56556 339684 56568
rect 339639 56528 339684 56556
rect 339678 56516 339684 56528
rect 339736 56516 339742 56568
rect 296806 56216 296812 56228
rect 296767 56188 296812 56216
rect 296806 56176 296812 56188
rect 296864 56176 296870 56228
rect 262677 55267 262735 55273
rect 262677 55233 262689 55267
rect 262723 55264 262735 55267
rect 262766 55264 262772 55276
rect 262723 55236 262772 55264
rect 262723 55233 262735 55236
rect 262677 55227 262735 55233
rect 262766 55224 262772 55236
rect 262824 55224 262830 55276
rect 294230 55264 294236 55276
rect 294191 55236 294236 55264
rect 294230 55224 294236 55236
rect 294288 55224 294294 55276
rect 317506 55224 317512 55276
rect 317564 55264 317570 55276
rect 317690 55264 317696 55276
rect 317564 55236 317696 55264
rect 317564 55224 317570 55236
rect 317690 55224 317696 55236
rect 317748 55224 317754 55276
rect 300949 55199 301007 55205
rect 300949 55165 300961 55199
rect 300995 55165 301007 55199
rect 300949 55159 301007 55165
rect 300964 55128 300992 55159
rect 301222 55128 301228 55140
rect 300964 55100 301228 55128
rect 301222 55088 301228 55100
rect 301280 55088 301286 55140
rect 244366 53796 244372 53848
rect 244424 53836 244430 53848
rect 244458 53836 244464 53848
rect 244424 53808 244464 53836
rect 244424 53796 244430 53808
rect 244458 53796 244464 53808
rect 244516 53796 244522 53848
rect 265250 53836 265256 53848
rect 265211 53808 265256 53836
rect 265250 53796 265256 53808
rect 265308 53796 265314 53848
rect 232225 53091 232283 53097
rect 232225 53057 232237 53091
rect 232271 53088 232283 53091
rect 232314 53088 232320 53100
rect 232271 53060 232320 53088
rect 232271 53057 232283 53060
rect 232225 53051 232283 53057
rect 232314 53048 232320 53060
rect 232372 53048 232378 53100
rect 267826 52436 267832 52488
rect 267884 52476 267890 52488
rect 268010 52476 268016 52488
rect 267884 52448 268016 52476
rect 267884 52436 267890 52448
rect 268010 52436 268016 52448
rect 268068 52436 268074 52488
rect 270681 52411 270739 52417
rect 270681 52377 270693 52411
rect 270727 52408 270739 52411
rect 270865 52411 270923 52417
rect 270865 52408 270877 52411
rect 270727 52380 270877 52408
rect 270727 52377 270739 52380
rect 270681 52371 270739 52377
rect 270865 52377 270877 52380
rect 270911 52377 270923 52411
rect 270865 52371 270923 52377
rect 273622 51116 273628 51128
rect 273548 51088 273628 51116
rect 273548 51060 273576 51088
rect 273622 51076 273628 51088
rect 273680 51076 273686 51128
rect 250070 51048 250076 51060
rect 250031 51020 250076 51048
rect 250070 51008 250076 51020
rect 250128 51008 250134 51060
rect 273530 51008 273536 51060
rect 273588 51008 273594 51060
rect 341337 50915 341395 50921
rect 341337 50881 341349 50915
rect 341383 50912 341395 50915
rect 341426 50912 341432 50924
rect 341383 50884 341432 50912
rect 341383 50881 341395 50884
rect 341337 50875 341395 50881
rect 341426 50872 341432 50884
rect 341484 50872 341490 50924
rect 2774 50124 2780 50176
rect 2832 50164 2838 50176
rect 4890 50164 4896 50176
rect 2832 50136 4896 50164
rect 2832 50124 2838 50136
rect 4890 50124 4896 50136
rect 4948 50124 4954 50176
rect 236270 48396 236276 48408
rect 236231 48368 236276 48396
rect 236270 48356 236276 48368
rect 236328 48356 236334 48408
rect 303890 48356 303896 48408
rect 303948 48356 303954 48408
rect 230750 48328 230756 48340
rect 230711 48300 230756 48328
rect 230750 48288 230756 48300
rect 230808 48288 230814 48340
rect 288710 48288 288716 48340
rect 288768 48328 288774 48340
rect 288986 48328 288992 48340
rect 288768 48300 288992 48328
rect 288768 48288 288774 48300
rect 288986 48288 288992 48300
rect 289044 48288 289050 48340
rect 295518 48328 295524 48340
rect 295479 48300 295524 48328
rect 295518 48288 295524 48300
rect 295576 48288 295582 48340
rect 303908 48272 303936 48356
rect 323302 48328 323308 48340
rect 323263 48300 323308 48328
rect 323302 48288 323308 48300
rect 323360 48288 323366 48340
rect 324682 48288 324688 48340
rect 324740 48328 324746 48340
rect 324774 48328 324780 48340
rect 324740 48300 324780 48328
rect 324740 48288 324746 48300
rect 324774 48288 324780 48300
rect 324832 48288 324838 48340
rect 358722 48328 358728 48340
rect 358683 48300 358728 48328
rect 358722 48288 358728 48300
rect 358780 48288 358786 48340
rect 367002 48328 367008 48340
rect 366963 48300 367008 48328
rect 367002 48288 367008 48300
rect 367060 48288 367066 48340
rect 389177 48331 389235 48337
rect 389177 48297 389189 48331
rect 389223 48328 389235 48331
rect 389266 48328 389272 48340
rect 389223 48300 389272 48328
rect 389223 48297 389235 48300
rect 389177 48291 389235 48297
rect 389266 48288 389272 48300
rect 389324 48288 389330 48340
rect 470594 48328 470600 48340
rect 470555 48300 470600 48328
rect 470594 48288 470600 48300
rect 470652 48288 470658 48340
rect 273530 48260 273536 48272
rect 273491 48232 273536 48260
rect 273530 48220 273536 48232
rect 273588 48220 273594 48272
rect 303890 48220 303896 48272
rect 303948 48220 303954 48272
rect 325878 48220 325884 48272
rect 325936 48220 325942 48272
rect 327166 48220 327172 48272
rect 327224 48260 327230 48272
rect 327350 48260 327356 48272
rect 327224 48232 327356 48260
rect 327224 48220 327230 48232
rect 327350 48220 327356 48232
rect 327408 48220 327414 48272
rect 325896 48192 325924 48220
rect 325970 48192 325976 48204
rect 325896 48164 325976 48192
rect 325970 48152 325976 48164
rect 326028 48152 326034 48204
rect 262766 47036 262772 47048
rect 262692 47008 262772 47036
rect 262692 46912 262720 47008
rect 262766 46996 262772 47008
rect 262824 46996 262830 47048
rect 268010 46968 268016 46980
rect 267752 46940 268016 46968
rect 267752 46912 267780 46940
rect 268010 46928 268016 46940
rect 268068 46928 268074 46980
rect 285950 46968 285956 46980
rect 285911 46940 285956 46968
rect 285950 46928 285956 46940
rect 286008 46928 286014 46980
rect 302510 46968 302516 46980
rect 302471 46940 302516 46968
rect 302510 46928 302516 46940
rect 302568 46928 302574 46980
rect 339681 46971 339739 46977
rect 339681 46937 339693 46971
rect 339727 46968 339739 46971
rect 339954 46968 339960 46980
rect 339727 46940 339960 46968
rect 339727 46937 339739 46940
rect 339681 46931 339739 46937
rect 339954 46928 339960 46940
rect 340012 46928 340018 46980
rect 358722 46968 358728 46980
rect 358683 46940 358728 46968
rect 358722 46928 358728 46940
rect 358780 46928 358786 46980
rect 236270 46900 236276 46912
rect 236231 46872 236276 46900
rect 236270 46860 236276 46872
rect 236328 46860 236334 46912
rect 247126 46900 247132 46912
rect 247087 46872 247132 46900
rect 247126 46860 247132 46872
rect 247184 46860 247190 46912
rect 250073 46903 250131 46909
rect 250073 46869 250085 46903
rect 250119 46900 250131 46903
rect 250162 46900 250168 46912
rect 250119 46872 250168 46900
rect 250119 46869 250131 46872
rect 250073 46863 250131 46869
rect 250162 46860 250168 46872
rect 250220 46860 250226 46912
rect 251358 46900 251364 46912
rect 251319 46872 251364 46900
rect 251358 46860 251364 46872
rect 251416 46860 251422 46912
rect 262674 46860 262680 46912
rect 262732 46860 262738 46912
rect 267734 46860 267740 46912
rect 267792 46860 267798 46912
rect 306742 46860 306748 46912
rect 306800 46860 306806 46912
rect 323302 46900 323308 46912
rect 323263 46872 323308 46900
rect 323302 46860 323308 46872
rect 323360 46860 323366 46912
rect 324685 46903 324743 46909
rect 324685 46869 324697 46903
rect 324731 46900 324743 46903
rect 324774 46900 324780 46912
rect 324731 46872 324780 46900
rect 324731 46869 324743 46872
rect 324685 46863 324743 46869
rect 324774 46860 324780 46872
rect 324832 46860 324838 46912
rect 325970 46860 325976 46912
rect 326028 46900 326034 46912
rect 326062 46900 326068 46912
rect 326028 46872 326068 46900
rect 326028 46860 326034 46872
rect 326062 46860 326068 46872
rect 326120 46860 326126 46912
rect 327350 46900 327356 46912
rect 327311 46872 327356 46900
rect 327350 46860 327356 46872
rect 327408 46860 327414 46912
rect 330110 46900 330116 46912
rect 330071 46872 330116 46900
rect 330110 46860 330116 46872
rect 330168 46860 330174 46912
rect 338482 46860 338488 46912
rect 338540 46900 338546 46912
rect 338942 46900 338948 46912
rect 338540 46872 338948 46900
rect 338540 46860 338546 46872
rect 338942 46860 338948 46872
rect 339000 46860 339006 46912
rect 296806 46832 296812 46844
rect 296767 46804 296812 46832
rect 296806 46792 296812 46804
rect 296864 46792 296870 46844
rect 306760 46832 306788 46860
rect 306834 46832 306840 46844
rect 306760 46804 306840 46832
rect 306834 46792 306840 46804
rect 306892 46792 306898 46844
rect 294230 45500 294236 45552
rect 294288 45540 294294 45552
rect 294414 45540 294420 45552
rect 294288 45512 294420 45540
rect 294288 45500 294294 45512
rect 294414 45500 294420 45512
rect 294472 45500 294478 45552
rect 310882 45500 310888 45552
rect 310940 45540 310946 45552
rect 311066 45540 311072 45552
rect 310940 45512 311072 45540
rect 310940 45500 310946 45512
rect 311066 45500 311072 45512
rect 311124 45500 311130 45552
rect 317506 45500 317512 45552
rect 317564 45540 317570 45552
rect 317690 45540 317696 45552
rect 317564 45512 317696 45540
rect 317564 45500 317570 45512
rect 317690 45500 317696 45512
rect 317748 45500 317754 45552
rect 338482 45540 338488 45552
rect 338443 45512 338488 45540
rect 338482 45500 338488 45512
rect 338540 45500 338546 45552
rect 284662 44684 284668 44736
rect 284720 44724 284726 44736
rect 284757 44727 284815 44733
rect 284757 44724 284769 44727
rect 284720 44696 284769 44724
rect 284720 44684 284726 44696
rect 284757 44693 284769 44696
rect 284803 44693 284815 44727
rect 284757 44687 284815 44693
rect 266630 44140 266636 44192
rect 266688 44180 266694 44192
rect 266906 44180 266912 44192
rect 266688 44152 266912 44180
rect 266688 44140 266694 44152
rect 266906 44140 266912 44152
rect 266964 44140 266970 44192
rect 272150 44140 272156 44192
rect 272208 44180 272214 44192
rect 272426 44180 272432 44192
rect 272208 44152 272432 44180
rect 272208 44140 272214 44152
rect 272426 44140 272432 44152
rect 272484 44140 272490 44192
rect 296809 43979 296867 43985
rect 296809 43945 296821 43979
rect 296855 43976 296867 43979
rect 296898 43976 296904 43988
rect 296855 43948 296904 43976
rect 296855 43945 296867 43948
rect 296809 43939 296867 43945
rect 296898 43936 296904 43948
rect 296956 43936 296962 43988
rect 270678 42848 270684 42900
rect 270736 42888 270742 42900
rect 270865 42891 270923 42897
rect 270865 42888 270877 42891
rect 270736 42860 270877 42888
rect 270736 42848 270742 42860
rect 270865 42857 270877 42860
rect 270911 42857 270923 42891
rect 270865 42851 270923 42857
rect 303801 42075 303859 42081
rect 303801 42041 303813 42075
rect 303847 42072 303859 42075
rect 303890 42072 303896 42084
rect 303847 42044 303896 42072
rect 303847 42041 303859 42044
rect 303801 42035 303859 42041
rect 303890 42032 303896 42044
rect 303948 42032 303954 42084
rect 265250 41460 265256 41472
rect 265211 41432 265256 41460
rect 265250 41420 265256 41432
rect 265308 41420 265314 41472
rect 341426 41460 341432 41472
rect 341387 41432 341432 41460
rect 341426 41420 341432 41432
rect 341484 41420 341490 41472
rect 266630 41392 266636 41404
rect 266591 41364 266636 41392
rect 266630 41352 266636 41364
rect 266688 41352 266694 41404
rect 360286 41352 360292 41404
rect 360344 41392 360350 41404
rect 360470 41392 360476 41404
rect 360344 41364 360476 41392
rect 360344 41352 360350 41364
rect 360470 41352 360476 41364
rect 360528 41352 360534 41404
rect 377122 41324 377128 41336
rect 377083 41296 377128 41324
rect 377122 41284 377128 41296
rect 377180 41284 377186 41336
rect 241422 40264 241428 40316
rect 241480 40304 241486 40316
rect 245010 40304 245016 40316
rect 241480 40276 245016 40304
rect 241480 40264 241486 40276
rect 245010 40264 245016 40276
rect 245068 40264 245074 40316
rect 417878 40196 417884 40248
rect 417936 40236 417942 40248
rect 420362 40236 420368 40248
rect 417936 40208 420368 40236
rect 417936 40196 417942 40208
rect 420362 40196 420368 40208
rect 420420 40196 420426 40248
rect 437198 40196 437204 40248
rect 437256 40236 437262 40248
rect 437474 40236 437480 40248
rect 437256 40208 437480 40236
rect 437256 40196 437262 40208
rect 437474 40196 437480 40208
rect 437532 40196 437538 40248
rect 456518 40128 456524 40180
rect 456576 40168 456582 40180
rect 456886 40168 456892 40180
rect 456576 40140 456892 40168
rect 456576 40128 456582 40140
rect 456886 40128 456892 40140
rect 456944 40128 456950 40180
rect 253842 40060 253848 40112
rect 253900 40100 253906 40112
rect 262858 40100 262864 40112
rect 253900 40072 262864 40100
rect 253900 40060 253906 40072
rect 262858 40060 262864 40072
rect 262916 40060 262922 40112
rect 230750 38740 230756 38752
rect 230711 38712 230756 38740
rect 230750 38700 230756 38712
rect 230808 38700 230814 38752
rect 232222 38740 232228 38752
rect 232183 38712 232228 38740
rect 232222 38700 232228 38712
rect 232280 38700 232286 38752
rect 377030 38700 377036 38752
rect 377088 38740 377094 38752
rect 377125 38743 377183 38749
rect 377125 38740 377137 38743
rect 377088 38712 377137 38740
rect 377088 38700 377094 38712
rect 377125 38709 377137 38712
rect 377171 38709 377183 38743
rect 377125 38703 377183 38709
rect 273530 38672 273536 38684
rect 273491 38644 273536 38672
rect 273530 38632 273536 38644
rect 273588 38632 273594 38684
rect 295518 38632 295524 38684
rect 295576 38632 295582 38684
rect 295536 38536 295564 38632
rect 341426 38604 341432 38616
rect 341387 38576 341432 38604
rect 341426 38564 341432 38576
rect 341484 38564 341490 38616
rect 367002 38604 367008 38616
rect 366963 38576 367008 38604
rect 367002 38564 367008 38576
rect 367060 38564 367066 38616
rect 377122 38564 377128 38616
rect 377180 38604 377186 38616
rect 377306 38604 377312 38616
rect 377180 38576 377312 38604
rect 377180 38564 377186 38576
rect 377306 38564 377312 38576
rect 377364 38564 377370 38616
rect 295610 38536 295616 38548
rect 295536 38508 295616 38536
rect 295610 38496 295616 38508
rect 295668 38496 295674 38548
rect 327350 38536 327356 38548
rect 327311 38508 327356 38536
rect 327350 38496 327356 38508
rect 327408 38496 327414 38548
rect 286042 37380 286048 37392
rect 285968 37352 286048 37380
rect 285968 37324 285996 37352
rect 286042 37340 286048 37352
rect 286100 37340 286106 37392
rect 299845 37383 299903 37389
rect 299845 37349 299857 37383
rect 299891 37380 299903 37383
rect 300026 37380 300032 37392
rect 299891 37352 300032 37380
rect 299891 37349 299903 37352
rect 299845 37343 299903 37349
rect 300026 37340 300032 37352
rect 300084 37340 300090 37392
rect 230750 37312 230756 37324
rect 230711 37284 230756 37312
rect 230750 37272 230756 37284
rect 230808 37272 230814 37324
rect 236273 37315 236331 37321
rect 236273 37281 236285 37315
rect 236319 37312 236331 37315
rect 236454 37312 236460 37324
rect 236319 37284 236460 37312
rect 236319 37281 236331 37284
rect 236273 37275 236331 37281
rect 236454 37272 236460 37284
rect 236512 37272 236518 37324
rect 250070 37312 250076 37324
rect 250031 37284 250076 37312
rect 250070 37272 250076 37284
rect 250128 37272 250134 37324
rect 251361 37315 251419 37321
rect 251361 37281 251373 37315
rect 251407 37312 251419 37315
rect 251450 37312 251456 37324
rect 251407 37284 251456 37312
rect 251407 37281 251419 37284
rect 251361 37275 251419 37281
rect 251450 37272 251456 37284
rect 251508 37272 251514 37324
rect 285950 37272 285956 37324
rect 286008 37272 286014 37324
rect 323302 37312 323308 37324
rect 323263 37284 323308 37312
rect 323302 37272 323308 37284
rect 323360 37272 323366 37324
rect 324682 37312 324688 37324
rect 324643 37284 324688 37312
rect 324682 37272 324688 37284
rect 324740 37272 324746 37324
rect 330110 37312 330116 37324
rect 330071 37284 330116 37312
rect 330110 37272 330116 37284
rect 330168 37272 330174 37324
rect 339770 37272 339776 37324
rect 339828 37312 339834 37324
rect 339954 37312 339960 37324
rect 339828 37284 339960 37312
rect 339828 37272 339834 37284
rect 339954 37272 339960 37284
rect 340012 37272 340018 37324
rect 358722 37272 358728 37324
rect 358780 37312 358786 37324
rect 358814 37312 358820 37324
rect 358780 37284 358820 37312
rect 358780 37272 358786 37284
rect 358814 37272 358820 37284
rect 358872 37272 358878 37324
rect 288710 37244 288716 37256
rect 288671 37216 288716 37244
rect 288710 37204 288716 37216
rect 288768 37204 288774 37256
rect 265250 35952 265256 35964
rect 265211 35924 265256 35952
rect 265250 35912 265256 35924
rect 265308 35912 265314 35964
rect 3142 35844 3148 35896
rect 3200 35884 3206 35896
rect 6178 35884 6184 35896
rect 3200 35856 6184 35884
rect 3200 35844 3206 35856
rect 6178 35844 6184 35856
rect 6236 35844 6242 35896
rect 251450 35884 251456 35896
rect 251411 35856 251456 35884
rect 251450 35844 251456 35856
rect 251508 35844 251514 35896
rect 244366 34484 244372 34536
rect 244424 34524 244430 34536
rect 244550 34524 244556 34536
rect 244424 34496 244556 34524
rect 244424 34484 244430 34496
rect 244550 34484 244556 34496
rect 244608 34484 244614 34536
rect 247126 34524 247132 34536
rect 247087 34496 247132 34524
rect 247126 34484 247132 34496
rect 247184 34484 247190 34536
rect 272242 34484 272248 34536
rect 272300 34524 272306 34536
rect 272426 34524 272432 34536
rect 272300 34496 272432 34524
rect 272300 34484 272306 34496
rect 272426 34484 272432 34496
rect 272484 34484 272490 34536
rect 266630 34456 266636 34468
rect 266591 34428 266636 34456
rect 266630 34416 266636 34428
rect 266688 34416 266694 34468
rect 303801 32419 303859 32425
rect 303801 32385 303813 32419
rect 303847 32416 303859 32419
rect 303890 32416 303896 32428
rect 303847 32388 303896 32416
rect 303847 32385 303859 32388
rect 303801 32379 303859 32385
rect 303890 32376 303896 32388
rect 303948 32376 303954 32428
rect 372706 31872 372712 31884
rect 372667 31844 372712 31872
rect 372706 31832 372712 31844
rect 372764 31832 372770 31884
rect 239122 31804 239128 31816
rect 239048 31776 239128 31804
rect 239048 31748 239076 31776
rect 239122 31764 239128 31776
rect 239180 31764 239186 31816
rect 317506 31764 317512 31816
rect 317564 31804 317570 31816
rect 317690 31804 317696 31816
rect 317564 31776 317696 31804
rect 317564 31764 317570 31776
rect 317690 31764 317696 31776
rect 317748 31764 317754 31816
rect 360470 31804 360476 31816
rect 360304 31776 360476 31804
rect 360304 31748 360332 31776
rect 360470 31764 360476 31776
rect 360528 31764 360534 31816
rect 389358 31764 389364 31816
rect 389416 31764 389422 31816
rect 239030 31696 239036 31748
rect 239088 31696 239094 31748
rect 360286 31696 360292 31748
rect 360344 31696 360350 31748
rect 389376 31668 389404 31764
rect 389450 31668 389456 31680
rect 389376 31640 389456 31668
rect 389450 31628 389456 31640
rect 389508 31628 389514 31680
rect 248414 29180 248420 29232
rect 248472 29220 248478 29232
rect 257890 29220 257896 29232
rect 248472 29192 257896 29220
rect 248472 29180 248478 29192
rect 257890 29180 257896 29192
rect 257948 29180 257954 29232
rect 417878 29180 417884 29232
rect 417936 29220 417942 29232
rect 418798 29220 418804 29232
rect 417936 29192 418804 29220
rect 417936 29180 417942 29192
rect 418798 29180 418804 29192
rect 418856 29180 418862 29232
rect 456518 29180 456524 29232
rect 456576 29220 456582 29232
rect 456978 29220 456984 29232
rect 456576 29192 456984 29220
rect 456576 29180 456582 29192
rect 456978 29180 456984 29192
rect 457036 29180 457042 29232
rect 437198 29112 437204 29164
rect 437256 29152 437262 29164
rect 437474 29152 437480 29164
rect 437256 29124 437480 29152
rect 437256 29112 437262 29124
rect 437474 29112 437480 29124
rect 437532 29112 437538 29164
rect 301314 29084 301320 29096
rect 301240 29056 301320 29084
rect 284754 29016 284760 29028
rect 284715 28988 284760 29016
rect 284754 28976 284760 28988
rect 284812 28976 284818 29028
rect 285950 28976 285956 29028
rect 286008 29016 286014 29028
rect 286042 29016 286048 29028
rect 286008 28988 286048 29016
rect 286008 28976 286014 28988
rect 286042 28976 286048 28988
rect 286100 28976 286106 29028
rect 295518 28976 295524 29028
rect 295576 29016 295582 29028
rect 295610 29016 295616 29028
rect 295576 28988 295616 29016
rect 295576 28976 295582 28988
rect 295610 28976 295616 28988
rect 295668 28976 295674 29028
rect 301240 28960 301268 29056
rect 301314 29044 301320 29056
rect 301372 29044 301378 29096
rect 367002 29084 367008 29096
rect 366963 29056 367008 29084
rect 367002 29044 367008 29056
rect 367060 29044 367066 29096
rect 367094 29044 367100 29096
rect 367152 29084 367158 29096
rect 376662 29084 376668 29096
rect 367152 29056 376668 29084
rect 367152 29044 367158 29056
rect 376662 29044 376668 29056
rect 376720 29044 376726 29096
rect 492766 29044 492772 29096
rect 492824 29084 492830 29096
rect 502242 29084 502248 29096
rect 492824 29056 502248 29084
rect 492824 29044 492830 29056
rect 502242 29044 502248 29056
rect 502300 29044 502306 29096
rect 327166 28976 327172 29028
rect 327224 29016 327230 29028
rect 327350 29016 327356 29028
rect 327224 28988 327356 29016
rect 327224 28976 327230 28988
rect 327350 28976 327356 28988
rect 327408 28976 327414 29028
rect 341150 28976 341156 29028
rect 341208 29016 341214 29028
rect 341426 29016 341432 29028
rect 341208 28988 341432 29016
rect 341208 28976 341214 28988
rect 341426 28976 341432 28988
rect 341484 28976 341490 29028
rect 372706 29016 372712 29028
rect 372667 28988 372712 29016
rect 372706 28976 372712 28988
rect 372764 28976 372770 29028
rect 232222 28908 232228 28960
rect 232280 28948 232286 28960
rect 232314 28948 232320 28960
rect 232280 28920 232320 28948
rect 232280 28908 232286 28920
rect 232314 28908 232320 28920
rect 232372 28908 232378 28960
rect 236362 28948 236368 28960
rect 236323 28920 236368 28948
rect 236362 28908 236368 28920
rect 236420 28908 236426 28960
rect 301222 28908 301228 28960
rect 301280 28908 301286 28960
rect 323210 28908 323216 28960
rect 323268 28948 323274 28960
rect 323394 28948 323400 28960
rect 323268 28920 323400 28948
rect 323268 28908 323274 28920
rect 323394 28908 323400 28920
rect 323452 28908 323458 28960
rect 357618 28908 357624 28960
rect 357676 28948 357682 28960
rect 357802 28948 357808 28960
rect 357676 28920 357808 28948
rect 357676 28908 357682 28920
rect 357802 28908 357808 28920
rect 357860 28908 357866 28960
rect 367002 28948 367008 28960
rect 366963 28920 367008 28948
rect 367002 28908 367008 28920
rect 367060 28908 367066 28960
rect 375834 28948 375840 28960
rect 375795 28920 375840 28948
rect 375834 28908 375840 28920
rect 375892 28908 375898 28960
rect 377122 28948 377128 28960
rect 377083 28920 377128 28948
rect 377122 28908 377128 28920
rect 377180 28908 377186 28960
rect 307662 28840 307668 28892
rect 307720 28880 307726 28892
rect 315942 28880 315948 28892
rect 307720 28852 315948 28880
rect 307720 28840 307726 28852
rect 315942 28840 315948 28852
rect 316000 28840 316006 28892
rect 259730 27616 259736 27668
rect 259788 27656 259794 27668
rect 259822 27656 259828 27668
rect 259788 27628 259828 27656
rect 259788 27616 259794 27628
rect 259822 27616 259828 27628
rect 259880 27616 259886 27668
rect 288713 27659 288771 27665
rect 288713 27625 288725 27659
rect 288759 27656 288771 27659
rect 288802 27656 288808 27668
rect 288759 27628 288808 27656
rect 288759 27625 288771 27628
rect 288713 27619 288771 27625
rect 288802 27616 288808 27628
rect 288860 27616 288866 27668
rect 338485 27659 338543 27665
rect 338485 27625 338497 27659
rect 338531 27656 338543 27659
rect 338666 27656 338672 27668
rect 338531 27628 338672 27656
rect 338531 27625 338543 27628
rect 338485 27619 338543 27625
rect 338666 27616 338672 27628
rect 338724 27616 338730 27668
rect 265161 27591 265219 27597
rect 265161 27557 265173 27591
rect 265207 27588 265219 27591
rect 265250 27588 265256 27600
rect 265207 27560 265256 27588
rect 265207 27557 265219 27560
rect 265161 27551 265219 27557
rect 265250 27548 265256 27560
rect 265308 27548 265314 27600
rect 285953 27591 286011 27597
rect 285953 27557 285965 27591
rect 285999 27588 286011 27591
rect 286042 27588 286048 27600
rect 285999 27560 286048 27588
rect 285999 27557 286011 27560
rect 285953 27551 286011 27557
rect 286042 27548 286048 27560
rect 286100 27548 286106 27600
rect 295518 27588 295524 27600
rect 295479 27560 295524 27588
rect 295518 27548 295524 27560
rect 295576 27548 295582 27600
rect 330113 27591 330171 27597
rect 330113 27557 330125 27591
rect 330159 27588 330171 27591
rect 330202 27588 330208 27600
rect 330159 27560 330208 27588
rect 330159 27557 330171 27560
rect 330113 27551 330171 27557
rect 330202 27548 330208 27560
rect 330260 27548 330266 27600
rect 358541 27591 358599 27597
rect 358541 27557 358553 27591
rect 358587 27588 358599 27591
rect 358630 27588 358636 27600
rect 358587 27560 358636 27588
rect 358587 27557 358599 27560
rect 358541 27551 358599 27557
rect 358630 27548 358636 27560
rect 358688 27548 358694 27600
rect 301133 27523 301191 27529
rect 301133 27489 301145 27523
rect 301179 27520 301191 27523
rect 301222 27520 301228 27532
rect 301179 27492 301228 27520
rect 301179 27489 301191 27492
rect 301133 27483 301191 27489
rect 301222 27480 301228 27492
rect 301280 27480 301286 27532
rect 247034 26324 247040 26376
rect 247092 26364 247098 26376
rect 247126 26364 247132 26376
rect 247092 26336 247132 26364
rect 247092 26324 247098 26336
rect 247126 26324 247132 26336
rect 247184 26324 247190 26376
rect 251450 26296 251456 26308
rect 251411 26268 251456 26296
rect 251450 26256 251456 26268
rect 251508 26256 251514 26308
rect 249978 26188 249984 26240
rect 250036 26228 250042 26240
rect 250162 26228 250168 26240
rect 250036 26200 250168 26228
rect 250036 26188 250042 26200
rect 250162 26188 250168 26200
rect 250220 26188 250226 26240
rect 288802 26228 288808 26240
rect 288763 26200 288808 26228
rect 288802 26188 288808 26200
rect 288860 26188 288866 26240
rect 310882 26228 310888 26240
rect 310843 26200 310888 26228
rect 310882 26188 310888 26200
rect 310940 26188 310946 26240
rect 266722 24936 266728 24948
rect 266648 24908 266728 24936
rect 266648 24812 266676 24908
rect 266722 24896 266728 24908
rect 266780 24896 266786 24948
rect 244369 24803 244427 24809
rect 244369 24769 244381 24803
rect 244415 24800 244427 24803
rect 244458 24800 244464 24812
rect 244415 24772 244464 24800
rect 244415 24769 244427 24772
rect 244369 24763 244427 24769
rect 244458 24760 244464 24772
rect 244516 24760 244522 24812
rect 266630 24760 266636 24812
rect 266688 24760 266694 24812
rect 337105 24327 337163 24333
rect 337105 24293 337117 24327
rect 337151 24324 337163 24327
rect 337194 24324 337200 24336
rect 337151 24296 337200 24324
rect 337151 24293 337163 24296
rect 337105 24287 337163 24293
rect 337194 24284 337200 24296
rect 337252 24284 337258 24336
rect 270494 22176 270500 22228
rect 270552 22216 270558 22228
rect 270770 22216 270776 22228
rect 270552 22188 270776 22216
rect 270552 22176 270558 22188
rect 270770 22176 270776 22188
rect 270828 22176 270834 22228
rect 247218 22148 247224 22160
rect 247144 22120 247224 22148
rect 247144 22092 247172 22120
rect 247218 22108 247224 22120
rect 247276 22108 247282 22160
rect 268010 22108 268016 22160
rect 268068 22148 268074 22160
rect 272242 22148 272248 22160
rect 268068 22120 272248 22148
rect 268068 22108 268074 22120
rect 272242 22108 272248 22120
rect 272300 22108 272306 22160
rect 374362 22108 374368 22160
rect 374420 22108 374426 22160
rect 247126 22040 247132 22092
rect 247184 22040 247190 22092
rect 372706 22040 372712 22092
rect 372764 22040 372770 22092
rect 372724 22012 372752 22040
rect 374380 22024 374408 22108
rect 377122 22080 377128 22092
rect 377083 22052 377128 22080
rect 377122 22040 377128 22052
rect 377180 22040 377186 22092
rect 372798 22012 372804 22024
rect 372724 21984 372804 22012
rect 372798 21972 372804 21984
rect 372856 21972 372862 22024
rect 374362 21972 374368 22024
rect 374420 21972 374426 22024
rect 239030 19388 239036 19440
rect 239088 19388 239094 19440
rect 236362 19360 236368 19372
rect 236323 19332 236368 19360
rect 236362 19320 236368 19332
rect 236420 19320 236426 19372
rect 239048 19304 239076 19388
rect 302510 19320 302516 19372
rect 302568 19360 302574 19372
rect 302602 19360 302608 19372
rect 302568 19332 302608 19360
rect 302568 19320 302574 19332
rect 302602 19320 302608 19332
rect 302660 19320 302666 19372
rect 306742 19320 306748 19372
rect 306800 19360 306806 19372
rect 306834 19360 306840 19372
rect 306800 19332 306840 19360
rect 306800 19320 306806 19332
rect 306834 19320 306840 19332
rect 306892 19320 306898 19372
rect 337102 19360 337108 19372
rect 337063 19332 337108 19360
rect 337102 19320 337108 19332
rect 337160 19320 337166 19372
rect 338666 19320 338672 19372
rect 338724 19360 338730 19372
rect 338850 19360 338856 19372
rect 338724 19332 338856 19360
rect 338724 19320 338730 19332
rect 338850 19320 338856 19332
rect 338908 19320 338914 19372
rect 367002 19360 367008 19372
rect 366963 19332 367008 19360
rect 367002 19320 367008 19332
rect 367060 19320 367066 19372
rect 375834 19360 375840 19372
rect 375795 19332 375840 19360
rect 375834 19320 375840 19332
rect 375892 19320 375898 19372
rect 239030 19252 239036 19304
rect 239088 19252 239094 19304
rect 366910 19292 366916 19304
rect 366871 19264 366916 19292
rect 366910 19252 366916 19264
rect 366968 19252 366974 19304
rect 366818 19184 366824 19236
rect 366876 19224 366882 19236
rect 367002 19224 367008 19236
rect 366876 19196 367008 19224
rect 366876 19184 366882 19196
rect 367002 19184 367008 19196
rect 367060 19184 367066 19236
rect 267826 18068 267832 18080
rect 267752 18040 267832 18068
rect 267752 18012 267780 18040
rect 267826 18028 267832 18040
rect 267884 18028 267890 18080
rect 284846 18068 284852 18080
rect 284680 18040 284852 18068
rect 284680 18012 284708 18040
rect 284846 18028 284852 18040
rect 284904 18028 284910 18080
rect 265158 18000 265164 18012
rect 265119 17972 265164 18000
rect 265158 17960 265164 17972
rect 265216 17960 265222 18012
rect 267734 17960 267740 18012
rect 267792 17960 267798 18012
rect 284662 17960 284668 18012
rect 284720 17960 284726 18012
rect 285950 18000 285956 18012
rect 285911 17972 285956 18000
rect 285950 17960 285956 17972
rect 286008 17960 286014 18012
rect 299842 18000 299848 18012
rect 299803 17972 299848 18000
rect 299842 17960 299848 17972
rect 299900 17960 299906 18012
rect 301130 18000 301136 18012
rect 301091 17972 301136 18000
rect 301130 17960 301136 17972
rect 301188 17960 301194 18012
rect 324498 17960 324504 18012
rect 324556 18000 324562 18012
rect 324682 18000 324688 18012
rect 324556 17972 324688 18000
rect 324556 17960 324562 17972
rect 324682 17960 324688 17972
rect 324740 17960 324746 18012
rect 327258 17932 327264 17944
rect 327219 17904 327264 17932
rect 327258 17892 327264 17904
rect 327316 17892 327322 17944
rect 389358 17932 389364 17944
rect 389319 17904 389364 17932
rect 389358 17892 389364 17904
rect 389416 17892 389422 17944
rect 456518 16804 456524 16856
rect 456576 16844 456582 16856
rect 458818 16844 458824 16856
rect 456576 16816 458824 16844
rect 456576 16804 456582 16816
rect 458818 16804 458824 16816
rect 458876 16804 458882 16856
rect 417878 16736 417884 16788
rect 417936 16776 417942 16788
rect 418154 16776 418160 16788
rect 417936 16748 418160 16776
rect 417936 16736 417942 16748
rect 418154 16736 418160 16748
rect 418212 16736 418218 16788
rect 437198 16736 437204 16788
rect 437256 16776 437262 16788
rect 437474 16776 437480 16788
rect 437256 16748 437480 16776
rect 437256 16736 437262 16748
rect 437474 16736 437480 16748
rect 437532 16736 437538 16788
rect 336734 16668 336740 16720
rect 336792 16708 336798 16720
rect 338206 16708 338212 16720
rect 336792 16680 338212 16708
rect 336792 16668 336798 16680
rect 338206 16668 338212 16680
rect 338264 16668 338270 16720
rect 251082 16600 251088 16652
rect 251140 16640 251146 16652
rect 259362 16640 259368 16652
rect 251140 16612 259368 16640
rect 251140 16600 251146 16612
rect 259362 16600 259368 16612
rect 259420 16600 259426 16652
rect 270586 16600 270592 16652
rect 270644 16600 270650 16652
rect 288802 16600 288808 16652
rect 288860 16640 288866 16652
rect 310882 16640 310888 16652
rect 288860 16612 288905 16640
rect 310843 16612 310888 16640
rect 288860 16600 288866 16612
rect 310882 16600 310888 16612
rect 310940 16600 310946 16652
rect 270604 16516 270632 16600
rect 273438 16572 273444 16584
rect 273399 16544 273444 16572
rect 273438 16532 273444 16544
rect 273496 16532 273502 16584
rect 270586 16464 270592 16516
rect 270644 16464 270650 16516
rect 114462 15104 114468 15156
rect 114520 15144 114526 15156
rect 276106 15144 276112 15156
rect 114520 15116 276112 15144
rect 114520 15104 114526 15116
rect 276106 15104 276112 15116
rect 276164 15104 276170 15156
rect 110322 15036 110328 15088
rect 110380 15076 110386 15088
rect 274726 15076 274732 15088
rect 110380 15048 274732 15076
rect 110380 15036 110386 15048
rect 274726 15036 274732 15048
rect 274784 15036 274790 15088
rect 107470 14968 107476 15020
rect 107528 15008 107534 15020
rect 273346 15008 273352 15020
rect 107528 14980 273352 15008
rect 107528 14968 107534 14980
rect 273346 14968 273352 14980
rect 273404 14968 273410 15020
rect 103422 14900 103428 14952
rect 103480 14940 103486 14952
rect 271966 14940 271972 14952
rect 103480 14912 271972 14940
rect 103480 14900 103486 14912
rect 271966 14900 271972 14912
rect 272024 14900 272030 14952
rect 99282 14832 99288 14884
rect 99340 14872 99346 14884
rect 270586 14872 270592 14884
rect 99340 14844 270592 14872
rect 99340 14832 99346 14844
rect 270586 14832 270592 14844
rect 270644 14832 270650 14884
rect 96522 14764 96528 14816
rect 96580 14804 96586 14816
rect 269206 14804 269212 14816
rect 96580 14776 269212 14804
rect 96580 14764 96586 14776
rect 269206 14764 269212 14776
rect 269264 14764 269270 14816
rect 92382 14696 92388 14748
rect 92440 14736 92446 14748
rect 266446 14736 266452 14748
rect 92440 14708 266452 14736
rect 92440 14696 92446 14708
rect 266446 14696 266452 14708
rect 266504 14696 266510 14748
rect 89622 14628 89628 14680
rect 89680 14668 89686 14680
rect 265066 14668 265072 14680
rect 89680 14640 265072 14668
rect 89680 14628 89686 14640
rect 265066 14628 265072 14640
rect 265124 14628 265130 14680
rect 85482 14560 85488 14612
rect 85540 14600 85546 14612
rect 263686 14600 263692 14612
rect 85540 14572 263692 14600
rect 85540 14560 85546 14572
rect 263686 14560 263692 14572
rect 263744 14560 263750 14612
rect 82722 14492 82728 14544
rect 82780 14532 82786 14544
rect 262582 14532 262588 14544
rect 82780 14504 262588 14532
rect 82780 14492 82786 14504
rect 262582 14492 262588 14504
rect 262640 14492 262646 14544
rect 78582 14424 78588 14476
rect 78640 14464 78646 14476
rect 260926 14464 260932 14476
rect 78640 14436 260932 14464
rect 78640 14424 78646 14436
rect 260926 14424 260932 14436
rect 260984 14424 260990 14476
rect 117222 14356 117228 14408
rect 117280 14396 117286 14408
rect 277670 14396 277676 14408
rect 117280 14368 277676 14396
rect 117280 14356 117286 14368
rect 277670 14356 277676 14368
rect 277728 14356 277734 14408
rect 121362 14288 121368 14340
rect 121420 14328 121426 14340
rect 278866 14328 278872 14340
rect 121420 14300 278872 14328
rect 121420 14288 121426 14300
rect 278866 14288 278872 14300
rect 278924 14288 278930 14340
rect 125410 14220 125416 14272
rect 125468 14260 125474 14272
rect 280246 14260 280252 14272
rect 125468 14232 280252 14260
rect 125468 14220 125474 14232
rect 280246 14220 280252 14232
rect 280304 14220 280310 14272
rect 186222 13744 186228 13796
rect 186280 13784 186286 13796
rect 306558 13784 306564 13796
rect 186280 13756 306564 13784
rect 186280 13744 186286 13756
rect 306558 13744 306564 13756
rect 306616 13744 306622 13796
rect 183462 13676 183468 13728
rect 183520 13716 183526 13728
rect 303890 13716 303896 13728
rect 183520 13688 303896 13716
rect 183520 13676 183526 13688
rect 303890 13676 303896 13688
rect 303948 13676 303954 13728
rect 179322 13608 179328 13660
rect 179380 13648 179386 13660
rect 302510 13648 302516 13660
rect 179380 13620 302516 13648
rect 179380 13608 179386 13620
rect 302510 13608 302516 13620
rect 302568 13608 302574 13660
rect 176562 13540 176568 13592
rect 176620 13580 176626 13592
rect 301130 13580 301136 13592
rect 176620 13552 301136 13580
rect 176620 13540 176626 13552
rect 301130 13540 301136 13552
rect 301188 13540 301194 13592
rect 172422 13472 172428 13524
rect 172480 13512 172486 13524
rect 299842 13512 299848 13524
rect 172480 13484 299848 13512
rect 172480 13472 172486 13484
rect 299842 13472 299848 13484
rect 299900 13472 299906 13524
rect 168282 13404 168288 13456
rect 168340 13444 168346 13456
rect 298278 13444 298284 13456
rect 168340 13416 298284 13444
rect 168340 13404 168346 13416
rect 298278 13404 298284 13416
rect 298336 13404 298342 13456
rect 165522 13336 165528 13388
rect 165580 13376 165586 13388
rect 296898 13376 296904 13388
rect 165580 13348 296904 13376
rect 165580 13336 165586 13348
rect 296898 13336 296904 13348
rect 296956 13336 296962 13388
rect 160002 13268 160008 13320
rect 160060 13308 160066 13320
rect 294230 13308 294236 13320
rect 160060 13280 294236 13308
rect 160060 13268 160066 13280
rect 294230 13268 294236 13280
rect 294288 13268 294294 13320
rect 74442 13200 74448 13252
rect 74500 13240 74506 13252
rect 259638 13240 259644 13252
rect 74500 13212 259644 13240
rect 74500 13200 74506 13212
rect 259638 13200 259644 13212
rect 259696 13200 259702 13252
rect 71682 13132 71688 13184
rect 71740 13172 71746 13184
rect 258166 13172 258172 13184
rect 71740 13144 258172 13172
rect 71740 13132 71746 13144
rect 258166 13132 258172 13144
rect 258224 13132 258230 13184
rect 31662 13064 31668 13116
rect 31720 13104 31726 13116
rect 241606 13104 241612 13116
rect 31720 13076 241612 13104
rect 31720 13064 31726 13076
rect 241606 13064 241612 13076
rect 241664 13064 241670 13116
rect 190362 12996 190368 13048
rect 190420 13036 190426 13048
rect 307938 13036 307944 13048
rect 190420 13008 307944 13036
rect 190420 12996 190426 13008
rect 307938 12996 307944 13008
rect 307996 12996 308002 13048
rect 206922 12928 206928 12980
rect 206980 12968 206986 12980
rect 314838 12968 314844 12980
rect 206980 12940 314844 12968
rect 206980 12928 206986 12940
rect 314838 12928 314844 12940
rect 314896 12928 314902 12980
rect 211062 12860 211068 12912
rect 211120 12900 211126 12912
rect 316218 12900 316224 12912
rect 211120 12872 316224 12900
rect 211120 12860 211126 12872
rect 316218 12860 316224 12872
rect 316276 12860 316282 12912
rect 213822 12792 213828 12844
rect 213880 12832 213886 12844
rect 317598 12832 317604 12844
rect 213880 12804 317604 12832
rect 213880 12792 213886 12804
rect 317598 12792 317604 12804
rect 317656 12792 317662 12844
rect 217962 12724 217968 12776
rect 218020 12764 218026 12776
rect 318978 12764 318984 12776
rect 218020 12736 318984 12764
rect 218020 12724 218026 12736
rect 318978 12724 318984 12736
rect 319036 12724 319042 12776
rect 220722 12656 220728 12708
rect 220780 12696 220786 12708
rect 320266 12696 320272 12708
rect 220780 12668 320272 12696
rect 220780 12656 220786 12668
rect 320266 12656 320272 12668
rect 320324 12656 320330 12708
rect 224862 12588 224868 12640
rect 224920 12628 224926 12640
rect 321738 12628 321744 12640
rect 224920 12600 321744 12628
rect 224920 12588 224926 12600
rect 321738 12588 321744 12600
rect 321796 12588 321802 12640
rect 229002 12520 229008 12572
rect 229060 12560 229066 12572
rect 323118 12560 323124 12572
rect 229060 12532 323124 12560
rect 229060 12520 229066 12532
rect 323118 12520 323124 12532
rect 323176 12520 323182 12572
rect 230661 12495 230719 12501
rect 230661 12461 230673 12495
rect 230707 12492 230719 12495
rect 230750 12492 230756 12504
rect 230707 12464 230756 12492
rect 230707 12461 230719 12464
rect 230661 12455 230719 12461
rect 230750 12452 230756 12464
rect 230808 12452 230814 12504
rect 323302 12492 323308 12504
rect 323136 12464 323308 12492
rect 323136 12436 323164 12464
rect 323302 12452 323308 12464
rect 323360 12452 323366 12504
rect 325970 12492 325976 12504
rect 325896 12464 325976 12492
rect 325896 12436 325924 12464
rect 325970 12452 325976 12464
rect 326028 12452 326034 12504
rect 337102 12492 337108 12504
rect 337028 12464 337108 12492
rect 337028 12436 337056 12464
rect 337102 12452 337108 12464
rect 337160 12452 337166 12504
rect 169662 12384 169668 12436
rect 169720 12424 169726 12436
rect 299566 12424 299572 12436
rect 169720 12396 299572 12424
rect 169720 12384 169726 12396
rect 299566 12384 299572 12396
rect 299624 12384 299630 12436
rect 323118 12384 323124 12436
rect 323176 12384 323182 12436
rect 325878 12384 325884 12436
rect 325936 12384 325942 12436
rect 337010 12384 337016 12436
rect 337068 12384 337074 12436
rect 166902 12316 166908 12368
rect 166960 12356 166966 12368
rect 298186 12356 298192 12368
rect 166960 12328 298192 12356
rect 166960 12316 166966 12328
rect 298186 12316 298192 12328
rect 298244 12316 298250 12368
rect 366910 12356 366916 12368
rect 366871 12328 366916 12356
rect 366910 12316 366916 12328
rect 366968 12316 366974 12368
rect 162762 12248 162768 12300
rect 162820 12288 162826 12300
rect 295521 12291 295579 12297
rect 295521 12288 295533 12291
rect 162820 12260 295533 12288
rect 162820 12248 162826 12260
rect 295521 12257 295533 12260
rect 295567 12257 295579 12291
rect 295521 12251 295579 12257
rect 155862 12180 155868 12232
rect 155920 12220 155926 12232
rect 292758 12220 292764 12232
rect 155920 12192 292764 12220
rect 155920 12180 155926 12192
rect 292758 12180 292764 12192
rect 292816 12180 292822 12232
rect 151722 12112 151728 12164
rect 151780 12152 151786 12164
rect 291470 12152 291476 12164
rect 151780 12124 291476 12152
rect 151780 12112 151786 12124
rect 291470 12112 291476 12124
rect 291528 12112 291534 12164
rect 148962 12044 148968 12096
rect 149020 12084 149026 12096
rect 289998 12084 290004 12096
rect 149020 12056 290004 12084
rect 149020 12044 149026 12056
rect 289998 12044 290004 12056
rect 290056 12044 290062 12096
rect 144822 11976 144828 12028
rect 144880 12016 144886 12028
rect 288802 12016 288808 12028
rect 144880 11988 288808 12016
rect 144880 11976 144886 11988
rect 288802 11976 288808 11988
rect 288860 11976 288866 12028
rect 142062 11908 142068 11960
rect 142120 11948 142126 11960
rect 287330 11948 287336 11960
rect 142120 11920 287336 11948
rect 142120 11908 142126 11920
rect 287330 11908 287336 11920
rect 287388 11908 287394 11960
rect 128262 11840 128268 11892
rect 128320 11880 128326 11892
rect 281534 11880 281540 11892
rect 128320 11852 281540 11880
rect 128320 11840 128326 11852
rect 281534 11840 281540 11852
rect 281592 11840 281598 11892
rect 126882 11772 126888 11824
rect 126940 11812 126946 11824
rect 281626 11812 281632 11824
rect 126940 11784 281632 11812
rect 126940 11772 126946 11784
rect 281626 11772 281632 11784
rect 281684 11772 281690 11824
rect 23382 11704 23388 11756
rect 23440 11744 23446 11756
rect 238938 11744 238944 11756
rect 23440 11716 238944 11744
rect 23440 11704 23446 11716
rect 238938 11704 238944 11716
rect 238996 11704 239002 11756
rect 173802 11636 173808 11688
rect 173860 11676 173866 11688
rect 300946 11676 300952 11688
rect 173860 11648 300952 11676
rect 173860 11636 173866 11648
rect 300946 11636 300952 11648
rect 301004 11636 301010 11688
rect 176470 11568 176476 11620
rect 176528 11608 176534 11620
rect 302326 11608 302332 11620
rect 176528 11580 302332 11608
rect 176528 11568 176534 11580
rect 302326 11568 302332 11580
rect 302384 11568 302390 11620
rect 180702 11500 180708 11552
rect 180760 11540 180766 11552
rect 303706 11540 303712 11552
rect 180760 11512 303712 11540
rect 180760 11500 180766 11512
rect 303706 11500 303712 11512
rect 303764 11500 303770 11552
rect 184842 11432 184848 11484
rect 184900 11472 184906 11484
rect 305086 11472 305092 11484
rect 184900 11444 305092 11472
rect 184900 11432 184906 11444
rect 305086 11432 305092 11444
rect 305144 11432 305150 11484
rect 187602 11364 187608 11416
rect 187660 11404 187666 11416
rect 306466 11404 306472 11416
rect 187660 11376 306472 11404
rect 187660 11364 187666 11376
rect 306466 11364 306472 11376
rect 306524 11364 306530 11416
rect 191742 11296 191748 11348
rect 191800 11336 191806 11348
rect 308030 11336 308036 11348
rect 191800 11308 308036 11336
rect 191800 11296 191806 11308
rect 308030 11296 308036 11308
rect 308088 11296 308094 11348
rect 194502 11228 194508 11280
rect 194560 11268 194566 11280
rect 309410 11268 309416 11280
rect 194560 11240 309416 11268
rect 194560 11228 194566 11240
rect 309410 11228 309416 11240
rect 309468 11228 309474 11280
rect 198642 11160 198648 11212
rect 198700 11200 198706 11212
rect 310882 11200 310888 11212
rect 198700 11172 310888 11200
rect 198700 11160 198706 11172
rect 310882 11160 310888 11172
rect 310940 11160 310946 11212
rect 230658 11132 230664 11144
rect 230619 11104 230664 11132
rect 230658 11092 230664 11104
rect 230716 11092 230722 11144
rect 113082 10956 113088 11008
rect 113140 10996 113146 11008
rect 276014 10996 276020 11008
rect 113140 10968 276020 10996
rect 113140 10956 113146 10968
rect 276014 10956 276020 10968
rect 276072 10956 276078 11008
rect 108942 10888 108948 10940
rect 109000 10928 109006 10940
rect 273441 10931 273499 10937
rect 273441 10928 273453 10931
rect 109000 10900 273453 10928
rect 109000 10888 109006 10900
rect 273441 10897 273453 10900
rect 273487 10897 273499 10931
rect 273441 10891 273499 10897
rect 106182 10820 106188 10872
rect 106240 10860 106246 10872
rect 268010 10860 268016 10872
rect 106240 10832 268016 10860
rect 106240 10820 106246 10832
rect 268010 10820 268016 10832
rect 268068 10820 268074 10872
rect 102042 10752 102048 10804
rect 102100 10792 102106 10804
rect 270494 10792 270500 10804
rect 102100 10764 270500 10792
rect 102100 10752 102106 10764
rect 270494 10752 270500 10764
rect 270552 10752 270558 10804
rect 99190 10684 99196 10736
rect 99248 10724 99254 10736
rect 269298 10724 269304 10736
rect 99248 10696 269304 10724
rect 99248 10684 99254 10696
rect 269298 10684 269304 10696
rect 269356 10684 269362 10736
rect 95142 10616 95148 10668
rect 95200 10656 95206 10668
rect 267734 10656 267740 10668
rect 95200 10628 267740 10656
rect 95200 10616 95206 10628
rect 267734 10616 267740 10628
rect 267792 10616 267798 10668
rect 91002 10548 91008 10600
rect 91060 10588 91066 10600
rect 266630 10588 266636 10600
rect 91060 10560 266636 10588
rect 91060 10548 91066 10560
rect 266630 10548 266636 10560
rect 266688 10548 266694 10600
rect 64782 10480 64788 10532
rect 64840 10520 64846 10532
rect 255590 10520 255596 10532
rect 64840 10492 255596 10520
rect 64840 10480 64846 10492
rect 255590 10480 255596 10492
rect 255648 10480 255654 10532
rect 60642 10412 60648 10464
rect 60700 10452 60706 10464
rect 254026 10452 254032 10464
rect 60700 10424 254032 10452
rect 60700 10412 60706 10424
rect 254026 10412 254032 10424
rect 254084 10412 254090 10464
rect 56502 10344 56508 10396
rect 56560 10384 56566 10396
rect 252646 10384 252652 10396
rect 56560 10356 252652 10384
rect 56560 10344 56566 10356
rect 252646 10344 252652 10356
rect 252704 10344 252710 10396
rect 53742 10276 53748 10328
rect 53800 10316 53806 10328
rect 251266 10316 251272 10328
rect 53800 10288 251272 10316
rect 53800 10276 53806 10288
rect 251266 10276 251272 10288
rect 251324 10276 251330 10328
rect 117130 10208 117136 10260
rect 117188 10248 117194 10260
rect 277578 10248 277584 10260
rect 117188 10220 277584 10248
rect 117188 10208 117194 10220
rect 277578 10208 277584 10220
rect 277636 10208 277642 10260
rect 119982 10140 119988 10192
rect 120040 10180 120046 10192
rect 278958 10180 278964 10192
rect 120040 10152 278964 10180
rect 120040 10140 120046 10152
rect 278958 10140 278964 10152
rect 279016 10140 279022 10192
rect 124122 10072 124128 10124
rect 124180 10112 124186 10124
rect 280338 10112 280344 10124
rect 124180 10084 280344 10112
rect 124180 10072 124186 10084
rect 280338 10072 280344 10084
rect 280396 10072 280402 10124
rect 143442 10004 143448 10056
rect 143500 10044 143506 10056
rect 288526 10044 288532 10056
rect 143500 10016 288532 10044
rect 143500 10004 143506 10016
rect 288526 10004 288532 10016
rect 288584 10004 288590 10056
rect 147582 9936 147588 9988
rect 147640 9976 147646 9988
rect 289814 9976 289820 9988
rect 147640 9948 289820 9976
rect 147640 9936 147646 9948
rect 289814 9936 289820 9948
rect 289872 9936 289878 9988
rect 151630 9868 151636 9920
rect 151688 9908 151694 9920
rect 291286 9908 291292 9920
rect 151688 9880 291292 9908
rect 151688 9868 151694 9880
rect 291286 9868 291292 9880
rect 291344 9868 291350 9920
rect 154482 9800 154488 9852
rect 154540 9840 154546 9852
rect 292850 9840 292856 9852
rect 154540 9812 292856 9840
rect 154540 9800 154546 9812
rect 292850 9800 292856 9812
rect 292908 9800 292914 9852
rect 158622 9732 158628 9784
rect 158680 9772 158686 9784
rect 294046 9772 294052 9784
rect 158680 9744 294052 9772
rect 158680 9732 158686 9744
rect 294046 9732 294052 9744
rect 294104 9732 294110 9784
rect 306742 9772 306748 9784
rect 306668 9744 306748 9772
rect 306668 9716 306696 9744
rect 306742 9732 306748 9744
rect 306800 9732 306806 9784
rect 161382 9664 161388 9716
rect 161440 9704 161446 9716
rect 295426 9704 295432 9716
rect 161440 9676 295432 9704
rect 161440 9664 161446 9676
rect 295426 9664 295432 9676
rect 295484 9664 295490 9716
rect 306650 9664 306656 9716
rect 306708 9664 306714 9716
rect 330110 9704 330116 9716
rect 330071 9676 330116 9704
rect 330110 9664 330116 9676
rect 330168 9664 330174 9716
rect 358538 9704 358544 9716
rect 358499 9676 358544 9704
rect 358538 9664 358544 9676
rect 358596 9664 358602 9716
rect 203886 9596 203892 9648
rect 203944 9636 203950 9648
rect 313366 9636 313372 9648
rect 203944 9608 313372 9636
rect 203944 9596 203950 9608
rect 313366 9596 313372 9608
rect 313424 9596 313430 9648
rect 327258 9636 327264 9648
rect 327219 9608 327264 9636
rect 327258 9596 327264 9608
rect 327316 9596 327322 9648
rect 200390 9528 200396 9580
rect 200448 9568 200454 9580
rect 311986 9568 311992 9580
rect 200448 9540 311992 9568
rect 200448 9528 200454 9540
rect 311986 9528 311992 9540
rect 312044 9528 312050 9580
rect 196802 9460 196808 9512
rect 196860 9500 196866 9512
rect 310606 9500 310612 9512
rect 196860 9472 310612 9500
rect 196860 9460 196866 9472
rect 310606 9460 310612 9472
rect 310664 9460 310670 9512
rect 193214 9392 193220 9444
rect 193272 9432 193278 9444
rect 309226 9432 309232 9444
rect 193272 9404 309232 9432
rect 193272 9392 193278 9404
rect 309226 9392 309232 9404
rect 309284 9392 309290 9444
rect 139670 9324 139676 9376
rect 139728 9364 139734 9376
rect 287146 9364 287152 9376
rect 139728 9336 287152 9364
rect 139728 9324 139734 9336
rect 287146 9324 287152 9336
rect 287204 9324 287210 9376
rect 136082 9256 136088 9308
rect 136140 9296 136146 9308
rect 285858 9296 285864 9308
rect 136140 9268 285864 9296
rect 136140 9256 136146 9268
rect 285858 9256 285864 9268
rect 285916 9256 285922 9308
rect 49326 9188 49332 9240
rect 49384 9228 49390 9240
rect 249886 9228 249892 9240
rect 49384 9200 249892 9228
rect 49384 9188 49390 9200
rect 249886 9188 249892 9200
rect 249944 9188 249950 9240
rect 253842 9188 253848 9240
rect 253900 9228 253906 9240
rect 334158 9228 334164 9240
rect 253900 9200 334164 9228
rect 253900 9188 253906 9200
rect 334158 9188 334164 9200
rect 334216 9188 334222 9240
rect 44542 9120 44548 9172
rect 44600 9160 44606 9172
rect 247126 9160 247132 9172
rect 44600 9132 247132 9160
rect 44600 9120 44606 9132
rect 247126 9120 247132 9132
rect 247184 9120 247190 9172
rect 250346 9120 250352 9172
rect 250404 9160 250410 9172
rect 332778 9160 332784 9172
rect 250404 9132 332784 9160
rect 250404 9120 250410 9132
rect 332778 9120 332784 9132
rect 332836 9120 332842 9172
rect 27890 9052 27896 9104
rect 27948 9092 27954 9104
rect 233878 9092 233884 9104
rect 27948 9064 233884 9092
rect 27948 9052 27954 9064
rect 233878 9052 233884 9064
rect 233936 9052 233942 9104
rect 243170 9052 243176 9104
rect 243228 9092 243234 9104
rect 330018 9092 330024 9104
rect 243228 9064 330024 9092
rect 243228 9052 243234 9064
rect 330018 9052 330024 9064
rect 330076 9052 330082 9104
rect 18322 8984 18328 9036
rect 18380 9024 18386 9036
rect 236178 9024 236184 9036
rect 18380 8996 236184 9024
rect 18380 8984 18386 8996
rect 236178 8984 236184 8996
rect 236236 8984 236242 9036
rect 239582 8984 239588 9036
rect 239640 9024 239646 9036
rect 328638 9024 328644 9036
rect 239640 8996 328644 9024
rect 239640 8984 239646 8996
rect 328638 8984 328644 8996
rect 328696 8984 328702 9036
rect 13630 8916 13636 8968
rect 13688 8956 13694 8968
rect 234798 8956 234804 8968
rect 13688 8928 234804 8956
rect 13688 8916 13694 8928
rect 234798 8916 234804 8928
rect 234856 8916 234862 8968
rect 235994 8916 236000 8968
rect 236052 8956 236058 8968
rect 325878 8956 325884 8968
rect 236052 8928 325884 8956
rect 236052 8916 236058 8928
rect 325878 8916 325884 8928
rect 325936 8916 325942 8968
rect 207474 8848 207480 8900
rect 207532 8888 207538 8900
rect 314930 8888 314936 8900
rect 207532 8860 314936 8888
rect 207532 8848 207538 8860
rect 314930 8848 314936 8860
rect 314988 8848 314994 8900
rect 210970 8780 210976 8832
rect 211028 8820 211034 8832
rect 316126 8820 316132 8832
rect 211028 8792 316132 8820
rect 211028 8780 211034 8792
rect 316126 8780 316132 8792
rect 316184 8780 316190 8832
rect 214650 8712 214656 8764
rect 214708 8752 214714 8764
rect 317506 8752 317512 8764
rect 214708 8724 317512 8752
rect 214708 8712 214714 8724
rect 317506 8712 317512 8724
rect 317564 8712 317570 8764
rect 218146 8644 218152 8696
rect 218204 8684 218210 8696
rect 318886 8684 318892 8696
rect 218204 8656 318892 8684
rect 218204 8644 218210 8656
rect 318886 8644 318892 8656
rect 318944 8644 318950 8696
rect 221734 8576 221740 8628
rect 221792 8616 221798 8628
rect 320174 8616 320180 8628
rect 221792 8588 320180 8616
rect 221792 8576 221798 8588
rect 320174 8576 320180 8588
rect 320232 8576 320238 8628
rect 225322 8508 225328 8560
rect 225380 8548 225386 8560
rect 321646 8548 321652 8560
rect 225380 8520 321652 8548
rect 225380 8508 225386 8520
rect 321646 8508 321652 8520
rect 321704 8508 321710 8560
rect 228910 8440 228916 8492
rect 228968 8480 228974 8492
rect 323118 8480 323124 8492
rect 228968 8452 323124 8480
rect 228968 8440 228974 8452
rect 323118 8440 323124 8452
rect 323176 8440 323182 8492
rect 232498 8372 232504 8424
rect 232556 8412 232562 8424
rect 324498 8412 324504 8424
rect 232556 8384 324504 8412
rect 232556 8372 232562 8384
rect 324498 8372 324504 8384
rect 324556 8372 324562 8424
rect 244366 8344 244372 8356
rect 244327 8316 244372 8344
rect 244366 8304 244372 8316
rect 244424 8304 244430 8356
rect 246758 8304 246764 8356
rect 246816 8344 246822 8356
rect 331398 8344 331404 8356
rect 246816 8316 331404 8344
rect 246816 8304 246822 8316
rect 331398 8304 331404 8316
rect 331456 8304 331462 8356
rect 389361 8347 389419 8353
rect 389361 8313 389373 8347
rect 389407 8344 389419 8347
rect 389450 8344 389456 8356
rect 389407 8316 389456 8344
rect 389407 8313 389419 8316
rect 389361 8307 389419 8313
rect 389450 8304 389456 8316
rect 389508 8304 389514 8356
rect 468754 8304 468760 8356
rect 468812 8344 468818 8356
rect 469030 8344 469036 8356
rect 468812 8316 469036 8344
rect 468812 8304 468818 8316
rect 469030 8304 469036 8316
rect 469088 8304 469094 8356
rect 87322 8236 87328 8288
rect 87380 8276 87386 8288
rect 265158 8276 265164 8288
rect 87380 8248 265164 8276
rect 87380 8236 87386 8248
rect 265158 8236 265164 8248
rect 265216 8236 265222 8288
rect 270494 8236 270500 8288
rect 270552 8276 270558 8288
rect 340966 8276 340972 8288
rect 270552 8248 340972 8276
rect 270552 8236 270558 8248
rect 340966 8236 340972 8248
rect 341024 8236 341030 8288
rect 445478 8236 445484 8288
rect 445536 8276 445542 8288
rect 523862 8276 523868 8288
rect 445536 8248 523868 8276
rect 445536 8236 445542 8248
rect 523862 8236 523868 8248
rect 523920 8236 523926 8288
rect 83826 8168 83832 8220
rect 83884 8208 83890 8220
rect 263870 8208 263876 8220
rect 83884 8180 263876 8208
rect 83884 8168 83890 8180
rect 263870 8168 263876 8180
rect 263928 8168 263934 8220
rect 266998 8168 267004 8220
rect 267056 8208 267062 8220
rect 339586 8208 339592 8220
rect 267056 8180 339592 8208
rect 267056 8168 267062 8180
rect 339586 8168 339592 8180
rect 339644 8168 339650 8220
rect 446950 8168 446956 8220
rect 447008 8208 447014 8220
rect 527450 8208 527456 8220
rect 447008 8180 527456 8208
rect 447008 8168 447014 8180
rect 527450 8168 527456 8180
rect 527508 8168 527514 8220
rect 2774 8100 2780 8152
rect 2832 8140 2838 8152
rect 4798 8140 4804 8152
rect 2832 8112 4804 8140
rect 2832 8100 2838 8112
rect 4798 8100 4804 8112
rect 4856 8100 4862 8152
rect 80238 8100 80244 8152
rect 80296 8140 80302 8152
rect 262398 8140 262404 8152
rect 80296 8112 262404 8140
rect 80296 8100 80302 8112
rect 262398 8100 262404 8112
rect 262456 8100 262462 8152
rect 263410 8100 263416 8152
rect 263468 8140 263474 8152
rect 338298 8140 338304 8152
rect 263468 8112 338304 8140
rect 263468 8100 263474 8112
rect 338298 8100 338304 8112
rect 338356 8100 338362 8152
rect 448238 8100 448244 8152
rect 448296 8140 448302 8152
rect 531038 8140 531044 8152
rect 448296 8112 531044 8140
rect 448296 8100 448302 8112
rect 531038 8100 531044 8112
rect 531096 8100 531102 8152
rect 40954 8032 40960 8084
rect 41012 8072 41018 8084
rect 245838 8072 245844 8084
rect 41012 8044 245844 8072
rect 41012 8032 41018 8044
rect 245838 8032 245844 8044
rect 245896 8032 245902 8084
rect 259822 8032 259828 8084
rect 259880 8072 259886 8084
rect 336918 8072 336924 8084
rect 259880 8044 336924 8072
rect 259880 8032 259886 8044
rect 336918 8032 336924 8044
rect 336976 8032 336982 8084
rect 450998 8032 451004 8084
rect 451056 8072 451062 8084
rect 534534 8072 534540 8084
rect 451056 8044 534540 8072
rect 451056 8032 451062 8044
rect 534534 8032 534540 8044
rect 534592 8032 534598 8084
rect 37366 7964 37372 8016
rect 37424 8004 37430 8016
rect 244366 8004 244372 8016
rect 37424 7976 244372 8004
rect 37424 7964 37430 7976
rect 244366 7964 244372 7976
rect 244424 7964 244430 8016
rect 256234 7964 256240 8016
rect 256292 8004 256298 8016
rect 334066 8004 334072 8016
rect 256292 7976 334072 8004
rect 256292 7964 256298 7976
rect 334066 7964 334072 7976
rect 334124 7964 334130 8016
rect 452470 7964 452476 8016
rect 452528 8004 452534 8016
rect 538122 8004 538128 8016
rect 452528 7976 538128 8004
rect 452528 7964 452534 7976
rect 538122 7964 538128 7976
rect 538180 7964 538186 8016
rect 33870 7896 33876 7948
rect 33928 7936 33934 7948
rect 242986 7936 242992 7948
rect 33928 7908 242992 7936
rect 33928 7896 33934 7908
rect 242986 7896 242992 7908
rect 243044 7896 243050 7948
rect 252646 7896 252652 7948
rect 252704 7936 252710 7948
rect 332686 7936 332692 7948
rect 252704 7908 332692 7936
rect 252704 7896 252710 7908
rect 332686 7896 332692 7908
rect 332744 7896 332750 7948
rect 453758 7896 453764 7948
rect 453816 7936 453822 7948
rect 541710 7936 541716 7948
rect 453816 7908 541716 7936
rect 453816 7896 453822 7908
rect 541710 7896 541716 7908
rect 541768 7896 541774 7948
rect 30282 7828 30288 7880
rect 30340 7868 30346 7880
rect 241790 7868 241796 7880
rect 30340 7840 241796 7868
rect 30340 7828 30346 7840
rect 241790 7828 241796 7840
rect 241848 7828 241854 7880
rect 249150 7828 249156 7880
rect 249208 7868 249214 7880
rect 331306 7868 331312 7880
rect 249208 7840 331312 7868
rect 249208 7828 249214 7840
rect 331306 7828 331312 7840
rect 331364 7828 331370 7880
rect 455230 7828 455236 7880
rect 455288 7868 455294 7880
rect 545298 7868 545304 7880
rect 455288 7840 545304 7868
rect 455288 7828 455294 7840
rect 545298 7828 545304 7840
rect 545356 7828 545362 7880
rect 26694 7760 26700 7812
rect 26752 7800 26758 7812
rect 240410 7800 240416 7812
rect 26752 7772 240416 7800
rect 26752 7760 26758 7772
rect 240410 7760 240416 7772
rect 240468 7760 240474 7812
rect 245562 7760 245568 7812
rect 245620 7800 245626 7812
rect 330110 7800 330116 7812
rect 245620 7772 330116 7800
rect 245620 7760 245626 7772
rect 330110 7760 330116 7772
rect 330168 7760 330174 7812
rect 456610 7760 456616 7812
rect 456668 7800 456674 7812
rect 548886 7800 548892 7812
rect 456668 7772 548892 7800
rect 456668 7760 456674 7772
rect 548886 7760 548892 7772
rect 548944 7760 548950 7812
rect 21910 7692 21916 7744
rect 21968 7732 21974 7744
rect 238846 7732 238852 7744
rect 21968 7704 238852 7732
rect 21968 7692 21974 7704
rect 238846 7692 238852 7704
rect 238904 7692 238910 7744
rect 241974 7692 241980 7744
rect 242032 7732 242038 7744
rect 328546 7732 328552 7744
rect 242032 7704 328552 7732
rect 242032 7692 242038 7704
rect 328546 7692 328552 7704
rect 328604 7692 328610 7744
rect 457990 7692 457996 7744
rect 458048 7732 458054 7744
rect 552382 7732 552388 7744
rect 458048 7704 552388 7732
rect 458048 7692 458054 7704
rect 552382 7692 552388 7704
rect 552440 7692 552446 7744
rect 8846 7624 8852 7676
rect 8904 7664 8910 7676
rect 227533 7667 227591 7673
rect 227533 7664 227545 7667
rect 8904 7636 227545 7664
rect 8904 7624 8910 7636
rect 227533 7633 227545 7636
rect 227579 7633 227591 7667
rect 230658 7664 230664 7676
rect 227533 7627 227591 7633
rect 227640 7636 230664 7664
rect 4062 7556 4068 7608
rect 4120 7596 4126 7608
rect 227640 7596 227668 7636
rect 230658 7624 230664 7636
rect 230716 7624 230722 7676
rect 234798 7624 234804 7676
rect 234856 7664 234862 7676
rect 325786 7664 325792 7676
rect 234856 7636 325792 7664
rect 234856 7624 234862 7636
rect 325786 7624 325792 7636
rect 325844 7624 325850 7676
rect 459370 7624 459376 7676
rect 459428 7664 459434 7676
rect 555970 7664 555976 7676
rect 459428 7636 555976 7664
rect 459428 7624 459434 7636
rect 555970 7624 555976 7636
rect 556028 7624 556034 7676
rect 4120 7568 227668 7596
rect 4120 7556 4126 7568
rect 227714 7556 227720 7608
rect 227772 7596 227778 7608
rect 229002 7596 229008 7608
rect 227772 7568 229008 7596
rect 227772 7556 227778 7568
rect 229002 7556 229008 7568
rect 229060 7556 229066 7608
rect 231302 7556 231308 7608
rect 231360 7596 231366 7608
rect 324406 7596 324412 7608
rect 231360 7568 324412 7596
rect 231360 7556 231366 7568
rect 324406 7556 324412 7568
rect 324464 7556 324470 7608
rect 460750 7556 460756 7608
rect 460808 7596 460814 7608
rect 559558 7596 559564 7608
rect 460808 7568 559564 7596
rect 460808 7556 460814 7568
rect 559558 7556 559564 7568
rect 559616 7556 559622 7608
rect 134886 7488 134892 7540
rect 134944 7528 134950 7540
rect 284570 7528 284576 7540
rect 134944 7500 284576 7528
rect 134944 7488 134950 7500
rect 284570 7488 284576 7500
rect 284628 7488 284634 7540
rect 444190 7488 444196 7540
rect 444248 7528 444254 7540
rect 520274 7528 520280 7540
rect 444248 7500 520280 7528
rect 444248 7488 444254 7500
rect 520274 7488 520280 7500
rect 520332 7488 520338 7540
rect 138474 7420 138480 7472
rect 138532 7460 138538 7472
rect 285950 7460 285956 7472
rect 138532 7432 285956 7460
rect 138532 7420 138538 7432
rect 285950 7420 285956 7432
rect 286008 7420 286014 7472
rect 442810 7420 442816 7472
rect 442868 7460 442874 7472
rect 516778 7460 516784 7472
rect 442868 7432 516784 7460
rect 442868 7420 442874 7432
rect 516778 7420 516784 7432
rect 516836 7420 516842 7472
rect 141970 7352 141976 7404
rect 142028 7392 142034 7404
rect 287054 7392 287060 7404
rect 142028 7364 287060 7392
rect 142028 7352 142034 7364
rect 287054 7352 287060 7364
rect 287112 7352 287118 7404
rect 441430 7352 441436 7404
rect 441488 7392 441494 7404
rect 513190 7392 513196 7404
rect 441488 7364 513196 7392
rect 441488 7352 441494 7364
rect 513190 7352 513196 7364
rect 513248 7352 513254 7404
rect 145650 7284 145656 7336
rect 145708 7324 145714 7336
rect 288434 7324 288440 7336
rect 145708 7296 288440 7324
rect 145708 7284 145714 7296
rect 288434 7284 288440 7296
rect 288492 7284 288498 7336
rect 440050 7284 440056 7336
rect 440108 7324 440114 7336
rect 509602 7324 509608 7336
rect 440108 7296 509608 7324
rect 440108 7284 440114 7296
rect 509602 7284 509608 7296
rect 509660 7284 509666 7336
rect 149238 7216 149244 7268
rect 149296 7256 149302 7268
rect 291194 7256 291200 7268
rect 149296 7228 291200 7256
rect 149296 7216 149302 7228
rect 291194 7216 291200 7228
rect 291252 7216 291258 7268
rect 152734 7148 152740 7200
rect 152792 7188 152798 7200
rect 292574 7188 292580 7200
rect 152792 7160 292580 7188
rect 152792 7148 152798 7160
rect 292574 7148 292580 7160
rect 292632 7148 292638 7200
rect 156322 7080 156328 7132
rect 156380 7120 156386 7132
rect 293954 7120 293960 7132
rect 156380 7092 293960 7120
rect 156380 7080 156386 7092
rect 293954 7080 293960 7092
rect 294012 7080 294018 7132
rect 159910 7012 159916 7064
rect 159968 7052 159974 7064
rect 295334 7052 295340 7064
rect 159968 7024 295340 7052
rect 159968 7012 159974 7024
rect 295334 7012 295340 7024
rect 295392 7012 295398 7064
rect 227533 6987 227591 6993
rect 227533 6953 227545 6987
rect 227579 6984 227591 6987
rect 233418 6984 233424 6996
rect 227579 6956 233424 6984
rect 227579 6953 227591 6956
rect 227533 6947 227591 6953
rect 233418 6944 233424 6956
rect 233476 6944 233482 6996
rect 238386 6944 238392 6996
rect 238444 6984 238450 6996
rect 327166 6984 327172 6996
rect 238444 6956 327172 6984
rect 238444 6944 238450 6956
rect 327166 6944 327172 6956
rect 327224 6944 327230 6996
rect 516686 6876 516692 6928
rect 516744 6916 516750 6928
rect 516870 6916 516876 6928
rect 516744 6888 516876 6916
rect 516744 6876 516750 6888
rect 516870 6876 516876 6888
rect 516928 6876 516934 6928
rect 170582 6808 170588 6860
rect 170640 6848 170646 6860
rect 299474 6848 299480 6860
rect 170640 6820 299480 6848
rect 170640 6808 170646 6820
rect 299474 6808 299480 6820
rect 299532 6808 299538 6860
rect 431770 6808 431776 6860
rect 431828 6848 431834 6860
rect 490558 6848 490564 6860
rect 431828 6820 490564 6848
rect 431828 6808 431834 6820
rect 490558 6808 490564 6820
rect 490616 6808 490622 6860
rect 167086 6740 167092 6792
rect 167144 6780 167150 6792
rect 298370 6780 298376 6792
rect 167144 6752 298376 6780
rect 167144 6740 167150 6752
rect 298370 6740 298376 6752
rect 298428 6740 298434 6792
rect 433150 6740 433156 6792
rect 433208 6780 433214 6792
rect 491754 6780 491760 6792
rect 433208 6752 491760 6780
rect 433208 6740 433214 6752
rect 491754 6740 491760 6752
rect 491812 6740 491818 6792
rect 163498 6672 163504 6724
rect 163556 6712 163562 6724
rect 296714 6712 296720 6724
rect 163556 6684 296720 6712
rect 163556 6672 163562 6684
rect 296714 6672 296720 6684
rect 296772 6672 296778 6724
rect 297358 6672 297364 6724
rect 297416 6712 297422 6724
rect 336826 6712 336832 6724
rect 297416 6684 336832 6712
rect 297416 6672 297422 6684
rect 336826 6672 336832 6684
rect 336884 6672 336890 6724
rect 434622 6672 434628 6724
rect 434680 6712 434686 6724
rect 495342 6712 495348 6724
rect 434680 6684 495348 6712
rect 434680 6672 434686 6684
rect 495342 6672 495348 6684
rect 495400 6672 495406 6724
rect 131390 6604 131396 6656
rect 131448 6644 131454 6656
rect 283006 6644 283012 6656
rect 131448 6616 283012 6644
rect 131448 6604 131454 6616
rect 283006 6604 283012 6616
rect 283064 6604 283070 6656
rect 295886 6604 295892 6656
rect 295944 6644 295950 6656
rect 335446 6644 335452 6656
rect 295944 6616 335452 6644
rect 295944 6604 295950 6616
rect 335446 6604 335452 6616
rect 335504 6604 335510 6656
rect 433242 6604 433248 6656
rect 433300 6644 433306 6656
rect 494146 6644 494152 6656
rect 433300 6616 494152 6644
rect 433300 6604 433306 6616
rect 494146 6604 494152 6616
rect 494204 6604 494210 6656
rect 76650 6536 76656 6588
rect 76708 6576 76714 6588
rect 261018 6576 261024 6588
rect 76708 6548 261024 6576
rect 76708 6536 76714 6548
rect 261018 6536 261024 6548
rect 261076 6536 261082 6588
rect 298094 6536 298100 6588
rect 298152 6576 298158 6588
rect 338390 6576 338396 6588
rect 298152 6548 338396 6576
rect 298152 6536 298158 6548
rect 338390 6536 338396 6548
rect 338448 6536 338454 6588
rect 435910 6536 435916 6588
rect 435968 6576 435974 6588
rect 497734 6576 497740 6588
rect 435968 6548 497740 6576
rect 435968 6536 435974 6548
rect 497734 6536 497740 6548
rect 497792 6536 497798 6588
rect 73062 6468 73068 6520
rect 73120 6508 73126 6520
rect 259454 6508 259460 6520
rect 73120 6480 259460 6508
rect 73120 6468 73126 6480
rect 259454 6468 259460 6480
rect 259512 6468 259518 6520
rect 289814 6468 289820 6520
rect 289872 6508 289878 6520
rect 339678 6508 339684 6520
rect 289872 6480 339684 6508
rect 289872 6468 289878 6480
rect 339678 6468 339684 6480
rect 339736 6468 339742 6520
rect 436002 6468 436008 6520
rect 436060 6508 436066 6520
rect 498930 6508 498936 6520
rect 436060 6480 498936 6508
rect 436060 6468 436066 6480
rect 498930 6468 498936 6480
rect 498988 6468 498994 6520
rect 69474 6400 69480 6452
rect 69532 6440 69538 6452
rect 258258 6440 258264 6452
rect 69532 6412 258264 6440
rect 69532 6400 69538 6412
rect 258258 6400 258264 6412
rect 258316 6400 258322 6452
rect 288434 6400 288440 6452
rect 288492 6440 288498 6452
rect 341242 6440 341248 6452
rect 288492 6412 341248 6440
rect 288492 6400 288498 6412
rect 341242 6400 341248 6412
rect 341300 6400 341306 6452
rect 437382 6400 437388 6452
rect 437440 6440 437446 6452
rect 501230 6440 501236 6452
rect 437440 6412 501236 6440
rect 437440 6400 437446 6412
rect 501230 6400 501236 6412
rect 501288 6400 501294 6452
rect 65978 6332 65984 6384
rect 66036 6372 66042 6384
rect 256786 6372 256792 6384
rect 66036 6344 256792 6372
rect 66036 6332 66042 6344
rect 256786 6332 256792 6344
rect 256844 6332 256850 6384
rect 288526 6332 288532 6384
rect 288584 6372 288590 6384
rect 343634 6372 343640 6384
rect 288584 6344 343640 6372
rect 288584 6332 288590 6344
rect 343634 6332 343640 6344
rect 343692 6332 343698 6384
rect 438670 6332 438676 6384
rect 438728 6372 438734 6384
rect 504818 6372 504824 6384
rect 438728 6344 504824 6372
rect 438728 6332 438734 6344
rect 504818 6332 504824 6344
rect 504876 6332 504882 6384
rect 62390 6264 62396 6316
rect 62448 6304 62454 6316
rect 255498 6304 255504 6316
rect 62448 6276 255504 6304
rect 62448 6264 62454 6276
rect 255498 6264 255504 6276
rect 255556 6264 255562 6316
rect 294322 6264 294328 6316
rect 294380 6304 294386 6316
rect 350626 6304 350632 6316
rect 294380 6276 350632 6304
rect 294380 6264 294386 6276
rect 350626 6264 350632 6276
rect 350684 6264 350690 6316
rect 437290 6264 437296 6316
rect 437348 6304 437354 6316
rect 502426 6304 502432 6316
rect 437348 6276 502432 6304
rect 437348 6264 437354 6276
rect 502426 6264 502432 6276
rect 502484 6264 502490 6316
rect 58802 6196 58808 6248
rect 58860 6236 58866 6248
rect 253934 6236 253940 6248
rect 58860 6208 253940 6236
rect 58860 6196 58866 6208
rect 253934 6196 253940 6208
rect 253992 6196 253998 6248
rect 280062 6196 280068 6248
rect 280120 6236 280126 6248
rect 345198 6236 345204 6248
rect 280120 6208 345204 6236
rect 280120 6196 280126 6208
rect 345198 6196 345204 6208
rect 345256 6196 345262 6248
rect 438762 6196 438768 6248
rect 438820 6236 438826 6248
rect 506014 6236 506020 6248
rect 438820 6208 506020 6236
rect 438820 6196 438826 6208
rect 506014 6196 506020 6208
rect 506072 6196 506078 6248
rect 55214 6128 55220 6180
rect 55272 6168 55278 6180
rect 251358 6168 251364 6180
rect 55272 6140 251364 6168
rect 55272 6128 55278 6140
rect 251358 6128 251364 6140
rect 251416 6128 251422 6180
rect 274082 6128 274088 6180
rect 274140 6168 274146 6180
rect 342346 6168 342352 6180
rect 274140 6140 342352 6168
rect 274140 6128 274146 6140
rect 342346 6128 342352 6140
rect 342404 6128 342410 6180
rect 440142 6128 440148 6180
rect 440200 6168 440206 6180
rect 508406 6168 508412 6180
rect 440200 6140 508412 6168
rect 440200 6128 440206 6140
rect 508406 6128 508412 6140
rect 508464 6128 508470 6180
rect 174170 6060 174176 6112
rect 174228 6100 174234 6112
rect 300854 6100 300860 6112
rect 174228 6072 300860 6100
rect 174228 6060 174234 6072
rect 300854 6060 300860 6072
rect 300912 6060 300918 6112
rect 430390 6060 430396 6112
rect 430448 6100 430454 6112
rect 486970 6100 486976 6112
rect 430448 6072 486976 6100
rect 430448 6060 430454 6072
rect 486970 6060 486976 6072
rect 487028 6060 487034 6112
rect 177758 5992 177764 6044
rect 177816 6032 177822 6044
rect 302234 6032 302240 6044
rect 177816 6004 302240 6032
rect 177816 5992 177822 6004
rect 302234 5992 302240 6004
rect 302292 5992 302298 6044
rect 431862 5992 431868 6044
rect 431920 6032 431926 6044
rect 488166 6032 488172 6044
rect 431920 6004 488172 6032
rect 431920 5992 431926 6004
rect 488166 5992 488172 6004
rect 488224 5992 488230 6044
rect 181346 5924 181352 5976
rect 181404 5964 181410 5976
rect 303614 5964 303620 5976
rect 181404 5936 303620 5964
rect 181404 5924 181410 5936
rect 303614 5924 303620 5936
rect 303672 5924 303678 5976
rect 430482 5924 430488 5976
rect 430540 5964 430546 5976
rect 484578 5964 484584 5976
rect 430540 5936 484584 5964
rect 430540 5924 430546 5936
rect 484578 5924 484584 5936
rect 484636 5924 484642 5976
rect 184842 5856 184848 5908
rect 184900 5896 184906 5908
rect 304994 5896 305000 5908
rect 184900 5868 305000 5896
rect 184900 5856 184906 5868
rect 304994 5856 305000 5868
rect 305052 5856 305058 5908
rect 429102 5856 429108 5908
rect 429160 5896 429166 5908
rect 483474 5896 483480 5908
rect 429160 5868 483480 5896
rect 429160 5856 429166 5868
rect 483474 5856 483480 5868
rect 483532 5856 483538 5908
rect 188430 5788 188436 5840
rect 188488 5828 188494 5840
rect 306650 5828 306656 5840
rect 188488 5800 306656 5828
rect 188488 5788 188494 5800
rect 306650 5788 306656 5800
rect 306708 5788 306714 5840
rect 427722 5788 427728 5840
rect 427780 5828 427786 5840
rect 479886 5828 479892 5840
rect 427780 5800 479892 5828
rect 427780 5788 427786 5800
rect 479886 5788 479892 5800
rect 479944 5788 479950 5840
rect 192018 5720 192024 5772
rect 192076 5760 192082 5772
rect 307754 5760 307760 5772
rect 192076 5732 307760 5760
rect 192076 5720 192082 5732
rect 307754 5720 307760 5732
rect 307812 5720 307818 5772
rect 426342 5720 426348 5772
rect 426400 5760 426406 5772
rect 476298 5760 476304 5772
rect 426400 5732 476304 5760
rect 426400 5720 426406 5732
rect 476298 5720 476304 5732
rect 476356 5720 476362 5772
rect 195606 5652 195612 5704
rect 195664 5692 195670 5704
rect 309134 5692 309140 5704
rect 195664 5664 309140 5692
rect 195664 5652 195670 5664
rect 309134 5652 309140 5664
rect 309192 5652 309198 5704
rect 199194 5584 199200 5636
rect 199252 5624 199258 5636
rect 310514 5624 310520 5636
rect 199252 5596 310520 5624
rect 199252 5584 199258 5596
rect 310514 5584 310520 5596
rect 310572 5584 310578 5636
rect 470594 5584 470600 5636
rect 470652 5624 470658 5636
rect 471517 5627 471575 5633
rect 471517 5624 471529 5627
rect 470652 5596 471529 5624
rect 470652 5584 470658 5596
rect 471517 5593 471529 5596
rect 471563 5593 471575 5627
rect 471517 5587 471575 5593
rect 202690 5516 202696 5568
rect 202748 5556 202754 5568
rect 313274 5556 313280 5568
rect 202748 5528 313280 5556
rect 202748 5516 202754 5528
rect 313274 5516 313280 5528
rect 313332 5516 313338 5568
rect 319533 5559 319591 5565
rect 319533 5525 319545 5559
rect 319579 5556 319591 5559
rect 327074 5556 327080 5568
rect 319579 5528 327080 5556
rect 319579 5525 319591 5528
rect 319533 5519 319591 5525
rect 327074 5516 327080 5528
rect 327132 5516 327138 5568
rect 468938 5516 468944 5568
rect 468996 5556 469002 5568
rect 471425 5559 471483 5565
rect 471425 5556 471437 5559
rect 468996 5528 471437 5556
rect 468996 5516 469002 5528
rect 471425 5525 471437 5528
rect 471471 5525 471483 5559
rect 471425 5519 471483 5525
rect 137278 5448 137284 5500
rect 137336 5488 137342 5500
rect 285674 5488 285680 5500
rect 137336 5460 285680 5488
rect 137336 5448 137342 5460
rect 285674 5448 285680 5460
rect 285732 5448 285738 5500
rect 287701 5491 287759 5497
rect 287701 5457 287713 5491
rect 287747 5488 287759 5491
rect 297085 5491 297143 5497
rect 297085 5488 297097 5491
rect 287747 5460 297097 5488
rect 287747 5457 287759 5460
rect 287701 5451 287759 5457
rect 297085 5457 297097 5460
rect 297131 5457 297143 5491
rect 297085 5451 297143 5457
rect 297818 5448 297824 5500
rect 297876 5488 297882 5500
rect 352098 5488 352104 5500
rect 297876 5460 352104 5488
rect 297876 5448 297882 5460
rect 352098 5448 352104 5460
rect 352156 5448 352162 5500
rect 452562 5448 452568 5500
rect 452620 5488 452626 5500
rect 540514 5488 540520 5500
rect 452620 5460 540520 5488
rect 452620 5448 452626 5460
rect 540514 5448 540520 5460
rect 540572 5448 540578 5500
rect 133782 5380 133788 5432
rect 133840 5420 133846 5432
rect 284294 5420 284300 5432
rect 133840 5392 284300 5420
rect 133840 5380 133846 5392
rect 284294 5380 284300 5392
rect 284352 5380 284358 5432
rect 290734 5380 290740 5432
rect 290792 5420 290798 5432
rect 349338 5420 349344 5432
rect 290792 5392 349344 5420
rect 290792 5380 290798 5392
rect 349338 5380 349344 5392
rect 349396 5380 349402 5432
rect 408402 5380 408408 5432
rect 408460 5420 408466 5432
rect 433518 5420 433524 5432
rect 408460 5392 433524 5420
rect 408460 5380 408466 5392
rect 433518 5380 433524 5392
rect 433576 5380 433582 5432
rect 453850 5380 453856 5432
rect 453908 5420 453914 5432
rect 544102 5420 544108 5432
rect 453908 5392 544108 5420
rect 453908 5380 453914 5392
rect 544102 5380 544108 5392
rect 544160 5380 544166 5432
rect 130194 5312 130200 5364
rect 130252 5352 130258 5364
rect 283190 5352 283196 5364
rect 130252 5324 283196 5352
rect 130252 5312 130258 5324
rect 283190 5312 283196 5324
rect 283248 5312 283254 5364
rect 287146 5312 287152 5364
rect 287204 5352 287210 5364
rect 347958 5352 347964 5364
rect 287204 5324 347964 5352
rect 287204 5312 287210 5324
rect 347958 5312 347964 5324
rect 348016 5312 348022 5364
rect 412358 5312 412364 5364
rect 412416 5352 412422 5364
rect 440602 5352 440608 5364
rect 412416 5324 440608 5352
rect 412416 5312 412422 5324
rect 440602 5312 440608 5324
rect 440660 5312 440666 5364
rect 455322 5312 455328 5364
rect 455380 5352 455386 5364
rect 547690 5352 547696 5364
rect 455380 5324 547696 5352
rect 455380 5312 455386 5324
rect 547690 5312 547696 5324
rect 547748 5312 547754 5364
rect 67174 5244 67180 5296
rect 67232 5284 67238 5296
rect 256970 5284 256976 5296
rect 67232 5256 256976 5284
rect 67232 5244 67238 5256
rect 256970 5244 256976 5256
rect 257028 5244 257034 5296
rect 268381 5287 268439 5293
rect 268381 5253 268393 5287
rect 268427 5284 268439 5287
rect 278041 5287 278099 5293
rect 278041 5284 278053 5287
rect 268427 5256 278053 5284
rect 268427 5253 268439 5256
rect 268381 5247 268439 5253
rect 278041 5253 278053 5256
rect 278087 5253 278099 5287
rect 278041 5247 278099 5253
rect 283650 5244 283656 5296
rect 283708 5284 283714 5296
rect 346578 5284 346584 5296
rect 283708 5256 346584 5284
rect 283708 5244 283714 5256
rect 346578 5244 346584 5256
rect 346636 5244 346642 5296
rect 413830 5244 413836 5296
rect 413888 5284 413894 5296
rect 444190 5284 444196 5296
rect 413888 5256 444196 5284
rect 413888 5244 413894 5256
rect 444190 5244 444196 5256
rect 444248 5244 444254 5296
rect 459462 5244 459468 5296
rect 459520 5284 459526 5296
rect 466089 5287 466147 5293
rect 459520 5256 466040 5284
rect 459520 5244 459526 5256
rect 48130 5176 48136 5228
rect 48188 5216 48194 5228
rect 248506 5216 248512 5228
rect 48188 5188 248512 5216
rect 48188 5176 48194 5188
rect 248506 5176 248512 5188
rect 248564 5176 248570 5228
rect 251450 5176 251456 5228
rect 251508 5216 251514 5228
rect 332594 5216 332600 5228
rect 251508 5188 332600 5216
rect 251508 5176 251514 5188
rect 332594 5176 332600 5188
rect 332652 5176 332658 5228
rect 415302 5176 415308 5228
rect 415360 5216 415366 5228
rect 447778 5216 447784 5228
rect 415360 5188 447784 5216
rect 415360 5176 415366 5188
rect 447778 5176 447784 5188
rect 447836 5176 447842 5228
rect 460842 5176 460848 5228
rect 460900 5216 460906 5228
rect 466012 5216 466040 5256
rect 466089 5253 466101 5287
rect 466135 5284 466147 5287
rect 551186 5284 551192 5296
rect 466135 5256 551192 5284
rect 466135 5253 466147 5256
rect 466089 5247 466147 5253
rect 551186 5244 551192 5256
rect 551244 5244 551250 5296
rect 554774 5216 554780 5228
rect 460900 5188 465948 5216
rect 466012 5188 554780 5216
rect 460900 5176 460906 5188
rect 17218 5108 17224 5160
rect 17276 5148 17282 5160
rect 236086 5148 236092 5160
rect 17276 5120 236092 5148
rect 17276 5108 17282 5120
rect 236086 5108 236092 5120
rect 236144 5108 236150 5160
rect 247954 5108 247960 5160
rect 248012 5148 248018 5160
rect 331214 5148 331220 5160
rect 248012 5120 331220 5148
rect 248012 5108 248018 5120
rect 331214 5108 331220 5120
rect 331272 5108 331278 5160
rect 416498 5108 416504 5160
rect 416556 5148 416562 5160
rect 451274 5148 451280 5160
rect 416556 5120 451280 5148
rect 416556 5108 416562 5120
rect 451274 5108 451280 5120
rect 451332 5108 451338 5160
rect 461213 5151 461271 5157
rect 461213 5117 461225 5151
rect 461259 5148 461271 5151
rect 461259 5120 462268 5148
rect 461259 5117 461271 5120
rect 461213 5111 461271 5117
rect 12434 5040 12440 5092
rect 12492 5080 12498 5092
rect 234706 5080 234712 5092
rect 12492 5052 234712 5080
rect 12492 5040 12498 5052
rect 234706 5040 234712 5052
rect 234764 5040 234770 5092
rect 244366 5040 244372 5092
rect 244424 5080 244430 5092
rect 324133 5083 324191 5089
rect 324133 5080 324145 5083
rect 244424 5052 324145 5080
rect 244424 5040 244430 5052
rect 324133 5049 324145 5052
rect 324179 5049 324191 5083
rect 324133 5043 324191 5049
rect 327169 5083 327227 5089
rect 327169 5049 327181 5083
rect 327215 5080 327227 5083
rect 329834 5080 329840 5092
rect 327215 5052 329840 5080
rect 327215 5049 327227 5052
rect 327169 5043 327227 5049
rect 329834 5040 329840 5052
rect 329892 5040 329898 5092
rect 337102 5040 337108 5092
rect 337160 5080 337166 5092
rect 368566 5080 368572 5092
rect 337160 5052 368572 5080
rect 337160 5040 337166 5052
rect 368566 5040 368572 5052
rect 368624 5040 368630 5092
rect 417970 5040 417976 5092
rect 418028 5080 418034 5092
rect 454862 5080 454868 5092
rect 418028 5052 454868 5080
rect 418028 5040 418034 5052
rect 454862 5040 454868 5052
rect 454920 5040 454926 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 232130 5012 232136 5024
rect 7708 4984 232136 5012
rect 7708 4972 7714 4984
rect 232130 4972 232136 4984
rect 232188 4972 232194 5024
rect 240778 4972 240784 5024
rect 240836 5012 240842 5024
rect 249061 5015 249119 5021
rect 249061 5012 249073 5015
rect 240836 4984 249073 5012
rect 240836 4972 240842 4984
rect 249061 4981 249073 4984
rect 249107 4981 249119 5015
rect 249061 4975 249119 4981
rect 258721 5015 258779 5021
rect 258721 4981 258733 5015
rect 258767 5012 258779 5015
rect 268381 5015 268439 5021
rect 268381 5012 268393 5015
rect 258767 4984 268393 5012
rect 258767 4981 258779 4984
rect 258721 4975 258779 4981
rect 268381 4981 268393 4984
rect 268427 4981 268439 5015
rect 268381 4975 268439 4981
rect 278041 5015 278099 5021
rect 278041 4981 278053 5015
rect 278087 5012 278099 5015
rect 287701 5015 287759 5021
rect 287701 5012 287713 5015
rect 278087 4984 287713 5012
rect 278087 4981 278099 4984
rect 278041 4975 278099 4981
rect 287701 4981 287713 4984
rect 287747 4981 287759 5015
rect 287701 4975 287759 4981
rect 297085 5015 297143 5021
rect 297085 4981 297097 5015
rect 297131 5012 297143 5015
rect 307021 5015 307079 5021
rect 307021 5012 307033 5015
rect 297131 4984 307033 5012
rect 297131 4981 297143 4984
rect 297085 4975 297143 4981
rect 307021 4981 307033 4984
rect 307067 4981 307079 5015
rect 307021 4975 307079 4981
rect 315942 4972 315948 5024
rect 316000 5012 316006 5024
rect 325145 5015 325203 5021
rect 325145 5012 325157 5015
rect 316000 4984 325157 5012
rect 316000 4972 316006 4984
rect 325145 4981 325157 4984
rect 325191 4981 325203 5015
rect 325145 4975 325203 4981
rect 325602 4972 325608 5024
rect 325660 5012 325666 5024
rect 338114 5012 338120 5024
rect 325660 4984 338120 5012
rect 325660 4972 325666 4984
rect 338114 4972 338120 4984
rect 338172 4972 338178 5024
rect 419442 4972 419448 5024
rect 419500 5012 419506 5024
rect 458450 5012 458456 5024
rect 419500 4984 458456 5012
rect 419500 4972 419506 4984
rect 458450 4972 458456 4984
rect 458508 4972 458514 5024
rect 462240 5012 462268 5120
rect 463510 5108 463516 5160
rect 463568 5148 463574 5160
rect 465920 5148 465948 5188
rect 554774 5176 554780 5188
rect 554832 5176 554838 5228
rect 558362 5148 558368 5160
rect 463568 5120 465856 5148
rect 465920 5120 558368 5148
rect 463568 5108 463574 5120
rect 464982 5040 464988 5092
rect 465040 5080 465046 5092
rect 465828 5080 465856 5120
rect 558362 5108 558368 5120
rect 558420 5108 558426 5160
rect 471333 5083 471391 5089
rect 465040 5052 465764 5080
rect 465828 5052 471284 5080
rect 465040 5040 465046 5052
rect 465626 5012 465632 5024
rect 462240 4984 465632 5012
rect 465626 4972 465632 4984
rect 465684 4972 465690 5024
rect 465736 5012 465764 5052
rect 471256 5012 471284 5052
rect 471333 5049 471345 5083
rect 471379 5080 471391 5083
rect 561950 5080 561956 5092
rect 471379 5052 561956 5080
rect 471379 5049 471391 5052
rect 471333 5043 471391 5049
rect 561950 5040 561956 5052
rect 562008 5040 562014 5092
rect 565538 5012 565544 5024
rect 465736 4984 471192 5012
rect 471256 4984 565544 5012
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 230566 4944 230572 4956
rect 2924 4916 230572 4944
rect 2924 4904 2930 4916
rect 230566 4904 230572 4916
rect 230624 4904 230630 4956
rect 237190 4904 237196 4956
rect 237248 4944 237254 4956
rect 319533 4947 319591 4953
rect 319533 4944 319545 4947
rect 237248 4916 319545 4944
rect 237248 4904 237254 4916
rect 319533 4913 319545 4916
rect 319579 4913 319591 4947
rect 319533 4907 319591 4913
rect 320913 4947 320971 4953
rect 320913 4913 320925 4947
rect 320959 4944 320971 4947
rect 326341 4947 326399 4953
rect 326341 4944 326353 4947
rect 320959 4916 326353 4944
rect 320959 4913 320971 4916
rect 320913 4907 320971 4913
rect 326341 4913 326353 4916
rect 326387 4913 326399 4947
rect 328730 4944 328736 4956
rect 326341 4907 326399 4913
rect 326540 4916 328736 4944
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 230474 4876 230480 4888
rect 1728 4848 223160 4876
rect 1728 4836 1734 4848
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 220265 4811 220323 4817
rect 220265 4808 220277 4811
rect 624 4780 220277 4808
rect 624 4768 630 4780
rect 220265 4777 220277 4780
rect 220311 4777 220323 4811
rect 223132 4808 223160 4848
rect 227732 4848 230480 4876
rect 227732 4808 227760 4848
rect 230474 4836 230480 4848
rect 230532 4836 230538 4888
rect 233694 4836 233700 4888
rect 233752 4876 233758 4888
rect 320637 4879 320695 4885
rect 320637 4876 320649 4879
rect 233752 4848 320649 4876
rect 233752 4836 233758 4848
rect 320637 4845 320649 4848
rect 320683 4845 320695 4879
rect 320637 4839 320695 4845
rect 320821 4879 320879 4885
rect 320821 4845 320833 4879
rect 320867 4876 320879 4879
rect 325694 4876 325700 4888
rect 320867 4848 325700 4876
rect 320867 4845 320879 4848
rect 320821 4839 320879 4845
rect 325694 4836 325700 4848
rect 325752 4836 325758 4888
rect 223132 4780 227760 4808
rect 220265 4771 220323 4777
rect 230106 4768 230112 4820
rect 230164 4808 230170 4820
rect 325145 4811 325203 4817
rect 230164 4780 320220 4808
rect 230164 4768 230170 4780
rect 212258 4700 212264 4752
rect 212316 4740 212322 4752
rect 316034 4740 316040 4752
rect 212316 4712 316040 4740
rect 212316 4700 212322 4712
rect 316034 4700 316040 4712
rect 316092 4700 316098 4752
rect 318702 4700 318708 4752
rect 318760 4740 318766 4752
rect 320085 4743 320143 4749
rect 320085 4740 320097 4743
rect 318760 4712 320097 4740
rect 318760 4700 318766 4712
rect 320085 4709 320097 4712
rect 320131 4709 320143 4743
rect 320192 4740 320220 4780
rect 325145 4777 325157 4811
rect 325191 4808 325203 4811
rect 326540 4808 326568 4916
rect 328730 4904 328736 4916
rect 328788 4904 328794 4956
rect 333606 4904 333612 4956
rect 333664 4944 333670 4956
rect 367186 4944 367192 4956
rect 333664 4916 367192 4944
rect 333664 4904 333670 4916
rect 367186 4904 367192 4916
rect 367244 4904 367250 4956
rect 420730 4904 420736 4956
rect 420788 4944 420794 4956
rect 454681 4947 454739 4953
rect 454681 4944 454693 4947
rect 420788 4916 454693 4944
rect 420788 4904 420794 4916
rect 454681 4913 454693 4916
rect 454727 4913 454739 4947
rect 454681 4907 454739 4913
rect 458082 4904 458088 4956
rect 458140 4944 458146 4956
rect 466089 4947 466147 4953
rect 466089 4944 466101 4947
rect 458140 4916 466101 4944
rect 458140 4904 458146 4916
rect 466089 4913 466101 4916
rect 466135 4913 466147 4947
rect 466089 4907 466147 4913
rect 466178 4904 466184 4956
rect 466236 4944 466242 4956
rect 471164 4944 471192 4984
rect 565538 4972 565544 4984
rect 565596 4972 565602 5024
rect 569034 4944 569040 4956
rect 466236 4916 471100 4944
rect 471164 4916 569040 4944
rect 466236 4904 466242 4916
rect 327074 4836 327080 4888
rect 327132 4876 327138 4888
rect 361666 4876 361672 4888
rect 327132 4848 361672 4876
rect 327132 4836 327138 4848
rect 361666 4836 361672 4848
rect 361724 4836 361730 4888
rect 422202 4836 422208 4888
rect 422260 4876 422266 4888
rect 461213 4879 461271 4885
rect 461213 4876 461225 4879
rect 422260 4848 461225 4876
rect 422260 4836 422266 4848
rect 461213 4845 461225 4848
rect 461259 4845 461271 4879
rect 469122 4876 469128 4888
rect 461213 4839 461271 4845
rect 461596 4848 469128 4876
rect 325191 4780 326568 4808
rect 326617 4811 326675 4817
rect 325191 4777 325203 4780
rect 325145 4771 325203 4777
rect 326617 4777 326629 4811
rect 326663 4808 326675 4811
rect 327169 4811 327227 4817
rect 327169 4808 327181 4811
rect 326663 4780 327181 4808
rect 326663 4777 326675 4780
rect 326617 4771 326675 4777
rect 327169 4777 327181 4780
rect 327215 4777 327227 4811
rect 327169 4771 327227 4777
rect 328454 4768 328460 4820
rect 328512 4808 328518 4820
rect 363046 4808 363052 4820
rect 328512 4780 363052 4808
rect 328512 4768 328518 4780
rect 363046 4768 363052 4780
rect 363104 4768 363110 4820
rect 423582 4768 423588 4820
rect 423640 4808 423646 4820
rect 461596 4808 461624 4848
rect 469122 4836 469128 4848
rect 469180 4836 469186 4888
rect 471072 4876 471100 4916
rect 569034 4904 569040 4916
rect 569092 4904 569098 4956
rect 572622 4876 572628 4888
rect 471072 4848 572628 4876
rect 572622 4836 572628 4848
rect 572680 4836 572686 4888
rect 423640 4780 461624 4808
rect 423640 4768 423646 4780
rect 462130 4768 462136 4820
rect 462188 4808 462194 4820
rect 471333 4811 471391 4817
rect 471333 4808 471345 4811
rect 462188 4780 471345 4808
rect 462188 4768 462194 4780
rect 471333 4777 471345 4780
rect 471379 4777 471391 4811
rect 471333 4771 471391 4777
rect 471425 4811 471483 4817
rect 471425 4777 471437 4811
rect 471471 4808 471483 4811
rect 579798 4808 579804 4820
rect 471471 4780 579804 4808
rect 471471 4777 471483 4780
rect 471425 4771 471483 4777
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 324314 4740 324320 4752
rect 320192 4712 324320 4740
rect 320085 4703 320143 4709
rect 324314 4700 324320 4712
rect 324372 4700 324378 4752
rect 358998 4740 359004 4752
rect 324424 4712 359004 4740
rect 215846 4632 215852 4684
rect 215904 4672 215910 4684
rect 317414 4672 317420 4684
rect 215904 4644 317420 4672
rect 215904 4632 215910 4644
rect 317414 4632 317420 4644
rect 317472 4632 317478 4684
rect 321554 4672 321560 4684
rect 318904 4644 321560 4672
rect 219342 4564 219348 4616
rect 219400 4604 219406 4616
rect 318794 4604 318800 4616
rect 219400 4576 318800 4604
rect 219400 4564 219406 4576
rect 318794 4564 318800 4576
rect 318852 4564 318858 4616
rect 222930 4496 222936 4548
rect 222988 4536 222994 4548
rect 318904 4536 318932 4644
rect 321554 4632 321560 4644
rect 321612 4632 321618 4684
rect 324222 4632 324228 4684
rect 324280 4672 324286 4684
rect 324424 4672 324452 4712
rect 358998 4700 359004 4712
rect 359056 4700 359062 4752
rect 451090 4700 451096 4752
rect 451148 4740 451154 4752
rect 536926 4740 536932 4752
rect 451148 4712 536932 4740
rect 451148 4700 451154 4712
rect 536926 4700 536932 4712
rect 536984 4700 536990 4752
rect 324280 4644 324452 4672
rect 326341 4675 326399 4681
rect 324280 4632 324286 4644
rect 326341 4641 326353 4675
rect 326387 4641 326399 4675
rect 326341 4635 326399 4641
rect 322934 4604 322940 4616
rect 222988 4508 318932 4536
rect 319456 4576 322940 4604
rect 222988 4496 222994 4508
rect 226518 4428 226524 4480
rect 226576 4468 226582 4480
rect 319456 4468 319484 4576
rect 322934 4564 322940 4576
rect 322992 4564 322998 4616
rect 324133 4607 324191 4613
rect 324133 4573 324145 4607
rect 324179 4604 324191 4607
rect 326249 4607 326307 4613
rect 326249 4604 326261 4607
rect 324179 4576 326261 4604
rect 324179 4573 324191 4576
rect 324133 4567 324191 4573
rect 326249 4573 326261 4576
rect 326295 4573 326307 4607
rect 326356 4604 326384 4635
rect 326522 4632 326528 4684
rect 326580 4672 326586 4684
rect 360470 4672 360476 4684
rect 326580 4644 360476 4672
rect 326580 4632 326586 4644
rect 360470 4632 360476 4644
rect 360528 4632 360534 4684
rect 449802 4632 449808 4684
rect 449860 4672 449866 4684
rect 533430 4672 533436 4684
rect 449860 4644 533436 4672
rect 449860 4632 449866 4644
rect 533430 4632 533436 4644
rect 533488 4632 533494 4684
rect 333974 4604 333980 4616
rect 326356 4576 333980 4604
rect 326249 4567 326307 4573
rect 333974 4564 333980 4576
rect 334032 4564 334038 4616
rect 448330 4564 448336 4616
rect 448388 4604 448394 4616
rect 529842 4604 529848 4616
rect 448388 4576 529848 4604
rect 448388 4564 448394 4576
rect 529842 4564 529848 4576
rect 529900 4564 529906 4616
rect 320085 4539 320143 4545
rect 320085 4505 320097 4539
rect 320131 4536 320143 4539
rect 320913 4539 320971 4545
rect 320913 4536 320925 4539
rect 320131 4508 320925 4536
rect 320131 4505 320143 4508
rect 320085 4499 320143 4505
rect 320913 4505 320925 4508
rect 320959 4505 320971 4539
rect 320913 4499 320971 4505
rect 322842 4496 322848 4548
rect 322900 4536 322906 4548
rect 337010 4536 337016 4548
rect 322900 4508 337016 4536
rect 322900 4496 322906 4508
rect 337010 4496 337016 4508
rect 337068 4496 337074 4548
rect 350537 4539 350595 4545
rect 350537 4505 350549 4539
rect 350583 4536 350595 4539
rect 353478 4536 353484 4548
rect 350583 4508 353484 4536
rect 350583 4505 350595 4508
rect 350537 4499 350595 4505
rect 353478 4496 353484 4508
rect 353536 4496 353542 4548
rect 447042 4496 447048 4548
rect 447100 4536 447106 4548
rect 526254 4536 526260 4548
rect 447100 4508 526260 4536
rect 447100 4496 447106 4508
rect 526254 4496 526260 4508
rect 526312 4496 526318 4548
rect 226576 4440 319484 4468
rect 226576 4428 226582 4440
rect 320358 4428 320364 4480
rect 320416 4468 320422 4480
rect 335354 4468 335360 4480
rect 320416 4440 335360 4468
rect 320416 4428 320422 4440
rect 335354 4428 335360 4440
rect 335412 4428 335418 4480
rect 350169 4471 350227 4477
rect 350169 4437 350181 4471
rect 350215 4468 350227 4471
rect 352558 4468 352564 4480
rect 350215 4440 352564 4468
rect 350215 4437 350227 4440
rect 350169 4431 350227 4437
rect 352558 4428 352564 4440
rect 352616 4428 352622 4480
rect 445570 4428 445576 4480
rect 445628 4468 445634 4480
rect 522666 4468 522672 4480
rect 445628 4440 522672 4468
rect 445628 4428 445634 4440
rect 522666 4428 522672 4440
rect 522724 4428 522730 4480
rect 201494 4360 201500 4412
rect 201552 4400 201558 4412
rect 271138 4400 271144 4412
rect 201552 4372 271144 4400
rect 201552 4360 201558 4372
rect 271138 4360 271144 4372
rect 271196 4360 271202 4412
rect 301406 4360 301412 4412
rect 301464 4400 301470 4412
rect 350537 4403 350595 4409
rect 350537 4400 350549 4403
rect 301464 4372 350549 4400
rect 301464 4360 301470 4372
rect 350537 4369 350549 4372
rect 350583 4369 350595 4403
rect 350537 4363 350595 4369
rect 351273 4403 351331 4409
rect 351273 4369 351285 4403
rect 351319 4400 351331 4403
rect 355318 4400 355324 4412
rect 351319 4372 355324 4400
rect 351319 4369 351331 4372
rect 351273 4363 351331 4369
rect 355318 4360 355324 4372
rect 355376 4360 355382 4412
rect 376757 4403 376815 4409
rect 376757 4369 376769 4403
rect 376803 4400 376815 4403
rect 380158 4400 380164 4412
rect 376803 4372 380164 4400
rect 376803 4369 376815 4372
rect 376757 4363 376815 4369
rect 380158 4360 380164 4372
rect 380216 4360 380222 4412
rect 444282 4360 444288 4412
rect 444340 4400 444346 4412
rect 519078 4400 519084 4412
rect 444340 4372 519084 4400
rect 444340 4360 444346 4372
rect 519078 4360 519084 4372
rect 519136 4360 519142 4412
rect 205082 4292 205088 4344
rect 205140 4332 205146 4344
rect 272518 4332 272524 4344
rect 205140 4304 272524 4332
rect 205140 4292 205146 4304
rect 272518 4292 272524 4304
rect 272576 4292 272582 4344
rect 304994 4292 305000 4344
rect 305052 4332 305058 4344
rect 354950 4332 354956 4344
rect 305052 4304 354956 4332
rect 305052 4292 305058 4304
rect 354950 4292 354956 4304
rect 355008 4292 355014 4344
rect 442902 4292 442908 4344
rect 442960 4332 442966 4344
rect 515582 4332 515588 4344
rect 442960 4304 515588 4332
rect 442960 4292 442966 4304
rect 515582 4292 515588 4304
rect 515640 4292 515646 4344
rect 220265 4267 220323 4273
rect 220265 4233 220277 4267
rect 220311 4264 220323 4267
rect 229094 4264 229100 4276
rect 220311 4236 229100 4264
rect 220311 4233 220323 4236
rect 220265 4227 220323 4233
rect 229094 4224 229100 4236
rect 229152 4224 229158 4276
rect 249061 4267 249119 4273
rect 249061 4233 249073 4267
rect 249107 4264 249119 4267
rect 258721 4267 258779 4273
rect 258721 4264 258733 4267
rect 249107 4236 258733 4264
rect 249107 4233 249119 4236
rect 249061 4227 249119 4233
rect 258721 4233 258733 4236
rect 258767 4233 258779 4267
rect 258721 4227 258779 4233
rect 308582 4224 308588 4276
rect 308640 4264 308646 4276
rect 356146 4264 356152 4276
rect 308640 4236 356152 4264
rect 308640 4224 308646 4236
rect 356146 4224 356152 4236
rect 356204 4224 356210 4276
rect 441522 4224 441528 4276
rect 441580 4264 441586 4276
rect 511994 4264 512000 4276
rect 441580 4236 512000 4264
rect 441580 4224 441586 4236
rect 511994 4224 512000 4236
rect 512052 4224 512058 4276
rect 124214 4156 124220 4208
rect 124272 4196 124278 4208
rect 125410 4196 125416 4208
rect 124272 4168 125416 4196
rect 124272 4156 124278 4168
rect 125410 4156 125416 4168
rect 125468 4156 125474 4208
rect 140866 4156 140872 4208
rect 140924 4196 140930 4208
rect 142062 4196 142068 4208
rect 140924 4168 142068 4196
rect 140924 4156 140930 4168
rect 142062 4156 142068 4168
rect 142120 4156 142126 4208
rect 150434 4156 150440 4208
rect 150492 4196 150498 4208
rect 151630 4196 151636 4208
rect 150492 4168 151636 4196
rect 150492 4156 150498 4168
rect 151630 4156 151636 4168
rect 151688 4156 151694 4208
rect 158714 4156 158720 4208
rect 158772 4196 158778 4208
rect 160002 4196 160008 4208
rect 158772 4168 160008 4196
rect 158772 4156 158778 4168
rect 160002 4156 160008 4168
rect 160060 4156 160066 4208
rect 175366 4156 175372 4208
rect 175424 4196 175430 4208
rect 176562 4196 176568 4208
rect 175424 4168 176568 4196
rect 175424 4156 175430 4168
rect 176562 4156 176568 4168
rect 176620 4156 176626 4208
rect 209866 4156 209872 4208
rect 209924 4196 209930 4208
rect 211062 4196 211068 4208
rect 209924 4168 211068 4196
rect 209924 4156 209930 4168
rect 211062 4156 211068 4168
rect 211120 4156 211126 4208
rect 287609 4199 287667 4205
rect 284680 4168 285720 4196
rect 34974 4088 34980 4140
rect 35032 4128 35038 4140
rect 50338 4128 50344 4140
rect 35032 4100 50344 4128
rect 35032 4088 35038 4100
rect 50338 4088 50344 4100
rect 50396 4088 50402 4140
rect 57606 4088 57612 4140
rect 57664 4128 57670 4140
rect 250438 4128 250444 4140
rect 57664 4100 250444 4128
rect 57664 4088 57670 4100
rect 250438 4088 250444 4100
rect 250496 4088 250502 4140
rect 268102 4088 268108 4140
rect 268160 4128 268166 4140
rect 269022 4128 269028 4140
rect 268160 4100 269028 4128
rect 268160 4088 268166 4100
rect 269022 4088 269028 4100
rect 269080 4088 269086 4140
rect 278041 4131 278099 4137
rect 278041 4097 278053 4131
rect 278087 4128 278099 4131
rect 284680 4128 284708 4168
rect 278087 4100 284708 4128
rect 278087 4097 278099 4100
rect 278041 4091 278099 4097
rect 284754 4088 284760 4140
rect 284812 4128 284818 4140
rect 285582 4128 285588 4140
rect 284812 4100 285588 4128
rect 284812 4088 284818 4100
rect 285582 4088 285588 4100
rect 285640 4088 285646 4140
rect 285692 4128 285720 4168
rect 287609 4165 287621 4199
rect 287655 4196 287667 4199
rect 307021 4199 307079 4205
rect 287655 4168 287928 4196
rect 287655 4165 287667 4168
rect 287609 4159 287667 4165
rect 287900 4128 287928 4168
rect 307021 4165 307033 4199
rect 307067 4196 307079 4199
rect 312078 4196 312084 4208
rect 307067 4168 312084 4196
rect 307067 4165 307079 4168
rect 307021 4159 307079 4165
rect 312078 4156 312084 4168
rect 312136 4156 312142 4208
rect 312170 4156 312176 4208
rect 312228 4196 312234 4208
rect 357802 4196 357808 4208
rect 312228 4168 357808 4196
rect 312228 4156 312234 4168
rect 357802 4156 357808 4168
rect 357860 4156 357866 4208
rect 424962 4156 424968 4208
rect 425020 4196 425026 4208
rect 472710 4196 472716 4208
rect 425020 4168 472716 4196
rect 425020 4156 425026 4168
rect 472710 4156 472716 4168
rect 472768 4156 472774 4208
rect 295886 4128 295892 4140
rect 285692 4100 287836 4128
rect 287900 4100 295892 4128
rect 20714 4020 20720 4072
rect 20772 4060 20778 4072
rect 28258 4060 28264 4072
rect 20772 4032 28264 4060
rect 20772 4020 20778 4032
rect 28258 4020 28264 4032
rect 28316 4020 28322 4072
rect 50522 4020 50528 4072
rect 50580 4060 50586 4072
rect 249058 4060 249064 4072
rect 50580 4032 249064 4060
rect 50580 4020 50586 4032
rect 249058 4020 249064 4032
rect 249116 4020 249122 4072
rect 263873 4063 263931 4069
rect 263873 4029 263885 4063
rect 263919 4060 263931 4063
rect 282917 4063 282975 4069
rect 282917 4060 282929 4063
rect 263919 4032 282929 4060
rect 263919 4029 263931 4032
rect 263873 4023 263931 4029
rect 282917 4029 282929 4032
rect 282963 4029 282975 4063
rect 287808 4060 287836 4100
rect 295886 4088 295892 4100
rect 295944 4088 295950 4140
rect 296714 4088 296720 4140
rect 296772 4128 296778 4140
rect 297910 4128 297916 4140
rect 296772 4100 297916 4128
rect 296772 4088 296778 4100
rect 297910 4088 297916 4100
rect 297968 4088 297974 4140
rect 300302 4088 300308 4140
rect 300360 4128 300366 4140
rect 342898 4128 342904 4140
rect 300360 4100 342904 4128
rect 300360 4088 300366 4100
rect 342898 4088 342904 4100
rect 342956 4088 342962 4140
rect 343634 4088 343640 4140
rect 343692 4128 343698 4140
rect 344278 4128 344284 4140
rect 343692 4100 344284 4128
rect 343692 4088 343698 4100
rect 344278 4088 344284 4100
rect 344336 4088 344342 4140
rect 347866 4088 347872 4140
rect 347924 4128 347930 4140
rect 349062 4128 349068 4140
rect 347924 4100 349068 4128
rect 347924 4088 347930 4100
rect 349062 4088 349068 4100
rect 349120 4088 349126 4140
rect 349157 4131 349215 4137
rect 349157 4097 349169 4131
rect 349203 4128 349215 4131
rect 351273 4131 351331 4137
rect 351273 4128 351285 4131
rect 349203 4100 351285 4128
rect 349203 4097 349215 4100
rect 349157 4091 349215 4097
rect 351273 4097 351285 4100
rect 351319 4097 351331 4131
rect 351273 4091 351331 4097
rect 351362 4088 351368 4140
rect 351420 4128 351426 4140
rect 351822 4128 351828 4140
rect 351420 4100 351828 4128
rect 351420 4088 351426 4100
rect 351822 4088 351828 4100
rect 351880 4088 351886 4140
rect 352558 4088 352564 4140
rect 352616 4128 352622 4140
rect 354309 4131 354367 4137
rect 352616 4100 354260 4128
rect 352616 4088 352622 4100
rect 298094 4060 298100 4072
rect 287808 4032 298100 4060
rect 282917 4023 282975 4029
rect 298094 4020 298100 4032
rect 298152 4020 298158 4072
rect 302602 4020 302608 4072
rect 302660 4060 302666 4072
rect 309778 4060 309784 4072
rect 302660 4032 309784 4060
rect 302660 4020 302666 4032
rect 309778 4020 309784 4032
rect 309836 4020 309842 4072
rect 314562 4020 314568 4072
rect 314620 4060 314626 4072
rect 350626 4060 350632 4072
rect 314620 4032 350632 4060
rect 314620 4020 314626 4032
rect 350626 4020 350632 4032
rect 350684 4020 350690 4072
rect 46934 3952 46940 4004
rect 46992 3992 46998 4004
rect 248690 3992 248696 4004
rect 46992 3964 248696 3992
rect 46992 3952 46998 3964
rect 248690 3952 248696 3964
rect 248748 3952 248754 4004
rect 257430 3952 257436 4004
rect 257488 3992 257494 4004
rect 287609 3995 287667 4001
rect 287609 3992 287621 3995
rect 257488 3964 287621 3992
rect 257488 3952 257494 3964
rect 287609 3961 287621 3964
rect 287655 3961 287667 3995
rect 287609 3955 287667 3961
rect 287701 3995 287759 4001
rect 287701 3961 287713 3995
rect 287747 3992 287759 3995
rect 297358 3992 297364 4004
rect 287747 3964 297364 3992
rect 287747 3961 287759 3964
rect 287701 3955 287759 3961
rect 297358 3952 297364 3964
rect 297416 3952 297422 4004
rect 313366 3952 313372 4004
rect 313424 3992 313430 4004
rect 350534 3992 350540 4004
rect 313424 3964 350540 3992
rect 313424 3952 313430 3964
rect 350534 3952 350540 3964
rect 350592 3952 350598 4004
rect 354232 3992 354260 4100
rect 354309 4097 354321 4131
rect 354355 4128 354367 4131
rect 360841 4131 360899 4137
rect 360841 4128 360853 4131
rect 354355 4100 360853 4128
rect 354355 4097 354367 4100
rect 354309 4091 354367 4097
rect 360841 4097 360853 4100
rect 360887 4097 360899 4131
rect 360841 4091 360899 4097
rect 360930 4088 360936 4140
rect 360988 4128 360994 4140
rect 360988 4100 362448 4128
rect 360988 4088 360994 4100
rect 357434 4020 357440 4072
rect 357492 4060 357498 4072
rect 358078 4060 358084 4072
rect 357492 4032 358084 4060
rect 357492 4020 357498 4032
rect 358078 4020 358084 4032
rect 358136 4020 358142 4072
rect 358170 4020 358176 4072
rect 358228 4060 358234 4072
rect 362218 4060 362224 4072
rect 358228 4032 362224 4060
rect 358228 4020 358234 4032
rect 362218 4020 362224 4032
rect 362276 4020 362282 4072
rect 362420 4060 362448 4100
rect 363322 4088 363328 4140
rect 363380 4128 363386 4140
rect 364242 4128 364248 4140
rect 363380 4100 364248 4128
rect 363380 4088 363386 4100
rect 364242 4088 364248 4100
rect 364300 4088 364306 4140
rect 369210 4088 369216 4140
rect 369268 4128 369274 4140
rect 369762 4128 369768 4140
rect 369268 4100 369768 4128
rect 369268 4088 369274 4100
rect 369762 4088 369768 4100
rect 369820 4088 369826 4140
rect 370406 4088 370412 4140
rect 370464 4128 370470 4140
rect 371142 4128 371148 4140
rect 370464 4100 371148 4128
rect 370464 4088 370470 4100
rect 371142 4088 371148 4100
rect 371200 4088 371206 4140
rect 377582 4088 377588 4140
rect 377640 4128 377646 4140
rect 378042 4128 378048 4140
rect 377640 4100 378048 4128
rect 377640 4088 377646 4100
rect 378042 4088 378048 4100
rect 378100 4088 378106 4140
rect 378778 4088 378784 4140
rect 378836 4128 378842 4140
rect 385310 4128 385316 4140
rect 378836 4100 385316 4128
rect 378836 4088 378842 4100
rect 385310 4088 385316 4100
rect 385368 4088 385374 4140
rect 390830 4088 390836 4140
rect 390888 4128 390894 4140
rect 391842 4128 391848 4140
rect 390888 4100 391848 4128
rect 390888 4088 390894 4100
rect 391842 4088 391848 4100
rect 391900 4088 391906 4140
rect 393130 4088 393136 4140
rect 393188 4128 393194 4140
rect 395430 4128 395436 4140
rect 393188 4100 395436 4128
rect 393188 4088 393194 4100
rect 395430 4088 395436 4100
rect 395488 4088 395494 4140
rect 398098 4088 398104 4140
rect 398156 4128 398162 4140
rect 404906 4128 404912 4140
rect 398156 4100 404912 4128
rect 398156 4088 398162 4100
rect 404906 4088 404912 4100
rect 404964 4088 404970 4140
rect 411070 4088 411076 4140
rect 411128 4128 411134 4140
rect 438210 4128 438216 4140
rect 411128 4100 438216 4128
rect 411128 4088 411134 4100
rect 438210 4088 438216 4100
rect 438268 4088 438274 4140
rect 442258 4088 442264 4140
rect 442316 4128 442322 4140
rect 445573 4131 445631 4137
rect 445573 4128 445585 4131
rect 442316 4100 445585 4128
rect 442316 4088 442322 4100
rect 445573 4097 445585 4100
rect 445619 4097 445631 4131
rect 445573 4091 445631 4097
rect 445662 4088 445668 4140
rect 445720 4128 445726 4140
rect 521470 4128 521476 4140
rect 445720 4100 521476 4128
rect 445720 4088 445726 4100
rect 521470 4088 521476 4100
rect 521528 4088 521534 4140
rect 529198 4088 529204 4140
rect 529256 4128 529262 4140
rect 575014 4128 575020 4140
rect 529256 4100 575020 4128
rect 529256 4088 529262 4100
rect 575014 4088 575020 4100
rect 575072 4088 575078 4140
rect 377398 4060 377404 4072
rect 362420 4032 377404 4060
rect 377398 4020 377404 4032
rect 377456 4020 377462 4072
rect 379974 4020 379980 4072
rect 380032 4060 380038 4072
rect 380802 4060 380808 4072
rect 380032 4032 380808 4060
rect 380032 4020 380038 4032
rect 380802 4020 380808 4032
rect 380860 4020 380866 4072
rect 381170 4020 381176 4072
rect 381228 4060 381234 4072
rect 382182 4060 382188 4072
rect 381228 4032 382188 4060
rect 381228 4020 381234 4032
rect 382182 4020 382188 4032
rect 382240 4020 382246 4072
rect 383562 4020 383568 4072
rect 383620 4060 383626 4072
rect 384298 4060 384304 4072
rect 383620 4032 384304 4060
rect 383620 4020 383626 4032
rect 384298 4020 384304 4032
rect 384356 4020 384362 4072
rect 393222 4020 393228 4072
rect 393280 4060 393286 4072
rect 396626 4060 396632 4072
rect 393280 4032 396632 4060
rect 393280 4020 393286 4032
rect 396626 4020 396632 4032
rect 396684 4020 396690 4072
rect 411162 4020 411168 4072
rect 411220 4060 411226 4072
rect 439406 4060 439412 4072
rect 411220 4032 439412 4060
rect 411220 4020 411226 4032
rect 439406 4020 439412 4032
rect 439464 4020 439470 4072
rect 439498 4020 439504 4072
rect 439556 4060 439562 4072
rect 446309 4063 446367 4069
rect 446309 4060 446321 4063
rect 439556 4032 446321 4060
rect 439556 4020 439562 4032
rect 446309 4029 446321 4032
rect 446355 4029 446367 4063
rect 446309 4023 446367 4029
rect 448422 4020 448428 4072
rect 448480 4060 448486 4072
rect 528646 4060 528652 4072
rect 448480 4032 528652 4060
rect 448480 4020 448486 4032
rect 528646 4020 528652 4032
rect 528704 4020 528710 4072
rect 530578 4020 530584 4072
rect 530636 4060 530642 4072
rect 582190 4060 582196 4072
rect 530636 4032 582196 4060
rect 530636 4020 530642 4032
rect 582190 4020 582196 4032
rect 582248 4020 582254 4072
rect 359553 3995 359611 4001
rect 359553 3992 359565 3995
rect 354232 3964 359565 3992
rect 359553 3961 359565 3964
rect 359599 3961 359611 3995
rect 359553 3955 359611 3961
rect 369765 3995 369823 4001
rect 369765 3961 369777 3995
rect 369811 3992 369823 3995
rect 377122 3992 377128 4004
rect 369811 3964 377128 3992
rect 369811 3961 369823 3964
rect 369765 3955 369823 3961
rect 377122 3952 377128 3964
rect 377180 3952 377186 4004
rect 402790 3952 402796 4004
rect 402848 3992 402854 4004
rect 419166 3992 419172 4004
rect 402848 3964 419172 3992
rect 402848 3952 402854 3964
rect 419166 3952 419172 3964
rect 419224 3952 419230 4004
rect 421558 3952 421564 4004
rect 421616 3992 421622 4004
rect 450170 3992 450176 4004
rect 421616 3964 450176 3992
rect 421616 3952 421622 3964
rect 450170 3952 450176 3964
rect 450228 3952 450234 4004
rect 451182 3952 451188 4004
rect 451240 3992 451246 4004
rect 535730 3992 535736 4004
rect 451240 3964 535736 3992
rect 451240 3952 451246 3964
rect 535730 3952 535736 3964
rect 535788 3952 535794 4004
rect 45738 3884 45744 3936
rect 45796 3924 45802 3936
rect 247678 3924 247684 3936
rect 45796 3896 247684 3924
rect 45796 3884 45802 3896
rect 247678 3884 247684 3896
rect 247736 3884 247742 3936
rect 282454 3884 282460 3936
rect 282512 3924 282518 3936
rect 318889 3927 318947 3933
rect 318889 3924 318901 3927
rect 282512 3896 318901 3924
rect 282512 3884 282518 3896
rect 318889 3893 318901 3896
rect 318935 3893 318947 3927
rect 318889 3887 318947 3893
rect 318981 3927 319039 3933
rect 318981 3893 318993 3927
rect 319027 3924 319039 3927
rect 325602 3924 325608 3936
rect 319027 3896 325608 3924
rect 319027 3893 319039 3896
rect 318981 3887 319039 3893
rect 325602 3884 325608 3896
rect 325660 3884 325666 3936
rect 326430 3884 326436 3936
rect 326488 3924 326494 3936
rect 328454 3924 328460 3936
rect 326488 3896 328460 3924
rect 326488 3884 326494 3896
rect 328454 3884 328460 3896
rect 328512 3884 328518 3936
rect 328822 3884 328828 3936
rect 328880 3924 328886 3936
rect 354122 3924 354128 3936
rect 328880 3896 354128 3924
rect 328880 3884 328886 3896
rect 354122 3884 354128 3896
rect 354180 3884 354186 3936
rect 354214 3884 354220 3936
rect 354272 3924 354278 3936
rect 359090 3924 359096 3936
rect 354272 3896 359096 3924
rect 354272 3884 354278 3896
rect 359090 3884 359096 3896
rect 359148 3884 359154 3936
rect 359734 3884 359740 3936
rect 359792 3924 359798 3936
rect 360749 3927 360807 3933
rect 360749 3924 360761 3927
rect 359792 3896 360761 3924
rect 359792 3884 359798 3896
rect 360749 3893 360761 3896
rect 360795 3893 360807 3927
rect 360749 3887 360807 3893
rect 360841 3927 360899 3933
rect 360841 3893 360853 3927
rect 360887 3924 360899 3927
rect 374086 3924 374092 3936
rect 360887 3896 374092 3924
rect 360887 3893 360899 3896
rect 360841 3887 360899 3893
rect 374086 3884 374092 3896
rect 374144 3884 374150 3936
rect 412450 3884 412456 3936
rect 412508 3924 412514 3936
rect 441798 3924 441804 3936
rect 412508 3896 441804 3924
rect 412508 3884 412514 3896
rect 441798 3884 441804 3896
rect 441856 3884 441862 3936
rect 442350 3884 442356 3936
rect 442408 3924 442414 3936
rect 445481 3927 445539 3933
rect 445481 3924 445493 3927
rect 442408 3896 445493 3924
rect 442408 3884 442414 3896
rect 445481 3893 445493 3896
rect 445527 3893 445539 3927
rect 445481 3887 445539 3893
rect 445573 3927 445631 3933
rect 445573 3893 445585 3927
rect 445619 3924 445631 3927
rect 446306 3924 446312 3936
rect 445619 3896 446312 3924
rect 445619 3893 445631 3896
rect 445573 3887 445631 3893
rect 446306 3884 446312 3896
rect 446364 3884 446370 3936
rect 446401 3927 446459 3933
rect 446401 3893 446413 3927
rect 446447 3924 446459 3927
rect 453666 3924 453672 3936
rect 446447 3896 453672 3924
rect 446447 3893 446459 3896
rect 446401 3887 446459 3893
rect 453666 3884 453672 3896
rect 453724 3884 453730 3936
rect 453942 3884 453948 3936
rect 454000 3924 454006 3936
rect 542906 3924 542912 3936
rect 454000 3896 542912 3924
rect 454000 3884 454006 3896
rect 542906 3884 542912 3896
rect 542964 3884 542970 3936
rect 39758 3816 39764 3868
rect 39816 3856 39822 3868
rect 245930 3856 245936 3868
rect 39816 3828 245936 3856
rect 39816 3816 39822 3828
rect 245930 3816 245936 3828
rect 245988 3816 245994 3868
rect 264606 3816 264612 3868
rect 264664 3856 264670 3868
rect 278041 3859 278099 3865
rect 278041 3856 278053 3859
rect 264664 3828 278053 3856
rect 264664 3816 264670 3828
rect 278041 3825 278053 3828
rect 278087 3825 278099 3859
rect 278041 3819 278099 3825
rect 285950 3816 285956 3868
rect 286008 3856 286014 3868
rect 331401 3859 331459 3865
rect 331401 3856 331413 3859
rect 286008 3828 331413 3856
rect 286008 3816 286014 3828
rect 331401 3825 331413 3828
rect 331447 3825 331459 3859
rect 331401 3819 331459 3825
rect 332410 3816 332416 3868
rect 332468 3856 332474 3868
rect 333238 3856 333244 3868
rect 332468 3828 333244 3856
rect 332468 3816 332474 3828
rect 333238 3816 333244 3828
rect 333296 3816 333302 3868
rect 334710 3816 334716 3868
rect 334768 3856 334774 3868
rect 335262 3856 335268 3868
rect 334768 3828 335268 3856
rect 334768 3816 334774 3828
rect 335262 3816 335268 3828
rect 335320 3816 335326 3868
rect 338209 3859 338267 3865
rect 338209 3825 338221 3859
rect 338255 3856 338267 3859
rect 338758 3856 338764 3868
rect 338255 3828 338764 3856
rect 338255 3825 338267 3828
rect 338209 3819 338267 3825
rect 338758 3816 338764 3828
rect 338816 3816 338822 3868
rect 341518 3856 341524 3868
rect 338960 3828 341524 3856
rect 19518 3748 19524 3800
rect 19576 3788 19582 3800
rect 32398 3788 32404 3800
rect 19576 3760 32404 3788
rect 19576 3748 19582 3760
rect 32398 3748 32404 3760
rect 32456 3748 32462 3800
rect 38562 3748 38568 3800
rect 38620 3788 38626 3800
rect 245746 3788 245752 3800
rect 38620 3760 245752 3788
rect 38620 3748 38626 3760
rect 245746 3748 245752 3760
rect 245804 3748 245810 3800
rect 282917 3791 282975 3797
rect 282917 3757 282929 3791
rect 282963 3788 282975 3791
rect 287701 3791 287759 3797
rect 287701 3788 287713 3791
rect 282963 3760 287713 3788
rect 282963 3757 282975 3760
rect 282917 3751 282975 3757
rect 287701 3757 287713 3760
rect 287747 3757 287759 3791
rect 287701 3751 287759 3757
rect 289538 3748 289544 3800
rect 289596 3788 289602 3800
rect 332321 3791 332379 3797
rect 332321 3788 332333 3791
rect 289596 3760 332333 3788
rect 289596 3748 289602 3760
rect 332321 3757 332333 3760
rect 332367 3757 332379 3791
rect 332321 3751 332379 3757
rect 332505 3791 332563 3797
rect 332505 3757 332517 3791
rect 332551 3788 332563 3791
rect 338960 3788 338988 3828
rect 341518 3816 341524 3828
rect 341576 3816 341582 3868
rect 341886 3816 341892 3868
rect 341944 3856 341950 3868
rect 370130 3856 370136 3868
rect 341944 3828 370136 3856
rect 341944 3816 341950 3828
rect 370130 3816 370136 3828
rect 370188 3816 370194 3868
rect 372798 3816 372804 3868
rect 372856 3856 372862 3868
rect 373902 3856 373908 3868
rect 372856 3828 373908 3856
rect 372856 3816 372862 3828
rect 373902 3816 373908 3828
rect 373960 3816 373966 3868
rect 412542 3816 412548 3868
rect 412600 3856 412606 3868
rect 442994 3856 443000 3868
rect 412600 3828 443000 3856
rect 412600 3816 412606 3828
rect 442994 3816 443000 3828
rect 443052 3816 443058 3868
rect 443638 3816 443644 3868
rect 443696 3856 443702 3868
rect 446493 3859 446551 3865
rect 446493 3856 446505 3859
rect 443696 3828 446505 3856
rect 443696 3816 443702 3828
rect 446493 3825 446505 3828
rect 446539 3825 446551 3859
rect 446493 3819 446551 3825
rect 446582 3816 446588 3868
rect 446640 3856 446646 3868
rect 452470 3856 452476 3868
rect 446640 3828 452476 3856
rect 446640 3816 446646 3828
rect 452470 3816 452476 3828
rect 452528 3816 452534 3868
rect 460201 3859 460259 3865
rect 460201 3825 460213 3859
rect 460247 3825 460259 3859
rect 460201 3819 460259 3825
rect 466365 3859 466423 3865
rect 466365 3825 466377 3859
rect 466411 3856 466423 3859
rect 550082 3856 550088 3868
rect 466411 3828 550088 3856
rect 466411 3825 466423 3828
rect 466365 3819 466423 3825
rect 332551 3760 338988 3788
rect 332551 3757 332563 3760
rect 332505 3751 332563 3757
rect 343082 3748 343088 3800
rect 343140 3788 343146 3800
rect 361853 3791 361911 3797
rect 361853 3788 361865 3791
rect 343140 3760 361865 3788
rect 343140 3748 343146 3760
rect 361853 3757 361865 3760
rect 361899 3757 361911 3791
rect 368658 3788 368664 3800
rect 361853 3751 361911 3757
rect 361960 3760 368664 3788
rect 32674 3680 32680 3732
rect 32732 3720 32738 3732
rect 243078 3720 243084 3732
rect 32732 3692 243084 3720
rect 32732 3680 32738 3692
rect 243078 3680 243084 3692
rect 243136 3680 243142 3732
rect 287609 3723 287667 3729
rect 287609 3689 287621 3723
rect 287655 3720 287667 3723
rect 326341 3723 326399 3729
rect 326341 3720 326353 3723
rect 287655 3692 326353 3720
rect 287655 3689 287667 3692
rect 287609 3683 287667 3689
rect 326341 3689 326353 3692
rect 326387 3689 326399 3723
rect 326341 3683 326399 3689
rect 327626 3680 327632 3732
rect 327684 3720 327690 3732
rect 331401 3723 331459 3729
rect 327684 3692 331260 3720
rect 327684 3680 327690 3692
rect 24302 3612 24308 3664
rect 24360 3652 24366 3664
rect 239030 3652 239036 3664
rect 24360 3624 239036 3652
rect 24360 3612 24366 3624
rect 239030 3612 239036 3624
rect 239088 3612 239094 3664
rect 265802 3612 265808 3664
rect 265860 3652 265866 3664
rect 318705 3655 318763 3661
rect 318705 3652 318717 3655
rect 265860 3624 318717 3652
rect 265860 3612 265866 3624
rect 318705 3621 318717 3624
rect 318751 3621 318763 3655
rect 322842 3652 322848 3664
rect 318705 3615 318763 3621
rect 318812 3624 322848 3652
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 19978 3584 19984 3596
rect 11296 3556 19984 3584
rect 11296 3544 11302 3556
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 25498 3544 25504 3596
rect 25556 3584 25562 3596
rect 240318 3584 240324 3596
rect 25556 3556 240324 3584
rect 25556 3544 25562 3556
rect 240318 3544 240324 3556
rect 240376 3544 240382 3596
rect 262214 3544 262220 3596
rect 262272 3584 262278 3596
rect 318812 3584 318840 3624
rect 322842 3612 322848 3624
rect 322900 3612 322906 3664
rect 322937 3655 322995 3661
rect 322937 3621 322949 3655
rect 322983 3652 322995 3655
rect 326522 3652 326528 3664
rect 322983 3624 326528 3652
rect 322983 3621 322995 3624
rect 322937 3615 322995 3621
rect 326522 3612 326528 3624
rect 326580 3612 326586 3664
rect 262272 3556 318840 3584
rect 318889 3587 318947 3593
rect 262272 3544 262278 3556
rect 318889 3553 318901 3587
rect 318935 3584 318947 3587
rect 327718 3584 327724 3596
rect 318935 3556 327724 3584
rect 318935 3553 318947 3556
rect 318889 3547 318947 3553
rect 327718 3544 327724 3556
rect 327776 3544 327782 3596
rect 331232 3584 331260 3692
rect 331401 3689 331413 3723
rect 331447 3720 331459 3723
rect 338209 3723 338267 3729
rect 338209 3720 338221 3723
rect 331447 3692 338221 3720
rect 331447 3689 331459 3692
rect 331401 3683 331459 3689
rect 338209 3689 338221 3692
rect 338255 3689 338267 3723
rect 338209 3683 338267 3689
rect 338298 3680 338304 3732
rect 338356 3720 338362 3732
rect 361960 3720 361988 3760
rect 368658 3748 368664 3760
rect 368716 3748 368722 3800
rect 373994 3748 374000 3800
rect 374052 3788 374058 3800
rect 375282 3788 375288 3800
rect 374052 3760 375288 3788
rect 374052 3748 374058 3760
rect 375282 3748 375288 3760
rect 375340 3748 375346 3800
rect 376386 3748 376392 3800
rect 376444 3788 376450 3800
rect 381630 3788 381636 3800
rect 376444 3760 381636 3788
rect 376444 3748 376450 3760
rect 381630 3748 381636 3760
rect 381688 3748 381694 3800
rect 399478 3748 399484 3800
rect 399536 3788 399542 3800
rect 408494 3788 408500 3800
rect 399536 3760 408500 3788
rect 399536 3748 399542 3760
rect 408494 3748 408500 3760
rect 408552 3748 408558 3800
rect 416682 3748 416688 3800
rect 416740 3788 416746 3800
rect 420549 3791 420607 3797
rect 416740 3760 420500 3788
rect 416740 3748 416746 3760
rect 338356 3692 361988 3720
rect 362037 3723 362095 3729
rect 338356 3680 338362 3692
rect 362037 3689 362049 3723
rect 362083 3720 362095 3723
rect 372706 3720 372712 3732
rect 362083 3692 372712 3720
rect 362083 3689 362095 3692
rect 362037 3683 362095 3689
rect 372706 3680 372712 3692
rect 372764 3680 372770 3732
rect 376849 3723 376907 3729
rect 376849 3689 376861 3723
rect 376895 3720 376907 3723
rect 379698 3720 379704 3732
rect 376895 3692 379704 3720
rect 376895 3689 376907 3692
rect 376849 3683 376907 3689
rect 379698 3680 379704 3692
rect 379756 3680 379762 3732
rect 400030 3680 400036 3732
rect 400088 3720 400094 3732
rect 412082 3720 412088 3732
rect 400088 3692 412088 3720
rect 400088 3680 400094 3692
rect 412082 3680 412088 3692
rect 412140 3680 412146 3732
rect 413097 3723 413155 3729
rect 413097 3689 413109 3723
rect 413143 3720 413155 3723
rect 420362 3720 420368 3732
rect 413143 3692 420368 3720
rect 413143 3689 413155 3692
rect 413097 3683 413155 3689
rect 420362 3680 420368 3692
rect 420420 3680 420426 3732
rect 420472 3720 420500 3760
rect 420549 3757 420561 3791
rect 420595 3788 420607 3791
rect 445386 3788 445392 3800
rect 420595 3760 445392 3788
rect 420595 3757 420607 3760
rect 420549 3751 420607 3757
rect 445386 3748 445392 3760
rect 445444 3748 445450 3800
rect 445481 3791 445539 3797
rect 445481 3757 445493 3791
rect 445527 3788 445539 3791
rect 446677 3791 446735 3797
rect 446677 3788 446689 3791
rect 445527 3760 446689 3788
rect 445527 3757 445539 3760
rect 445481 3751 445539 3757
rect 446677 3757 446689 3760
rect 446723 3757 446735 3791
rect 446677 3751 446735 3757
rect 456702 3748 456708 3800
rect 456760 3788 456766 3800
rect 460216 3788 460244 3819
rect 550082 3816 550088 3828
rect 550140 3816 550146 3868
rect 456760 3760 460244 3788
rect 456760 3748 456766 3760
rect 460290 3748 460296 3800
rect 460348 3788 460354 3800
rect 463234 3788 463240 3800
rect 460348 3760 463240 3788
rect 460348 3748 460354 3760
rect 463234 3748 463240 3760
rect 463292 3748 463298 3800
rect 557166 3788 557172 3800
rect 463344 3760 557172 3788
rect 422297 3723 422355 3729
rect 422297 3720 422309 3723
rect 420472 3692 422309 3720
rect 422297 3689 422309 3692
rect 422343 3689 422355 3723
rect 422297 3683 422355 3689
rect 431865 3723 431923 3729
rect 431865 3689 431877 3723
rect 431911 3720 431923 3723
rect 441617 3723 441675 3729
rect 441617 3720 441629 3723
rect 431911 3692 441629 3720
rect 431911 3689 431923 3692
rect 431865 3683 431923 3689
rect 441617 3689 441629 3692
rect 441663 3689 441675 3723
rect 441617 3683 441675 3689
rect 449158 3680 449164 3732
rect 449216 3720 449222 3732
rect 456797 3723 456855 3729
rect 449216 3692 452516 3720
rect 449216 3680 449222 3692
rect 331306 3612 331312 3664
rect 331364 3652 331370 3664
rect 365806 3652 365812 3664
rect 331364 3624 365812 3652
rect 331364 3612 331370 3624
rect 365806 3612 365812 3624
rect 365864 3612 365870 3664
rect 375190 3612 375196 3664
rect 375248 3652 375254 3664
rect 383838 3652 383844 3664
rect 375248 3624 383844 3652
rect 375248 3612 375254 3624
rect 383838 3612 383844 3624
rect 383896 3612 383902 3664
rect 400122 3612 400128 3664
rect 400180 3652 400186 3664
rect 413186 3652 413192 3664
rect 400180 3624 413192 3652
rect 400180 3612 400186 3624
rect 413186 3612 413192 3624
rect 413244 3612 413250 3664
rect 413922 3612 413928 3664
rect 413980 3652 413986 3664
rect 413980 3624 415808 3652
rect 413980 3612 413986 3624
rect 363598 3584 363604 3596
rect 331232 3556 363604 3584
rect 363598 3544 363604 3556
rect 363656 3544 363662 3596
rect 365714 3544 365720 3596
rect 365772 3584 365778 3596
rect 366910 3584 366916 3596
rect 365772 3556 366916 3584
rect 365772 3544 365778 3556
rect 366910 3544 366916 3556
rect 366968 3544 366974 3596
rect 371602 3544 371608 3596
rect 371660 3584 371666 3596
rect 381538 3584 381544 3596
rect 371660 3556 381544 3584
rect 371660 3544 371666 3556
rect 381538 3544 381544 3556
rect 381596 3544 381602 3596
rect 402882 3544 402888 3596
rect 402940 3584 402946 3596
rect 413097 3587 413155 3593
rect 413097 3584 413109 3587
rect 402940 3556 413109 3584
rect 402940 3544 402946 3556
rect 413097 3553 413109 3556
rect 413143 3553 413155 3587
rect 415670 3584 415676 3596
rect 413097 3547 413155 3553
rect 413204 3556 415676 3584
rect 14826 3476 14832 3528
rect 14884 3516 14890 3528
rect 234890 3516 234896 3528
rect 14884 3488 234896 3516
rect 14884 3476 14890 3488
rect 234890 3476 234896 3488
rect 234948 3476 234954 3528
rect 258626 3476 258632 3528
rect 258684 3516 258690 3528
rect 320358 3516 320364 3528
rect 258684 3488 320364 3516
rect 258684 3476 258690 3488
rect 320358 3476 320364 3488
rect 320416 3476 320422 3528
rect 320450 3476 320456 3528
rect 320508 3516 320514 3528
rect 321462 3516 321468 3528
rect 320508 3488 321468 3516
rect 320508 3476 320514 3488
rect 321462 3476 321468 3488
rect 321520 3476 321526 3528
rect 324038 3476 324044 3528
rect 324096 3516 324102 3528
rect 363138 3516 363144 3528
rect 324096 3488 363144 3516
rect 324096 3476 324102 3488
rect 363138 3476 363144 3488
rect 363196 3476 363202 3528
rect 369118 3516 369124 3528
rect 363524 3488 369124 3516
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 10318 3448 10324 3460
rect 5316 3420 10324 3448
rect 5316 3408 5322 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 16022 3408 16028 3460
rect 16080 3448 16086 3460
rect 236270 3448 236276 3460
rect 16080 3420 236276 3448
rect 16080 3408 16086 3420
rect 236270 3408 236276 3420
rect 236328 3408 236334 3460
rect 255038 3408 255044 3460
rect 255096 3448 255102 3460
rect 318702 3448 318708 3460
rect 255096 3420 318708 3448
rect 255096 3408 255102 3420
rect 318702 3408 318708 3420
rect 318760 3408 318766 3460
rect 321646 3408 321652 3460
rect 321704 3448 321710 3460
rect 361850 3448 361856 3460
rect 321704 3420 361856 3448
rect 321704 3408 321710 3420
rect 361850 3408 361856 3420
rect 361908 3408 361914 3460
rect 361945 3451 362003 3457
rect 361945 3417 361957 3451
rect 361991 3448 362003 3451
rect 363524 3448 363552 3488
rect 369118 3476 369124 3488
rect 369176 3476 369182 3528
rect 376757 3519 376815 3525
rect 376757 3485 376769 3519
rect 376803 3485 376815 3519
rect 376757 3479 376815 3485
rect 361991 3420 363552 3448
rect 361991 3417 362003 3420
rect 361945 3411 362003 3417
rect 368014 3408 368020 3460
rect 368072 3448 368078 3460
rect 376772 3448 376800 3479
rect 388254 3476 388260 3528
rect 388312 3516 388318 3528
rect 389082 3516 389088 3528
rect 388312 3488 389088 3516
rect 388312 3476 388318 3488
rect 389082 3476 389088 3488
rect 389140 3476 389146 3528
rect 394602 3476 394608 3528
rect 394660 3516 394666 3528
rect 399018 3516 399024 3528
rect 394660 3488 399024 3516
rect 394660 3476 394666 3488
rect 399018 3476 399024 3488
rect 399076 3476 399082 3528
rect 402238 3476 402244 3528
rect 402296 3516 402302 3528
rect 413204 3516 413232 3556
rect 415670 3544 415676 3556
rect 415728 3544 415734 3596
rect 415780 3584 415808 3624
rect 420270 3612 420276 3664
rect 420328 3652 420334 3664
rect 423950 3652 423956 3664
rect 420328 3624 423956 3652
rect 420328 3612 420334 3624
rect 423950 3612 423956 3624
rect 424008 3612 424014 3664
rect 424410 3612 424416 3664
rect 424468 3652 424474 3664
rect 425241 3655 425299 3661
rect 425241 3652 425253 3655
rect 424468 3624 425253 3652
rect 424468 3612 424474 3624
rect 425241 3621 425253 3624
rect 425287 3621 425299 3655
rect 425241 3615 425299 3621
rect 427078 3612 427084 3664
rect 427136 3652 427142 3664
rect 431126 3652 431132 3664
rect 427136 3624 431132 3652
rect 427136 3612 427142 3624
rect 431126 3612 431132 3624
rect 431184 3612 431190 3664
rect 431221 3655 431279 3661
rect 431221 3621 431233 3655
rect 431267 3652 431279 3655
rect 446401 3655 446459 3661
rect 446401 3652 446413 3655
rect 431267 3624 446413 3652
rect 431267 3621 431279 3624
rect 431221 3615 431279 3621
rect 446401 3621 446413 3624
rect 446447 3621 446459 3655
rect 446401 3615 446459 3621
rect 446490 3612 446496 3664
rect 446548 3652 446554 3664
rect 451921 3655 451979 3661
rect 451921 3652 451933 3655
rect 446548 3624 451933 3652
rect 446548 3612 446554 3624
rect 451921 3621 451933 3624
rect 451967 3621 451979 3655
rect 452488 3652 452516 3692
rect 456797 3689 456809 3723
rect 456843 3720 456855 3723
rect 460109 3723 460167 3729
rect 460109 3720 460121 3723
rect 456843 3692 460121 3720
rect 456843 3689 456855 3692
rect 456797 3683 456855 3689
rect 460109 3689 460121 3692
rect 460155 3689 460167 3723
rect 460109 3683 460167 3689
rect 460198 3680 460204 3732
rect 460256 3720 460262 3732
rect 461765 3723 461823 3729
rect 460256 3692 461716 3720
rect 460256 3680 460262 3692
rect 461581 3655 461639 3661
rect 461581 3652 461593 3655
rect 452488 3624 461593 3652
rect 451921 3615 451979 3621
rect 461581 3621 461593 3624
rect 461627 3621 461639 3655
rect 461688 3652 461716 3692
rect 461765 3689 461777 3723
rect 461811 3720 461823 3723
rect 463145 3723 463203 3729
rect 463145 3720 463157 3723
rect 461811 3692 463157 3720
rect 461811 3689 461823 3692
rect 461765 3683 461823 3689
rect 463145 3689 463157 3692
rect 463191 3689 463203 3723
rect 463145 3683 463203 3689
rect 463344 3652 463372 3760
rect 557166 3748 557172 3760
rect 557224 3748 557230 3800
rect 564342 3720 564348 3732
rect 461688 3624 463372 3652
rect 463436 3692 564348 3720
rect 461581 3615 461639 3621
rect 420549 3587 420607 3593
rect 420549 3584 420561 3587
rect 415780 3556 420561 3584
rect 420549 3553 420561 3556
rect 420595 3553 420607 3587
rect 420549 3547 420607 3553
rect 420822 3544 420828 3596
rect 420880 3584 420886 3596
rect 460842 3584 460848 3596
rect 420880 3556 460848 3584
rect 420880 3544 420886 3556
rect 460842 3544 460848 3556
rect 460900 3544 460906 3596
rect 460937 3587 460995 3593
rect 460937 3553 460949 3587
rect 460983 3584 460995 3587
rect 461765 3587 461823 3593
rect 461765 3584 461777 3587
rect 460983 3556 461777 3584
rect 460983 3553 460995 3556
rect 460937 3547 460995 3553
rect 461765 3553 461777 3556
rect 461811 3553 461823 3587
rect 461765 3547 461823 3553
rect 462222 3544 462228 3596
rect 462280 3584 462286 3596
rect 463436 3584 463464 3692
rect 564342 3680 564348 3692
rect 564400 3680 564406 3732
rect 463602 3612 463608 3664
rect 463660 3652 463666 3664
rect 566734 3652 566740 3664
rect 463660 3624 566740 3652
rect 463660 3612 463666 3624
rect 566734 3612 566740 3624
rect 566792 3612 566798 3664
rect 462280 3556 463464 3584
rect 463513 3587 463571 3593
rect 462280 3544 462286 3556
rect 463513 3553 463525 3587
rect 463559 3584 463571 3587
rect 466089 3587 466147 3593
rect 466089 3584 466101 3587
rect 463559 3556 466101 3584
rect 463559 3553 463571 3556
rect 463513 3547 463571 3553
rect 466089 3553 466101 3556
rect 466135 3553 466147 3587
rect 466089 3547 466147 3553
rect 466362 3544 466368 3596
rect 466420 3584 466426 3596
rect 571426 3584 571432 3596
rect 466420 3556 571432 3584
rect 466420 3544 466426 3556
rect 571426 3544 571432 3556
rect 571484 3544 571490 3596
rect 402296 3488 413232 3516
rect 402296 3476 402302 3488
rect 413278 3476 413284 3528
rect 413336 3516 413342 3528
rect 414474 3516 414480 3528
rect 413336 3488 414480 3516
rect 413336 3476 413342 3488
rect 414474 3476 414480 3488
rect 414532 3476 414538 3528
rect 418062 3476 418068 3528
rect 418120 3516 418126 3528
rect 457254 3516 457260 3528
rect 418120 3488 457260 3516
rect 418120 3476 418126 3488
rect 457254 3476 457260 3488
rect 457312 3476 457318 3528
rect 460109 3519 460167 3525
rect 460109 3485 460121 3519
rect 460155 3516 460167 3519
rect 466181 3519 466239 3525
rect 466181 3516 466193 3519
rect 460155 3488 466193 3516
rect 460155 3485 460167 3488
rect 460109 3479 460167 3485
rect 466181 3485 466193 3488
rect 466227 3485 466239 3519
rect 466181 3479 466239 3485
rect 466270 3476 466276 3528
rect 466328 3516 466334 3528
rect 573818 3516 573824 3528
rect 466328 3488 573824 3516
rect 466328 3476 466334 3488
rect 573818 3476 573824 3488
rect 573876 3476 573882 3528
rect 368072 3420 376800 3448
rect 368072 3408 368078 3420
rect 382366 3408 382372 3460
rect 382424 3448 382430 3460
rect 386598 3448 386604 3460
rect 382424 3420 386604 3448
rect 382424 3408 382430 3420
rect 386598 3408 386604 3420
rect 386656 3408 386662 3460
rect 403618 3408 403624 3460
rect 403676 3448 403682 3460
rect 407298 3448 407304 3460
rect 403676 3420 407304 3448
rect 403676 3408 403682 3420
rect 407298 3408 407304 3420
rect 407356 3408 407362 3460
rect 422754 3448 422760 3460
rect 407408 3420 422760 3448
rect 29086 3340 29092 3392
rect 29144 3380 29150 3392
rect 35158 3380 35164 3392
rect 29144 3352 35164 3380
rect 29144 3340 29150 3352
rect 35158 3340 35164 3352
rect 35216 3340 35222 3392
rect 36170 3340 36176 3392
rect 36228 3380 36234 3392
rect 39298 3380 39304 3392
rect 36228 3352 39304 3380
rect 36228 3340 36234 3352
rect 39298 3340 39304 3352
rect 39356 3340 39362 3392
rect 45465 3383 45523 3389
rect 45465 3349 45477 3383
rect 45511 3380 45523 3383
rect 45511 3352 58296 3380
rect 45511 3349 45523 3352
rect 45465 3343 45523 3349
rect 10042 3272 10048 3324
rect 10100 3312 10106 3324
rect 13078 3312 13084 3324
rect 10100 3284 13084 3312
rect 10100 3272 10106 3284
rect 13078 3272 13084 3284
rect 13136 3272 13142 3324
rect 42150 3272 42156 3324
rect 42208 3312 42214 3324
rect 57238 3312 57244 3324
rect 42208 3284 57244 3312
rect 42208 3272 42214 3284
rect 57238 3272 57244 3284
rect 57296 3272 57302 3324
rect 58268 3312 58296 3352
rect 59998 3340 60004 3392
rect 60056 3380 60062 3392
rect 60642 3380 60648 3392
rect 60056 3352 60648 3380
rect 60056 3340 60062 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 63586 3340 63592 3392
rect 63644 3380 63650 3392
rect 64782 3380 64788 3392
rect 63644 3352 64788 3380
rect 63644 3340 63650 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 70670 3340 70676 3392
rect 70728 3380 70734 3392
rect 71682 3380 71688 3392
rect 70728 3352 71688 3380
rect 70728 3340 70734 3352
rect 71682 3340 71688 3352
rect 71740 3340 71746 3392
rect 251818 3380 251824 3392
rect 71792 3352 251824 3380
rect 61378 3312 61384 3324
rect 58268 3284 61384 3312
rect 61378 3272 61384 3284
rect 61436 3272 61442 3324
rect 52822 3204 52828 3256
rect 52880 3244 52886 3256
rect 53742 3244 53748 3256
rect 52880 3216 53748 3244
rect 52880 3204 52886 3216
rect 53742 3204 53748 3216
rect 53800 3204 53806 3256
rect 54018 3204 54024 3256
rect 54076 3244 54082 3256
rect 54076 3216 59676 3244
rect 54076 3204 54082 3216
rect 43346 3136 43352 3188
rect 43404 3176 43410 3188
rect 45465 3179 45523 3185
rect 45465 3176 45477 3179
rect 43404 3148 45477 3176
rect 43404 3136 43410 3148
rect 45465 3145 45477 3148
rect 45511 3145 45523 3179
rect 45465 3139 45523 3145
rect 59648 3108 59676 3216
rect 64782 3204 64788 3256
rect 64840 3244 64846 3256
rect 71792 3244 71820 3352
rect 251818 3340 251824 3352
rect 251876 3340 251882 3392
rect 282825 3383 282883 3389
rect 282825 3349 282837 3383
rect 282871 3380 282883 3383
rect 289814 3380 289820 3392
rect 282871 3352 289820 3380
rect 282871 3349 282883 3352
rect 282825 3343 282883 3349
rect 289814 3340 289820 3352
rect 289872 3340 289878 3392
rect 299106 3340 299112 3392
rect 299164 3380 299170 3392
rect 302878 3380 302884 3392
rect 299164 3352 302884 3380
rect 299164 3340 299170 3352
rect 302878 3340 302884 3352
rect 302936 3340 302942 3392
rect 310974 3340 310980 3392
rect 311032 3380 311038 3392
rect 311032 3352 341104 3380
rect 311032 3340 311038 3352
rect 71866 3272 71872 3324
rect 71924 3312 71930 3324
rect 253198 3312 253204 3324
rect 71924 3284 253204 3312
rect 71924 3272 71930 3284
rect 253198 3272 253204 3284
rect 253256 3272 253262 3324
rect 288434 3312 288440 3324
rect 276400 3284 288440 3312
rect 64840 3216 71820 3244
rect 71884 3216 74580 3244
rect 64840 3204 64846 3216
rect 61194 3136 61200 3188
rect 61252 3176 61258 3188
rect 61252 3148 67956 3176
rect 61252 3136 61258 3148
rect 66898 3108 66904 3120
rect 59648 3080 66904 3108
rect 66898 3068 66904 3080
rect 66956 3068 66962 3120
rect 67928 3108 67956 3148
rect 68278 3136 68284 3188
rect 68336 3176 68342 3188
rect 71884 3176 71912 3216
rect 68336 3148 71912 3176
rect 68336 3136 68342 3148
rect 71038 3108 71044 3120
rect 67928 3080 71044 3108
rect 71038 3068 71044 3080
rect 71096 3068 71102 3120
rect 74552 3040 74580 3216
rect 77846 3204 77852 3256
rect 77904 3244 77910 3256
rect 78582 3244 78588 3256
rect 77904 3216 78588 3244
rect 77904 3204 77910 3216
rect 78582 3204 78588 3216
rect 78640 3204 78646 3256
rect 81434 3204 81440 3256
rect 81492 3244 81498 3256
rect 82722 3244 82728 3256
rect 81492 3216 82728 3244
rect 81492 3204 81498 3216
rect 82722 3204 82728 3216
rect 82780 3204 82786 3256
rect 84838 3244 84844 3256
rect 82832 3216 84844 3244
rect 75454 3136 75460 3188
rect 75512 3176 75518 3188
rect 79318 3176 79324 3188
rect 75512 3148 79324 3176
rect 75512 3136 75518 3148
rect 79318 3136 79324 3148
rect 79376 3136 79382 3188
rect 82630 3136 82636 3188
rect 82688 3176 82694 3188
rect 82832 3176 82860 3216
rect 84838 3204 84844 3216
rect 84896 3204 84902 3256
rect 84930 3204 84936 3256
rect 84988 3244 84994 3256
rect 85482 3244 85488 3256
rect 84988 3216 85488 3244
rect 84988 3204 84994 3216
rect 85482 3204 85488 3216
rect 85540 3204 85546 3256
rect 88518 3204 88524 3256
rect 88576 3244 88582 3256
rect 89622 3244 89628 3256
rect 88576 3216 89628 3244
rect 88576 3204 88582 3216
rect 89622 3204 89628 3216
rect 89680 3204 89686 3256
rect 254578 3244 254584 3256
rect 89732 3216 254584 3244
rect 82688 3148 82860 3176
rect 82909 3179 82967 3185
rect 82688 3136 82694 3148
rect 82909 3145 82921 3179
rect 82955 3176 82967 3179
rect 89732 3176 89760 3216
rect 254578 3204 254584 3216
rect 254636 3204 254642 3256
rect 269298 3204 269304 3256
rect 269356 3244 269362 3256
rect 273257 3247 273315 3253
rect 273257 3244 273269 3247
rect 269356 3216 273269 3244
rect 269356 3204 269362 3216
rect 273257 3213 273269 3216
rect 273303 3213 273315 3247
rect 273257 3207 273315 3213
rect 255958 3176 255964 3188
rect 82955 3148 89760 3176
rect 94424 3148 255964 3176
rect 82955 3145 82967 3148
rect 82909 3139 82967 3145
rect 89714 3068 89720 3120
rect 89772 3108 89778 3120
rect 94424 3108 94452 3148
rect 255958 3136 255964 3148
rect 256016 3136 256022 3188
rect 272886 3136 272892 3188
rect 272944 3176 272950 3188
rect 276400 3176 276428 3284
rect 288434 3272 288440 3284
rect 288492 3272 288498 3324
rect 303798 3272 303804 3324
rect 303856 3312 303862 3324
rect 336185 3315 336243 3321
rect 336185 3312 336197 3315
rect 303856 3284 336197 3312
rect 303856 3272 303862 3284
rect 336185 3281 336197 3284
rect 336231 3281 336243 3315
rect 336185 3275 336243 3281
rect 339494 3272 339500 3324
rect 339552 3312 339558 3324
rect 340782 3312 340788 3324
rect 339552 3284 340788 3312
rect 339552 3272 339558 3284
rect 340782 3272 340788 3284
rect 340840 3272 340846 3324
rect 341076 3312 341104 3352
rect 341150 3340 341156 3392
rect 341208 3380 341214 3392
rect 349157 3383 349215 3389
rect 349157 3380 349169 3383
rect 341208 3352 349169 3380
rect 341208 3340 341214 3352
rect 349157 3349 349169 3352
rect 349203 3349 349215 3383
rect 349157 3343 349215 3349
rect 350534 3340 350540 3392
rect 350592 3380 350598 3392
rect 353662 3380 353668 3392
rect 350592 3352 353668 3380
rect 350592 3340 350598 3352
rect 353662 3340 353668 3352
rect 353720 3340 353726 3392
rect 353754 3340 353760 3392
rect 353812 3380 353818 3392
rect 375650 3380 375656 3392
rect 353812 3352 375656 3380
rect 353812 3340 353818 3352
rect 375650 3340 375656 3352
rect 375708 3340 375714 3392
rect 376680 3352 376800 3380
rect 345845 3315 345903 3321
rect 341076 3284 345796 3312
rect 276474 3204 276480 3256
rect 276532 3244 276538 3256
rect 288526 3244 288532 3256
rect 276532 3216 288532 3244
rect 276532 3204 276538 3216
rect 288526 3204 288532 3216
rect 288584 3204 288590 3256
rect 291930 3204 291936 3256
rect 291988 3244 291994 3256
rect 316678 3244 316684 3256
rect 291988 3216 316684 3244
rect 291988 3204 291994 3216
rect 316678 3204 316684 3216
rect 316736 3204 316742 3256
rect 318058 3204 318064 3256
rect 318116 3244 318122 3256
rect 345661 3247 345719 3253
rect 345661 3244 345673 3247
rect 318116 3216 345673 3244
rect 318116 3204 318122 3216
rect 345661 3213 345673 3216
rect 345707 3213 345719 3247
rect 345768 3244 345796 3284
rect 345845 3281 345857 3315
rect 345891 3312 345903 3315
rect 348418 3312 348424 3324
rect 345891 3284 348424 3312
rect 345891 3281 345903 3284
rect 345845 3275 345903 3281
rect 348418 3272 348424 3284
rect 348476 3272 348482 3324
rect 348970 3272 348976 3324
rect 349028 3312 349034 3324
rect 362037 3315 362095 3321
rect 362037 3312 362049 3315
rect 349028 3284 362049 3312
rect 349028 3272 349034 3284
rect 362037 3281 362049 3284
rect 362083 3281 362095 3315
rect 362037 3275 362095 3281
rect 362126 3272 362132 3324
rect 362184 3312 362190 3324
rect 362862 3312 362868 3324
rect 362184 3284 362868 3312
rect 362184 3272 362190 3284
rect 362862 3272 362868 3284
rect 362920 3272 362926 3324
rect 364518 3272 364524 3324
rect 364576 3312 364582 3324
rect 376680 3312 376708 3352
rect 376772 3321 376800 3352
rect 404262 3340 404268 3392
rect 404320 3380 404326 3392
rect 407408 3380 407436 3420
rect 422754 3408 422760 3420
rect 422812 3408 422818 3460
rect 424318 3408 424324 3460
rect 424376 3448 424382 3460
rect 425146 3448 425152 3460
rect 424376 3420 425152 3448
rect 424376 3408 424382 3420
rect 425146 3408 425152 3420
rect 425204 3408 425210 3460
rect 425241 3451 425299 3457
rect 425241 3417 425253 3451
rect 425287 3448 425299 3451
rect 467926 3448 467932 3460
rect 425287 3420 467932 3448
rect 425287 3417 425299 3420
rect 425241 3411 425299 3417
rect 467926 3408 467932 3420
rect 467984 3408 467990 3460
rect 469030 3408 469036 3460
rect 469088 3448 469094 3460
rect 578602 3448 578608 3460
rect 469088 3420 578608 3448
rect 469088 3408 469094 3420
rect 578602 3408 578608 3420
rect 578660 3408 578666 3460
rect 404320 3352 407436 3380
rect 404320 3340 404326 3352
rect 409782 3340 409788 3392
rect 409840 3380 409846 3392
rect 433889 3383 433947 3389
rect 433889 3380 433901 3383
rect 409840 3352 433901 3380
rect 409840 3340 409846 3352
rect 433889 3349 433901 3352
rect 433935 3349 433947 3383
rect 433889 3343 433947 3349
rect 433978 3340 433984 3392
rect 434036 3380 434042 3392
rect 435818 3380 435824 3392
rect 434036 3352 435824 3380
rect 434036 3340 434042 3352
rect 435818 3340 435824 3352
rect 435876 3340 435882 3392
rect 438118 3340 438124 3392
rect 438176 3380 438182 3392
rect 446401 3383 446459 3389
rect 446401 3380 446413 3383
rect 438176 3352 446413 3380
rect 438176 3340 438182 3352
rect 446401 3349 446413 3352
rect 446447 3349 446459 3383
rect 446401 3343 446459 3349
rect 446493 3383 446551 3389
rect 446493 3349 446505 3383
rect 446539 3380 446551 3383
rect 446539 3352 510108 3380
rect 446539 3349 446551 3352
rect 446493 3343 446551 3349
rect 364576 3284 376708 3312
rect 376757 3315 376815 3321
rect 364576 3272 364582 3284
rect 376757 3281 376769 3315
rect 376803 3281 376815 3315
rect 376757 3275 376815 3281
rect 394510 3272 394516 3324
rect 394568 3312 394574 3324
rect 400214 3312 400220 3324
rect 394568 3284 400220 3312
rect 394568 3272 394574 3284
rect 400214 3272 400220 3284
rect 400272 3272 400278 3324
rect 404998 3272 405004 3324
rect 405056 3312 405062 3324
rect 416866 3312 416872 3324
rect 405056 3284 416872 3312
rect 405056 3272 405062 3284
rect 416866 3272 416872 3284
rect 416924 3272 416930 3324
rect 420178 3272 420184 3324
rect 420236 3312 420242 3324
rect 446582 3312 446588 3324
rect 420236 3284 446588 3312
rect 420236 3272 420242 3284
rect 446582 3272 446588 3284
rect 446640 3272 446646 3324
rect 446677 3315 446735 3321
rect 446677 3281 446689 3315
rect 446723 3312 446735 3315
rect 503622 3312 503628 3324
rect 446723 3284 503628 3312
rect 446723 3281 446735 3284
rect 446677 3275 446735 3281
rect 503622 3272 503628 3284
rect 503680 3272 503686 3324
rect 510080 3312 510108 3352
rect 514018 3340 514024 3392
rect 514076 3380 514082 3392
rect 517882 3380 517888 3392
rect 514076 3352 517888 3380
rect 514076 3340 514082 3352
rect 517882 3340 517888 3352
rect 517940 3340 517946 3392
rect 525058 3380 525064 3392
rect 517992 3352 525064 3380
rect 514386 3312 514392 3324
rect 510080 3284 514392 3312
rect 514386 3272 514392 3284
rect 514444 3272 514450 3324
rect 516870 3272 516876 3324
rect 516928 3312 516934 3324
rect 517992 3312 518020 3352
rect 525058 3340 525064 3352
rect 525116 3340 525122 3392
rect 527818 3340 527824 3392
rect 527876 3380 527882 3392
rect 567838 3380 567844 3392
rect 527876 3352 567844 3380
rect 527876 3340 527882 3352
rect 567838 3340 567844 3352
rect 567896 3340 567902 3392
rect 577406 3312 577412 3324
rect 516928 3284 518020 3312
rect 518084 3284 577412 3312
rect 516928 3272 516934 3284
rect 350169 3247 350227 3253
rect 350169 3244 350181 3247
rect 345768 3216 350181 3244
rect 345661 3207 345719 3213
rect 350169 3213 350181 3216
rect 350215 3213 350227 3247
rect 350169 3207 350227 3213
rect 350258 3204 350264 3256
rect 350316 3244 350322 3256
rect 354309 3247 354367 3253
rect 354309 3244 354321 3247
rect 350316 3216 354321 3244
rect 350316 3204 350322 3216
rect 354309 3213 354321 3216
rect 354355 3213 354367 3247
rect 354309 3207 354367 3213
rect 354401 3247 354459 3253
rect 354401 3213 354413 3247
rect 354447 3244 354459 3247
rect 357250 3244 357256 3256
rect 354447 3216 357256 3244
rect 354447 3213 354459 3216
rect 354401 3207 354459 3213
rect 357250 3204 357256 3216
rect 357308 3204 357314 3256
rect 357342 3204 357348 3256
rect 357400 3244 357406 3256
rect 376018 3244 376024 3256
rect 357400 3216 376024 3244
rect 357400 3204 357406 3216
rect 376018 3204 376024 3216
rect 376076 3204 376082 3256
rect 409138 3204 409144 3256
rect 409196 3244 409202 3256
rect 432322 3244 432328 3256
rect 409196 3216 432328 3244
rect 409196 3204 409202 3216
rect 432322 3204 432328 3216
rect 432380 3204 432386 3256
rect 433889 3247 433947 3253
rect 433889 3213 433901 3247
rect 433935 3244 433947 3247
rect 437014 3244 437020 3256
rect 433935 3216 437020 3244
rect 433935 3213 433947 3216
rect 433889 3207 433947 3213
rect 437014 3204 437020 3216
rect 437072 3204 437078 3256
rect 441617 3247 441675 3253
rect 441617 3213 441629 3247
rect 441663 3244 441675 3247
rect 446214 3244 446220 3256
rect 441663 3216 446220 3244
rect 441663 3213 441675 3216
rect 441617 3207 441675 3213
rect 446214 3204 446220 3216
rect 446272 3204 446278 3256
rect 446309 3247 446367 3253
rect 446309 3213 446321 3247
rect 446355 3244 446367 3247
rect 496538 3244 496544 3256
rect 446355 3216 496544 3244
rect 446355 3213 446367 3216
rect 446309 3207 446367 3213
rect 496538 3204 496544 3216
rect 496596 3204 496602 3256
rect 512638 3204 512644 3256
rect 512696 3244 512702 3256
rect 518084 3244 518112 3284
rect 577406 3272 577412 3284
rect 577464 3272 577470 3324
rect 512696 3216 518112 3244
rect 518161 3247 518219 3253
rect 512696 3204 512702 3216
rect 518161 3213 518173 3247
rect 518207 3244 518219 3247
rect 570230 3244 570236 3256
rect 518207 3216 570236 3244
rect 518207 3213 518219 3216
rect 518161 3207 518219 3213
rect 570230 3204 570236 3216
rect 570288 3204 570294 3256
rect 290458 3176 290464 3188
rect 272944 3148 276428 3176
rect 278240 3148 290464 3176
rect 272944 3136 272950 3148
rect 89772 3080 94452 3108
rect 89772 3068 89778 3080
rect 94498 3068 94504 3120
rect 94556 3108 94562 3120
rect 95142 3108 95148 3120
rect 94556 3080 95148 3108
rect 94556 3068 94562 3080
rect 95142 3068 95148 3080
rect 95200 3068 95206 3120
rect 95694 3068 95700 3120
rect 95752 3108 95758 3120
rect 96522 3108 96528 3120
rect 95752 3080 96528 3108
rect 95752 3068 95758 3080
rect 96522 3068 96528 3080
rect 96580 3068 96586 3120
rect 98086 3068 98092 3120
rect 98144 3108 98150 3120
rect 99190 3108 99196 3120
rect 98144 3080 99196 3108
rect 98144 3068 98150 3080
rect 99190 3068 99196 3080
rect 99248 3068 99254 3120
rect 101582 3068 101588 3120
rect 101640 3108 101646 3120
rect 102042 3108 102048 3120
rect 101640 3080 102048 3108
rect 101640 3068 101646 3080
rect 102042 3068 102048 3080
rect 102100 3068 102106 3120
rect 102778 3068 102784 3120
rect 102836 3108 102842 3120
rect 103422 3108 103428 3120
rect 102836 3080 103428 3108
rect 102836 3068 102842 3080
rect 103422 3068 103428 3080
rect 103480 3068 103486 3120
rect 105170 3068 105176 3120
rect 105228 3108 105234 3120
rect 106182 3108 106188 3120
rect 105228 3080 106188 3108
rect 105228 3068 105234 3080
rect 106182 3068 106188 3080
rect 106240 3068 106246 3120
rect 106366 3068 106372 3120
rect 106424 3108 106430 3120
rect 107470 3108 107476 3120
rect 106424 3080 107476 3108
rect 106424 3068 106430 3080
rect 107470 3068 107476 3080
rect 107528 3068 107534 3120
rect 257338 3108 257344 3120
rect 108316 3080 257344 3108
rect 77938 3040 77944 3052
rect 74552 3012 77944 3040
rect 77938 3000 77944 3012
rect 77996 3000 78002 3052
rect 93302 3000 93308 3052
rect 93360 3040 93366 3052
rect 102594 3040 102600 3052
rect 93360 3012 102600 3040
rect 93360 3000 93366 3012
rect 102594 3000 102600 3012
rect 102652 3000 102658 3052
rect 79042 2932 79048 2984
rect 79100 2972 79106 2984
rect 82909 2975 82967 2981
rect 82909 2972 82921 2975
rect 79100 2944 82921 2972
rect 79100 2932 79106 2944
rect 82909 2941 82921 2944
rect 82955 2941 82967 2975
rect 82909 2935 82967 2941
rect 86126 2932 86132 2984
rect 86184 2972 86190 2984
rect 93857 2975 93915 2981
rect 93857 2972 93869 2975
rect 86184 2944 93869 2972
rect 86184 2932 86190 2944
rect 93857 2941 93869 2944
rect 93903 2941 93915 2975
rect 93857 2935 93915 2941
rect 96890 2932 96896 2984
rect 96948 2972 96954 2984
rect 108316 2972 108344 3080
rect 257338 3068 257344 3080
rect 257396 3068 257402 3120
rect 277670 3068 277676 3120
rect 277728 3108 277734 3120
rect 278240 3108 278268 3148
rect 290458 3136 290464 3148
rect 290516 3136 290522 3188
rect 295518 3136 295524 3188
rect 295576 3176 295582 3188
rect 319438 3176 319444 3188
rect 295576 3148 319444 3176
rect 295576 3136 295582 3148
rect 319438 3136 319444 3148
rect 319496 3136 319502 3188
rect 325234 3136 325240 3188
rect 325292 3176 325298 3188
rect 350534 3176 350540 3188
rect 325292 3148 350540 3176
rect 325292 3136 325298 3148
rect 350534 3136 350540 3148
rect 350592 3136 350598 3188
rect 350626 3136 350632 3188
rect 350684 3176 350690 3188
rect 358906 3176 358912 3188
rect 350684 3148 358912 3176
rect 350684 3136 350690 3148
rect 358906 3136 358912 3148
rect 358964 3136 358970 3188
rect 363693 3179 363751 3185
rect 363693 3145 363705 3179
rect 363739 3176 363751 3179
rect 367278 3176 367284 3188
rect 363739 3148 367284 3176
rect 363739 3145 363751 3148
rect 363693 3139 363751 3145
rect 367278 3136 367284 3148
rect 367336 3136 367342 3188
rect 407022 3136 407028 3188
rect 407080 3176 407086 3188
rect 429930 3176 429936 3188
rect 407080 3148 429936 3176
rect 407080 3136 407086 3148
rect 429930 3136 429936 3148
rect 429988 3136 429994 3188
rect 431218 3136 431224 3188
rect 431276 3176 431282 3188
rect 431276 3148 477632 3176
rect 431276 3136 431282 3148
rect 277728 3080 278268 3108
rect 277728 3068 277734 3080
rect 278866 3068 278872 3120
rect 278924 3108 278930 3120
rect 287609 3111 287667 3117
rect 287609 3108 287621 3111
rect 278924 3080 287621 3108
rect 278924 3068 278930 3080
rect 287609 3077 287621 3080
rect 287655 3077 287667 3111
rect 287609 3071 287667 3077
rect 309778 3068 309784 3120
rect 309836 3108 309842 3120
rect 335541 3111 335599 3117
rect 335541 3108 335553 3111
rect 309836 3080 335553 3108
rect 309836 3068 309842 3080
rect 335541 3077 335553 3080
rect 335587 3077 335599 3111
rect 345658 3108 345664 3120
rect 335541 3071 335599 3077
rect 336016 3080 345664 3108
rect 258810 3040 258816 3052
rect 96948 2944 108344 2972
rect 108408 3012 258816 3040
rect 96948 2932 96954 2944
rect 103974 2864 103980 2916
rect 104032 2904 104038 2916
rect 108408 2904 108436 3012
rect 258810 3000 258816 3012
rect 258868 3000 258874 3052
rect 273257 3043 273315 3049
rect 273257 3009 273269 3043
rect 273303 3040 273315 3043
rect 282825 3043 282883 3049
rect 282825 3040 282837 3043
rect 273303 3012 282837 3040
rect 273303 3009 273315 3012
rect 273257 3003 273315 3009
rect 282825 3009 282837 3012
rect 282871 3009 282883 3043
rect 282825 3003 282883 3009
rect 293126 3000 293132 3052
rect 293184 3040 293190 3052
rect 312538 3040 312544 3052
rect 293184 3012 312544 3040
rect 293184 3000 293190 3012
rect 312538 3000 312544 3012
rect 312596 3000 312602 3052
rect 315758 3000 315764 3052
rect 315816 3040 315822 3052
rect 324222 3040 324228 3052
rect 315816 3012 324228 3040
rect 315816 3000 315822 3012
rect 324222 3000 324228 3012
rect 324280 3000 324286 3052
rect 326341 3043 326399 3049
rect 326341 3009 326353 3043
rect 326387 3040 326399 3043
rect 335906 3040 335912 3052
rect 326387 3012 335912 3040
rect 326387 3009 326399 3012
rect 326341 3003 326399 3009
rect 335906 3000 335912 3012
rect 335964 3000 335970 3052
rect 112346 2932 112352 2984
rect 112404 2972 112410 2984
rect 113082 2972 113088 2984
rect 112404 2944 113088 2972
rect 112404 2932 112410 2944
rect 113082 2932 113088 2944
rect 113140 2932 113146 2984
rect 113542 2932 113548 2984
rect 113600 2972 113606 2984
rect 114462 2972 114468 2984
rect 113600 2944 114468 2972
rect 113600 2932 113606 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 115934 2932 115940 2984
rect 115992 2972 115998 2984
rect 116946 2972 116952 2984
rect 115992 2944 116952 2972
rect 115992 2932 115998 2944
rect 116946 2932 116952 2944
rect 117004 2932 117010 2984
rect 119430 2932 119436 2984
rect 119488 2972 119494 2984
rect 119982 2972 119988 2984
rect 119488 2944 119988 2972
rect 119488 2932 119494 2944
rect 119982 2932 119988 2944
rect 120040 2932 120046 2984
rect 120626 2932 120632 2984
rect 120684 2972 120690 2984
rect 121362 2972 121368 2984
rect 120684 2944 121368 2972
rect 120684 2932 120690 2944
rect 121362 2932 121368 2944
rect 121420 2932 121426 2984
rect 258718 2972 258724 2984
rect 121472 2944 258724 2972
rect 104032 2876 108436 2904
rect 104032 2864 104038 2876
rect 111150 2864 111156 2916
rect 111208 2904 111214 2916
rect 121472 2904 121500 2944
rect 258718 2932 258724 2944
rect 258776 2932 258782 2984
rect 316954 2932 316960 2984
rect 317012 2972 317018 2984
rect 336016 2972 336044 3080
rect 345658 3068 345664 3080
rect 345716 3068 345722 3120
rect 346670 3068 346676 3120
rect 346728 3108 346734 3120
rect 370498 3108 370504 3120
rect 346728 3080 370504 3108
rect 346728 3068 346734 3080
rect 370498 3068 370504 3080
rect 370556 3068 370562 3120
rect 405642 3068 405648 3120
rect 405700 3108 405706 3120
rect 426342 3108 426348 3120
rect 405700 3080 426348 3108
rect 405700 3068 405706 3080
rect 426342 3068 426348 3080
rect 426400 3068 426406 3120
rect 428458 3068 428464 3120
rect 428516 3108 428522 3120
rect 475102 3108 475108 3120
rect 428516 3080 475108 3108
rect 428516 3068 428522 3080
rect 475102 3068 475108 3080
rect 475160 3068 475166 3120
rect 475378 3068 475384 3120
rect 475436 3108 475442 3120
rect 477494 3108 477500 3120
rect 475436 3080 477500 3108
rect 475436 3068 475442 3080
rect 477494 3068 477500 3080
rect 477552 3068 477558 3120
rect 477604 3108 477632 3148
rect 505738 3136 505744 3188
rect 505796 3176 505802 3188
rect 563146 3176 563152 3188
rect 505796 3148 563152 3176
rect 505796 3136 505802 3148
rect 563146 3136 563152 3148
rect 563204 3136 563210 3188
rect 482278 3108 482284 3120
rect 477604 3080 482284 3108
rect 482278 3068 482284 3080
rect 482336 3068 482342 3120
rect 524966 3068 524972 3120
rect 525024 3108 525030 3120
rect 560754 3108 560760 3120
rect 525024 3080 560760 3108
rect 525024 3068 525030 3080
rect 560754 3068 560760 3080
rect 560812 3068 560818 3120
rect 336090 3000 336096 3052
rect 336148 3040 336154 3052
rect 363693 3043 363751 3049
rect 363693 3040 363705 3043
rect 336148 3012 363705 3040
rect 336148 3000 336154 3012
rect 363693 3009 363705 3012
rect 363739 3009 363751 3043
rect 363693 3003 363751 3009
rect 395890 3000 395896 3052
rect 395948 3040 395954 3052
rect 401318 3040 401324 3052
rect 395948 3012 401324 3040
rect 395948 3000 395954 3012
rect 401318 3000 401324 3012
rect 401376 3000 401382 3052
rect 406378 3000 406384 3052
rect 406436 3040 406442 3052
rect 410886 3040 410892 3052
rect 406436 3012 410892 3040
rect 406436 3000 406442 3012
rect 410886 3000 410892 3012
rect 410944 3000 410950 3052
rect 416590 3000 416596 3052
rect 416648 3040 416654 3052
rect 431221 3043 431279 3049
rect 431221 3040 431233 3043
rect 416648 3012 431233 3040
rect 416648 3000 416654 3012
rect 431221 3009 431233 3012
rect 431267 3009 431279 3043
rect 431221 3003 431279 3009
rect 431310 3000 431316 3052
rect 431368 3040 431374 3052
rect 459646 3040 459652 3052
rect 431368 3012 459652 3040
rect 431368 3000 431374 3012
rect 459646 3000 459652 3012
rect 459704 3000 459710 3052
rect 461581 3043 461639 3049
rect 461581 3009 461593 3043
rect 461627 3040 461639 3043
rect 489362 3040 489368 3052
rect 461627 3012 489368 3040
rect 461627 3009 461639 3012
rect 461581 3003 461639 3009
rect 489362 3000 489368 3012
rect 489420 3000 489426 3052
rect 509878 3000 509884 3052
rect 509936 3040 509942 3052
rect 518161 3043 518219 3049
rect 518161 3040 518173 3043
rect 509936 3012 518173 3040
rect 509936 3000 509942 3012
rect 518161 3009 518173 3012
rect 518207 3009 518219 3043
rect 518161 3003 518219 3009
rect 523678 3000 523684 3052
rect 523736 3040 523742 3052
rect 553578 3040 553584 3052
rect 523736 3012 553584 3040
rect 523736 3000 523742 3012
rect 553578 3000 553584 3012
rect 553636 3000 553642 3052
rect 317012 2944 336044 2972
rect 336185 2975 336243 2981
rect 317012 2932 317018 2944
rect 336185 2941 336197 2975
rect 336231 2972 336243 2975
rect 344370 2972 344376 2984
rect 336231 2944 344376 2972
rect 336231 2941 336243 2944
rect 336185 2935 336243 2941
rect 344370 2932 344376 2944
rect 344428 2932 344434 2984
rect 345474 2932 345480 2984
rect 345532 2972 345538 2984
rect 351178 2972 351184 2984
rect 345532 2944 351184 2972
rect 345532 2932 345538 2944
rect 351178 2932 351184 2944
rect 351236 2932 351242 2984
rect 354401 2975 354459 2981
rect 354401 2972 354413 2975
rect 352484 2944 354413 2972
rect 260098 2904 260104 2916
rect 111208 2876 121500 2904
rect 121564 2876 260104 2904
rect 111208 2864 111214 2876
rect 93857 2839 93915 2845
rect 93857 2805 93869 2839
rect 93903 2836 93915 2839
rect 95878 2836 95884 2848
rect 93903 2808 95884 2836
rect 93903 2805 93915 2808
rect 93857 2799 93915 2805
rect 95878 2796 95884 2808
rect 95936 2796 95942 2848
rect 114738 2796 114744 2848
rect 114796 2836 114802 2848
rect 121564 2836 121592 2876
rect 260098 2864 260104 2876
rect 260156 2864 260162 2916
rect 275278 2864 275284 2916
rect 275336 2904 275342 2916
rect 275922 2904 275928 2916
rect 275336 2876 275928 2904
rect 275336 2864 275342 2876
rect 275922 2864 275928 2876
rect 275980 2864 275986 2916
rect 319254 2864 319260 2916
rect 319312 2904 319318 2916
rect 322753 2907 322811 2913
rect 322753 2904 322765 2907
rect 319312 2876 322765 2904
rect 319312 2864 319318 2876
rect 322753 2873 322765 2876
rect 322799 2873 322811 2907
rect 322753 2867 322811 2873
rect 322842 2864 322848 2916
rect 322900 2904 322906 2916
rect 327074 2904 327080 2916
rect 322900 2876 327080 2904
rect 322900 2864 322906 2876
rect 327074 2864 327080 2876
rect 327132 2864 327138 2916
rect 335464 2876 344324 2904
rect 114796 2808 121592 2836
rect 114796 2796 114802 2808
rect 121822 2796 121828 2848
rect 121880 2836 121886 2848
rect 261478 2836 261484 2848
rect 121880 2808 261484 2836
rect 121880 2796 121886 2808
rect 261478 2796 261484 2808
rect 261536 2796 261542 2848
rect 330018 2796 330024 2848
rect 330076 2836 330082 2848
rect 335464 2836 335492 2876
rect 330076 2808 335492 2836
rect 335541 2839 335599 2845
rect 330076 2796 330082 2808
rect 335541 2805 335553 2839
rect 335587 2836 335599 2839
rect 339865 2839 339923 2845
rect 339865 2836 339877 2839
rect 335587 2808 339877 2836
rect 335587 2805 335599 2808
rect 335541 2799 335599 2805
rect 339865 2805 339877 2808
rect 339911 2805 339923 2839
rect 343634 2836 343640 2848
rect 339865 2799 339923 2805
rect 340340 2808 343640 2836
rect 339957 2771 340015 2777
rect 339957 2737 339969 2771
rect 340003 2768 340015 2771
rect 340340 2768 340368 2808
rect 343634 2796 343640 2808
rect 343692 2796 343698 2848
rect 344296 2836 344324 2876
rect 344554 2864 344560 2916
rect 344612 2904 344618 2916
rect 352484 2904 352512 2944
rect 354401 2941 354413 2944
rect 354447 2941 354459 2975
rect 354401 2935 354459 2941
rect 354950 2932 354956 2984
rect 355008 2972 355014 2984
rect 355962 2972 355968 2984
rect 355008 2944 355968 2972
rect 355008 2932 355014 2944
rect 355962 2932 355968 2944
rect 356020 2932 356026 2984
rect 356054 2932 356060 2984
rect 356112 2972 356118 2984
rect 356698 2972 356704 2984
rect 356112 2944 356704 2972
rect 356112 2932 356118 2944
rect 356698 2932 356704 2944
rect 356756 2932 356762 2984
rect 356790 2932 356796 2984
rect 356848 2972 356854 2984
rect 359458 2972 359464 2984
rect 356848 2944 359464 2972
rect 356848 2932 356854 2944
rect 359458 2932 359464 2944
rect 359516 2932 359522 2984
rect 359553 2975 359611 2981
rect 359553 2941 359565 2975
rect 359599 2972 359611 2975
rect 374362 2972 374368 2984
rect 359599 2944 374368 2972
rect 359599 2941 359611 2944
rect 359553 2935 359611 2941
rect 374362 2932 374368 2944
rect 374420 2932 374426 2984
rect 395982 2932 395988 2984
rect 396040 2972 396046 2984
rect 402514 2972 402520 2984
rect 396040 2944 402520 2972
rect 396040 2932 396046 2944
rect 402514 2932 402520 2944
rect 402572 2932 402578 2984
rect 417418 2932 417424 2984
rect 417476 2972 417482 2984
rect 428734 2972 428740 2984
rect 417476 2944 428740 2972
rect 417476 2932 417482 2944
rect 428734 2932 428740 2944
rect 428792 2932 428798 2984
rect 429838 2932 429844 2984
rect 429896 2972 429902 2984
rect 448974 2972 448980 2984
rect 429896 2944 448980 2972
rect 429896 2932 429902 2944
rect 448974 2932 448980 2944
rect 449032 2932 449038 2984
rect 451829 2975 451887 2981
rect 451829 2972 451841 2975
rect 451292 2944 451841 2972
rect 344612 2876 352512 2904
rect 360749 2907 360807 2913
rect 344612 2864 344618 2876
rect 360749 2873 360761 2907
rect 360795 2904 360807 2907
rect 369765 2907 369823 2913
rect 369765 2904 369777 2907
rect 360795 2876 369777 2904
rect 360795 2873 360807 2876
rect 360749 2867 360807 2873
rect 369765 2873 369777 2876
rect 369811 2873 369823 2907
rect 369765 2867 369823 2873
rect 385862 2864 385868 2916
rect 385920 2904 385926 2916
rect 387058 2904 387064 2916
rect 385920 2876 387064 2904
rect 385920 2864 385926 2876
rect 387058 2864 387064 2876
rect 387116 2864 387122 2916
rect 398190 2864 398196 2916
rect 398248 2904 398254 2916
rect 403710 2904 403716 2916
rect 398248 2876 403716 2904
rect 398248 2864 398254 2876
rect 403710 2864 403716 2876
rect 403768 2864 403774 2916
rect 451185 2907 451243 2913
rect 451185 2904 451197 2907
rect 446324 2876 451197 2904
rect 345569 2839 345627 2845
rect 345569 2836 345581 2839
rect 344296 2808 345581 2836
rect 345569 2805 345581 2808
rect 345615 2805 345627 2839
rect 345569 2799 345627 2805
rect 345661 2839 345719 2845
rect 345661 2805 345673 2839
rect 345707 2836 345719 2839
rect 356054 2836 356060 2848
rect 345707 2808 356060 2836
rect 345707 2805 345719 2808
rect 345661 2799 345719 2805
rect 356054 2796 356060 2808
rect 356112 2796 356118 2848
rect 356146 2796 356152 2848
rect 356204 2836 356210 2848
rect 375834 2836 375840 2848
rect 356204 2808 375840 2836
rect 356204 2796 356210 2808
rect 375834 2796 375840 2808
rect 375892 2796 375898 2848
rect 388438 2836 388444 2848
rect 387076 2808 388444 2836
rect 387076 2780 387104 2808
rect 388438 2796 388444 2808
rect 388496 2796 388502 2848
rect 422297 2839 422355 2845
rect 422297 2805 422309 2839
rect 422343 2836 422355 2839
rect 431865 2839 431923 2845
rect 431865 2836 431877 2839
rect 422343 2808 431877 2836
rect 422343 2805 422355 2808
rect 422297 2799 422355 2805
rect 431865 2805 431877 2808
rect 431911 2805 431923 2839
rect 431865 2799 431923 2805
rect 439590 2796 439596 2848
rect 439648 2836 439654 2848
rect 446324 2836 446352 2876
rect 451185 2873 451197 2876
rect 451231 2873 451243 2907
rect 451185 2867 451243 2873
rect 439648 2808 446352 2836
rect 446401 2839 446459 2845
rect 439648 2796 439654 2808
rect 446401 2805 446413 2839
rect 446447 2836 446459 2839
rect 451292 2836 451320 2944
rect 451829 2941 451841 2944
rect 451875 2941 451887 2975
rect 451829 2935 451887 2941
rect 451921 2975 451979 2981
rect 451921 2941 451933 2975
rect 451967 2972 451979 2975
rect 481082 2972 481088 2984
rect 451967 2944 481088 2972
rect 451967 2941 451979 2944
rect 451921 2935 451979 2941
rect 481082 2932 481088 2944
rect 481140 2932 481146 2984
rect 520918 2932 520924 2984
rect 520976 2972 520982 2984
rect 546494 2972 546500 2984
rect 520976 2944 546500 2972
rect 520976 2932 520982 2944
rect 546494 2932 546500 2944
rect 546552 2932 546558 2984
rect 451369 2907 451427 2913
rect 451369 2873 451381 2907
rect 451415 2904 451427 2907
rect 456797 2907 456855 2913
rect 456797 2904 456809 2907
rect 451415 2876 456809 2904
rect 451415 2873 451427 2876
rect 451369 2867 451427 2873
rect 456797 2873 456809 2876
rect 456843 2873 456855 2907
rect 456797 2867 456855 2873
rect 466365 2907 466423 2913
rect 466365 2873 466377 2907
rect 466411 2904 466423 2907
rect 473906 2904 473912 2916
rect 466411 2876 473912 2904
rect 466411 2873 466423 2876
rect 466365 2867 466423 2873
rect 473906 2864 473912 2876
rect 473964 2864 473970 2916
rect 521010 2864 521016 2916
rect 521068 2904 521074 2916
rect 539318 2904 539324 2916
rect 521068 2876 539324 2904
rect 521068 2864 521074 2876
rect 539318 2864 539324 2876
rect 539376 2864 539382 2916
rect 446447 2808 451320 2836
rect 451829 2839 451887 2845
rect 446447 2805 446459 2808
rect 446401 2799 446459 2805
rect 451829 2805 451841 2839
rect 451875 2836 451887 2839
rect 466822 2836 466828 2848
rect 451875 2808 466828 2836
rect 451875 2805 451887 2808
rect 451829 2799 451887 2805
rect 466822 2796 466828 2808
rect 466880 2796 466886 2848
rect 518158 2796 518164 2848
rect 518216 2836 518222 2848
rect 532234 2836 532240 2848
rect 518216 2808 532240 2836
rect 518216 2796 518222 2808
rect 532234 2796 532240 2808
rect 532292 2796 532298 2848
rect 340003 2740 340368 2768
rect 340003 2737 340015 2740
rect 339957 2731 340015 2737
rect 387058 2728 387064 2780
rect 387116 2728 387122 2780
rect 454681 2771 454739 2777
rect 454681 2737 454693 2771
rect 454727 2768 454739 2771
rect 462038 2768 462044 2780
rect 454727 2740 462044 2768
rect 454727 2737 454739 2740
rect 454681 2731 454739 2737
rect 462038 2728 462044 2740
rect 462096 2728 462102 2780
rect 261018 1232 261024 1284
rect 261076 1272 261082 1284
rect 263873 1275 263931 1281
rect 263873 1272 263885 1275
rect 261076 1244 263885 1272
rect 261076 1232 261082 1244
rect 263873 1241 263885 1244
rect 263919 1241 263931 1275
rect 263873 1235 263931 1241
rect 23106 552 23112 604
rect 23164 592 23170 604
rect 23382 592 23388 604
rect 23164 564 23388 592
rect 23164 552 23170 564
rect 23382 552 23388 564
rect 23440 552 23446 604
rect 164694 552 164700 604
rect 164752 592 164758 604
rect 165522 592 165528 604
rect 164752 564 165528 592
rect 164752 552 164758 564
rect 165522 552 165528 564
rect 165580 552 165586 604
rect 165890 552 165896 604
rect 165948 592 165954 604
rect 166902 592 166908 604
rect 165948 564 166908 592
rect 165948 552 165954 564
rect 166902 552 166908 564
rect 166960 552 166966 604
rect 169386 552 169392 604
rect 169444 592 169450 604
rect 169662 592 169668 604
rect 169444 564 169668 592
rect 169444 552 169450 564
rect 169662 552 169668 564
rect 169720 552 169726 604
rect 182542 552 182548 604
rect 182600 592 182606 604
rect 183462 592 183468 604
rect 182600 564 183468 592
rect 182600 552 182606 564
rect 183462 552 183468 564
rect 183520 552 183526 604
rect 183738 552 183744 604
rect 183796 592 183802 604
rect 184750 592 184756 604
rect 183796 564 184756 592
rect 183796 552 183802 564
rect 184750 552 184756 564
rect 184808 552 184814 604
rect 187234 552 187240 604
rect 187292 592 187298 604
rect 187602 592 187608 604
rect 187292 564 187608 592
rect 187292 552 187298 564
rect 187602 552 187608 564
rect 187660 552 187666 604
rect 189626 552 189632 604
rect 189684 592 189690 604
rect 190362 592 190368 604
rect 189684 564 190368 592
rect 189684 552 189690 564
rect 190362 552 190368 564
rect 190420 552 190426 604
rect 281258 552 281264 604
rect 281316 592 281322 604
rect 281442 592 281448 604
rect 281316 564 281448 592
rect 281316 552 281322 564
rect 281442 552 281448 564
rect 281500 552 281506 604
rect 384666 552 384672 604
rect 384724 592 384730 604
rect 384942 592 384948 604
rect 384724 564 384948 592
rect 384724 552 384730 564
rect 384942 552 384948 564
rect 385000 552 385006 604
rect 405918 552 405924 604
rect 405976 592 405982 604
rect 406102 592 406108 604
rect 405976 564 406108 592
rect 405976 552 405982 564
rect 406102 552 406108 564
rect 406160 552 406166 604
rect 463694 552 463700 604
rect 463752 592 463758 604
rect 464430 592 464436 604
rect 463752 564 464436 592
rect 463752 552 463758 564
rect 464430 552 464436 564
rect 464488 552 464494 604
rect 469214 552 469220 604
rect 469272 592 469278 604
rect 470318 592 470324 604
rect 469272 564 470324 592
rect 469272 552 469278 564
rect 470318 552 470324 564
rect 470376 552 470382 604
rect 471514 592 471520 604
rect 471475 564 471520 592
rect 471514 552 471520 564
rect 471572 552 471578 604
<< via1 >>
rect 202788 700952 202840 701004
rect 358820 700952 358872 701004
rect 170312 700884 170364 700936
rect 362960 700884 363012 700936
rect 328368 700816 328420 700868
rect 527180 700816 527232 700868
rect 329748 700748 329800 700800
rect 543464 700748 543516 700800
rect 154120 700680 154172 700732
rect 367100 700680 367152 700732
rect 137836 700612 137888 700664
rect 364340 700612 364392 700664
rect 105452 700544 105504 700596
rect 368480 700544 368532 700596
rect 89168 700476 89220 700528
rect 374000 700476 374052 700528
rect 72976 700408 73028 700460
rect 371240 700408 371292 700460
rect 40500 700340 40552 700392
rect 375380 700340 375432 700392
rect 24308 700272 24360 700324
rect 379520 700272 379572 700324
rect 218980 700204 219032 700256
rect 360200 700204 360252 700256
rect 336648 700136 336700 700188
rect 478512 700136 478564 700188
rect 335268 700068 335320 700120
rect 462320 700068 462372 700120
rect 235172 700000 235224 700052
rect 356060 700000 356112 700052
rect 267648 699932 267700 699984
rect 351920 699932 351972 699984
rect 283840 699864 283892 699916
rect 354680 699864 354732 699916
rect 343548 699796 343600 699848
rect 413652 699796 413704 699848
rect 340788 699728 340840 699780
rect 397460 699728 397512 699780
rect 300124 699660 300176 699712
rect 300768 699660 300820 699712
rect 332508 699660 332560 699712
rect 346400 699660 346452 699712
rect 347780 699660 347832 699712
rect 348792 699660 348844 699712
rect 321468 696940 321520 696992
rect 580172 696940 580224 696992
rect 429384 688576 429436 688628
rect 429844 688576 429896 688628
rect 559104 688576 559156 688628
rect 559656 688576 559708 688628
rect 364616 687760 364668 687812
rect 365168 687760 365220 687812
rect 324228 685856 324280 685908
rect 580172 685856 580224 685908
rect 364616 685788 364668 685840
rect 429292 684428 429344 684480
rect 559012 684428 559064 684480
rect 3516 681708 3568 681760
rect 382280 681708 382332 681760
rect 364524 676243 364576 676252
rect 364524 676209 364533 676243
rect 364533 676209 364567 676243
rect 364567 676209 364576 676243
rect 364524 676200 364576 676209
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 320088 673480 320140 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 386420 667904 386472 667956
rect 429660 666544 429712 666596
rect 494152 666544 494204 666596
rect 559380 666544 559432 666596
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 383660 652740 383712 652792
rect 315948 650020 316000 650072
rect 580172 650020 580224 650072
rect 429384 647232 429436 647284
rect 429476 647232 429528 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 429384 640364 429436 640416
rect 429476 640364 429528 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 317328 638936 317380 638988
rect 580172 638936 580224 638988
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 429292 630640 429344 630692
rect 429476 630640 429528 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 313188 626560 313240 626612
rect 580172 626560 580224 626612
rect 3424 623772 3476 623824
rect 387800 623772 387852 623824
rect 364616 618196 364668 618248
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 429292 611328 429344 611380
rect 429476 611328 429528 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 3424 609968 3476 610020
rect 391940 609968 391992 610020
rect 364524 608651 364576 608660
rect 364524 608617 364533 608651
rect 364533 608617 364567 608651
rect 364567 608617 364576 608651
rect 364524 608608 364576 608617
rect 429384 608583 429436 608592
rect 429384 608549 429393 608583
rect 429393 608549 429427 608583
rect 429427 608549 429436 608583
rect 429384 608540 429436 608549
rect 559104 608583 559156 608592
rect 559104 608549 559113 608583
rect 559113 608549 559147 608583
rect 559147 608549 559156 608583
rect 559104 608540 559156 608549
rect 309048 603100 309100 603152
rect 580172 603100 580224 603152
rect 429568 601672 429620 601724
rect 559288 601672 559340 601724
rect 364616 598927 364668 598936
rect 364616 598893 364625 598927
rect 364625 598893 364659 598927
rect 364659 598893 364668 598927
rect 364616 598884 364668 598893
rect 429568 598927 429620 598936
rect 429568 598893 429577 598927
rect 429577 598893 429611 598927
rect 429611 598893 429620 598927
rect 429568 598884 429620 598893
rect 559288 598927 559340 598936
rect 559288 598893 559297 598927
rect 559297 598893 559331 598927
rect 559331 598893 559340 598927
rect 559288 598884 559340 598893
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3240 594804 3292 594856
rect 390560 594804 390612 594856
rect 311808 592016 311860 592068
rect 580172 592016 580224 592068
rect 364708 589296 364760 589348
rect 429660 589296 429712 589348
rect 559380 589296 559432 589348
rect 344468 584672 344520 584724
rect 364708 584672 364760 584724
rect 300768 584604 300820 584656
rect 350816 584604 350868 584656
rect 338212 584536 338264 584588
rect 429660 584536 429712 584588
rect 331864 584468 331916 584520
rect 494244 584468 494296 584520
rect 325516 584400 325568 584452
rect 559380 584400 559432 584452
rect 298192 583652 298244 583704
rect 471244 583652 471296 583704
rect 256056 583584 256108 583636
rect 580540 583584 580592 583636
rect 245568 583516 245620 583568
rect 580264 583516 580316 583568
rect 6644 583448 6696 583500
rect 399208 583448 399260 583500
rect 4712 583380 4764 583432
rect 405556 583380 405608 583432
rect 10324 583312 10376 583364
rect 411904 583312 411956 583364
rect 6276 583244 6328 583296
rect 409788 583244 409840 583296
rect 3148 583176 3200 583228
rect 407672 583176 407724 583228
rect 13084 583108 13136 583160
rect 418160 583108 418212 583160
rect 14464 583040 14516 583092
rect 424508 583040 424560 583092
rect 3240 582972 3292 583024
rect 414020 582972 414072 583024
rect 5448 582904 5500 582956
rect 422392 582904 422444 582956
rect 15844 582836 15896 582888
rect 437112 582836 437164 582888
rect 4068 582768 4120 582820
rect 430856 582768 430908 582820
rect 5356 582700 5408 582752
rect 432972 582700 433024 582752
rect 3884 582632 3936 582684
rect 434996 582632 435048 582684
rect 17224 582564 17276 582616
rect 449808 582564 449860 582616
rect 5264 582496 5316 582548
rect 445576 582496 445628 582548
rect 3700 582428 3752 582480
rect 443460 582428 443512 582480
rect 5172 582360 5224 582412
rect 447692 582360 447744 582412
rect 302424 581680 302476 581732
rect 469588 581680 469640 581732
rect 296076 581612 296128 581664
rect 469772 581612 469824 581664
rect 289728 581544 289780 581596
rect 470508 581544 470560 581596
rect 287612 581476 287664 581528
rect 470416 581476 470468 581528
rect 283472 581408 283524 581460
rect 470324 581408 470376 581460
rect 281356 581340 281408 581392
rect 470232 581340 470284 581392
rect 275008 581272 275060 581324
rect 470140 581272 470192 581324
rect 268660 581204 268712 581256
rect 469956 581204 470008 581256
rect 304540 581136 304592 581188
rect 552664 581136 552716 581188
rect 264520 581068 264572 581120
rect 580908 581068 580960 581120
rect 4804 581000 4856 581052
rect 466644 581000 466696 581052
rect 300308 580320 300360 580372
rect 469680 580320 469732 580372
rect 262404 580252 262456 580304
rect 469864 580252 469916 580304
rect 306564 580184 306616 580236
rect 580172 580184 580224 580236
rect 6736 580116 6788 580168
rect 395068 580116 395120 580168
rect 6552 580048 6604 580100
rect 397092 580048 397144 580100
rect 6460 579980 6512 580032
rect 400956 579980 401008 580032
rect 6368 579912 6420 579964
rect 403164 579912 403216 579964
rect 3792 579844 3844 579896
rect 438860 579844 438912 579896
rect 5080 579776 5132 579828
rect 451556 579776 451608 579828
rect 4988 579708 5040 579760
rect 458272 579708 458324 579760
rect 6184 579640 6236 579692
rect 464252 579640 464304 579692
rect 271144 579368 271196 579420
rect 252100 579343 252152 579352
rect 252100 579309 252109 579343
rect 252109 579309 252143 579343
rect 252143 579309 252152 579343
rect 252100 579300 252152 579309
rect 254216 579343 254268 579352
rect 254216 579309 254225 579343
rect 254225 579309 254259 579343
rect 254259 579309 254268 579343
rect 254216 579300 254268 579309
rect 258448 579300 258500 579352
rect 260656 579300 260708 579352
rect 266912 579300 266964 579352
rect 273076 579300 273128 579352
rect 277308 579300 277360 579352
rect 279608 579300 279660 579352
rect 285680 579300 285732 579352
rect 292120 579300 292172 579352
rect 415676 579411 415728 579420
rect 415676 579377 415685 579411
rect 415685 579377 415719 579411
rect 415719 579377 415728 579411
rect 415676 579368 415728 579377
rect 428372 579411 428424 579420
rect 428372 579377 428381 579411
rect 428381 579377 428415 579411
rect 428415 579377 428424 579411
rect 428372 579368 428424 579377
rect 453580 579411 453632 579420
rect 453580 579377 453589 579411
rect 453589 579377 453623 579411
rect 453623 579377 453632 579411
rect 453580 579368 453632 579377
rect 455788 579411 455840 579420
rect 455788 579377 455797 579411
rect 455797 579377 455831 579411
rect 455831 579377 455840 579411
rect 455788 579368 455840 579377
rect 441068 579343 441120 579352
rect 441068 579309 441077 579343
rect 441077 579309 441111 579343
rect 441111 579309 441120 579343
rect 441068 579300 441120 579309
rect 579804 579164 579856 579216
rect 579896 579096 579948 579148
rect 580080 579028 580132 579080
rect 579988 578960 580040 579012
rect 580172 578892 580224 578944
rect 580816 578824 580868 578876
rect 580632 578756 580684 578808
rect 580724 578688 580776 578740
rect 580356 578620 580408 578672
rect 580448 578552 580500 578604
rect 3332 578484 3384 578536
rect 3976 578416 4028 578468
rect 3608 578348 3660 578400
rect 3424 578280 3476 578332
rect 3516 578212 3568 578264
rect 470048 577872 470100 577924
rect 3056 568284 3108 568336
rect 6736 568284 6788 568336
rect 579712 567128 579764 567180
rect 580908 567128 580960 567180
rect 579712 557608 579764 557660
rect 580908 557540 580960 557592
rect 469588 557472 469640 557524
rect 579712 557472 579764 557524
rect 3056 553324 3108 553376
rect 6644 553324 6696 553376
rect 579620 547816 579672 547868
rect 580908 547816 580960 547868
rect 552664 546388 552716 546440
rect 579712 546388 579764 546440
rect 3056 538636 3108 538688
rect 6552 538636 6604 538688
rect 579620 538228 579672 538280
rect 580908 538228 580960 538280
rect 469680 534012 469732 534064
rect 579712 534012 579764 534064
rect 579712 528504 579764 528556
rect 580908 528504 580960 528556
rect 579712 518916 579764 518968
rect 580908 518916 580960 518968
rect 469772 510552 469824 510604
rect 579712 510552 579764 510604
rect 3056 510212 3108 510264
rect 6460 510212 6512 510264
rect 579712 509192 579764 509244
rect 580908 509192 580960 509244
rect 579712 499604 579764 499656
rect 580908 499536 580960 499588
rect 471244 499468 471296 499520
rect 579712 499468 579764 499520
rect 2780 495524 2832 495576
rect 4712 495524 4764 495576
rect 579712 489812 579764 489864
rect 580908 489812 580960 489864
rect 2964 481108 3016 481160
rect 6368 481108 6420 481160
rect 579712 480224 579764 480276
rect 580908 480224 580960 480276
rect 579620 470500 579672 470552
rect 580908 470500 580960 470552
rect 470508 463632 470560 463684
rect 579712 463632 579764 463684
rect 579620 460912 579672 460964
rect 580908 460912 580960 460964
rect 579804 451188 579856 451240
rect 580908 451188 580960 451240
rect 579804 441600 579856 441652
rect 580908 441600 580960 441652
rect 470416 440172 470468 440224
rect 579804 440172 579856 440224
rect 3148 438812 3200 438864
rect 10324 438812 10376 438864
rect 579804 431876 579856 431928
rect 580908 431876 580960 431928
rect 3148 424056 3200 424108
rect 6276 424056 6328 424108
rect 579804 422288 579856 422340
rect 580908 422288 580960 422340
rect 470324 416712 470376 416764
rect 579804 416712 579856 416764
rect 579804 412564 579856 412616
rect 580908 412564 580960 412616
rect 579804 402976 579856 403028
rect 580908 402976 580960 403028
rect 470232 393252 470284 393304
rect 579896 393252 579948 393304
rect 579804 393184 579856 393236
rect 580908 393252 580960 393304
rect 579804 384276 579856 384328
rect 580908 384276 580960 384328
rect 3240 380808 3292 380860
rect 13084 380808 13136 380860
rect 579988 361224 580040 361276
rect 580908 361224 580960 361276
rect 579804 360136 579856 360188
rect 579988 360136 580040 360188
rect 470140 346332 470192 346384
rect 579804 346332 579856 346384
rect 580080 345040 580132 345092
rect 580908 345040 580960 345092
rect 580080 344904 580132 344956
rect 580908 344904 580960 344956
rect 71044 338036 71096 338088
rect 254952 338036 255004 338088
rect 284392 338079 284444 338088
rect 284392 338045 284401 338079
rect 284401 338045 284435 338079
rect 284435 338045 284444 338079
rect 284392 338036 284444 338045
rect 354404 338036 354456 338088
rect 358084 338036 358136 338088
rect 371516 338036 371568 338088
rect 376668 338036 376720 338088
rect 380348 338036 380400 338088
rect 406292 338036 406344 338088
rect 417424 338036 417476 338088
rect 419080 338036 419132 338088
rect 431408 338036 431460 338088
rect 435732 338036 435784 338088
rect 499580 338036 499632 338088
rect 66904 337968 66956 338020
rect 252008 337968 252060 338020
rect 306196 337968 306248 338020
rect 355876 337968 355928 338020
rect 364248 337968 364300 338020
rect 376760 337968 376812 338020
rect 61384 337900 61436 337952
rect 247592 337900 247644 337952
rect 303160 337900 303212 337952
rect 352932 337900 352984 337952
rect 355324 337900 355376 337952
rect 370044 337900 370096 337952
rect 371148 337900 371200 337952
rect 382280 337968 382332 338020
rect 404360 337968 404412 338020
rect 414664 337968 414716 338020
rect 429752 337968 429804 338020
rect 437204 337968 437256 338020
rect 442356 337968 442408 338020
rect 446036 337968 446088 338020
rect 451832 337968 451884 338020
rect 461676 337968 461728 338020
rect 400404 337900 400456 337952
rect 413284 337900 413336 337952
rect 413652 337900 413704 337952
rect 420184 337900 420236 337952
rect 420552 337900 420604 337952
rect 454776 337900 454828 337952
rect 460664 337900 460716 337952
rect 525064 337968 525116 338020
rect 467104 337900 467156 337952
rect 467748 337900 467800 337952
rect 468024 337900 468076 337952
rect 469128 337900 469180 337952
rect 527824 337900 527876 337952
rect 57244 337832 57296 337884
rect 247132 337832 247184 337884
rect 290464 337832 290516 337884
rect 347044 337832 347096 337884
rect 348424 337832 348476 337884
rect 365628 337832 365680 337884
rect 377404 337832 377456 337884
rect 398472 337832 398524 337884
rect 408776 337832 408828 337884
rect 414204 337832 414256 337884
rect 415308 337832 415360 337884
rect 50344 337764 50396 337816
rect 244188 337764 244240 337816
rect 259644 337764 259696 337816
rect 260104 337764 260156 337816
rect 288256 337764 288308 337816
rect 32404 337696 32456 337748
rect 237840 337696 237892 337748
rect 248512 337696 248564 337748
rect 249524 337696 249576 337748
rect 251456 337696 251508 337748
rect 252468 337696 252520 337748
rect 254584 337696 254636 337748
rect 262312 337696 262364 337748
rect 351920 337764 351972 337816
rect 358728 337764 358780 337816
rect 348516 337696 348568 337748
rect 39304 337628 39356 337680
rect 244648 337628 244700 337680
rect 260104 337628 260156 337680
rect 277032 337628 277084 337680
rect 285588 337628 285640 337680
rect 336096 337628 336148 337680
rect 344560 337628 344612 337680
rect 349988 337628 350040 337680
rect 35164 337560 35216 337612
rect 241704 337560 241756 337612
rect 255964 337560 256016 337612
rect 261392 337560 261444 337612
rect 279976 337560 280028 337612
rect 281448 337560 281500 337612
rect 345572 337560 345624 337612
rect 350172 337560 350224 337612
rect 28264 337492 28316 337544
rect 19984 337424 20036 337476
rect 234344 337424 234396 337476
rect 253204 337492 253256 337544
rect 259368 337492 259420 337544
rect 238300 337424 238352 337476
rect 258724 337424 258776 337476
rect 275560 337492 275612 337544
rect 275928 337492 275980 337544
rect 13084 337356 13136 337408
rect 233516 337356 233568 337408
rect 233884 337356 233936 337408
rect 241244 337356 241296 337408
rect 250444 337356 250496 337408
rect 253480 337356 253532 337408
rect 257344 337356 257396 337408
rect 269672 337424 269724 337476
rect 271788 337424 271840 337476
rect 341616 337492 341668 337544
rect 344376 337492 344428 337544
rect 354864 337628 354916 337680
rect 356704 337628 356756 337680
rect 360752 337628 360804 337680
rect 362868 337764 362920 337816
rect 378876 337764 378928 337816
rect 388444 337764 388496 337816
rect 389180 337764 389232 337816
rect 407304 337764 407356 337816
rect 416136 337764 416188 337816
rect 416688 337764 416740 337816
rect 417608 337832 417660 337884
rect 455604 337832 455656 337884
rect 457720 337832 457772 337884
rect 523684 337832 523736 337884
rect 420276 337764 420328 337816
rect 422024 337764 422076 337816
rect 438124 337764 438176 337816
rect 438676 337764 438728 337816
rect 369584 337696 369636 337748
rect 351184 337560 351236 337612
rect 375932 337696 375984 337748
rect 380164 337696 380216 337748
rect 381360 337696 381412 337748
rect 381544 337696 381596 337748
rect 382832 337696 382884 337748
rect 384948 337696 385000 337748
rect 388168 337696 388220 337748
rect 398932 337696 398984 337748
rect 351828 337492 351880 337544
rect 344100 337424 344152 337476
rect 349068 337424 349120 337476
rect 366916 337560 366968 337612
rect 376576 337628 376628 337680
rect 384304 337628 384356 337680
rect 387708 337628 387760 337680
rect 398012 337628 398064 337680
rect 399484 337628 399536 337680
rect 403348 337696 403400 337748
rect 406384 337628 406436 337680
rect 410248 337696 410300 337748
rect 411076 337696 411128 337748
rect 411260 337628 411312 337680
rect 412364 337628 412416 337680
rect 266728 337356 266780 337408
rect 269028 337356 269080 337408
rect 340236 337356 340288 337408
rect 340788 337356 340840 337408
rect 79324 337288 79376 337340
rect 260840 337288 260892 337340
rect 271328 337288 271380 337340
rect 132500 337220 132552 337272
rect 142068 337220 142120 337272
rect 151820 337220 151872 337272
rect 161388 337220 161440 337272
rect 171140 337220 171192 337272
rect 180708 337220 180760 337272
rect 190460 337220 190512 337272
rect 200028 337220 200080 337272
rect 209780 337220 209832 337272
rect 219348 337220 219400 337272
rect 229192 337220 229244 337272
rect 234620 337220 234672 337272
rect 257896 337220 257948 337272
rect 258816 337220 258868 337272
rect 272616 337220 272668 337272
rect 272800 337220 272852 337272
rect 309784 337288 309836 337340
rect 84844 337152 84896 337204
rect 263784 337152 263836 337204
rect 297916 337152 297968 337204
rect 77944 336948 77996 337000
rect 100668 337084 100720 337136
rect 271144 337084 271196 337136
rect 312728 337220 312780 337272
rect 361764 337288 361816 337340
rect 372068 337424 372120 337476
rect 373908 337492 373960 337544
rect 383292 337560 383344 337612
rect 404820 337560 404872 337612
rect 412732 337560 412784 337612
rect 413836 337560 413888 337612
rect 415584 337696 415636 337748
rect 416504 337696 416556 337748
rect 417056 337696 417108 337748
rect 417976 337696 418028 337748
rect 418528 337696 418580 337748
rect 419448 337696 419500 337748
rect 419540 337696 419592 337748
rect 420828 337696 420880 337748
rect 421472 337696 421524 337748
rect 422208 337696 422260 337748
rect 422484 337696 422536 337748
rect 424416 337696 424468 337748
rect 425428 337696 425480 337748
rect 428464 337696 428516 337748
rect 429384 337696 429436 337748
rect 430488 337696 430540 337748
rect 427084 337628 427136 337680
rect 432328 337696 432380 337748
rect 433156 337696 433208 337748
rect 433708 337696 433760 337748
rect 434628 337696 434680 337748
rect 435180 337696 435232 337748
rect 436008 337696 436060 337748
rect 436192 337696 436244 337748
rect 437388 337696 437440 337748
rect 439136 337696 439188 337748
rect 440148 337696 440200 337748
rect 440608 337764 440660 337816
rect 441528 337764 441580 337816
rect 442080 337764 442132 337816
rect 442908 337764 442960 337816
rect 444564 337764 444616 337816
rect 445668 337764 445720 337816
rect 448980 337764 449032 337816
rect 451372 337764 451424 337816
rect 452476 337764 452528 337816
rect 452844 337764 452896 337816
rect 453764 337764 453816 337816
rect 454316 337764 454368 337816
rect 455236 337764 455288 337816
rect 455788 337764 455840 337816
rect 456616 337764 456668 337816
rect 460204 337764 460256 337816
rect 460756 337764 460808 337816
rect 520924 337764 520976 337816
rect 506480 337696 506532 337748
rect 421196 337560 421248 337612
rect 426808 337560 426860 337612
rect 430856 337628 430908 337680
rect 431868 337628 431920 337680
rect 434720 337628 434772 337680
rect 435916 337628 435968 337680
rect 436652 337628 436704 337680
rect 437296 337628 437348 337680
rect 440240 337628 440292 337680
rect 443552 337628 443604 337680
rect 444288 337628 444340 337680
rect 445024 337628 445076 337680
rect 445576 337628 445628 337680
rect 446496 337628 446548 337680
rect 447048 337628 447100 337680
rect 448244 337628 448296 337680
rect 448428 337628 448480 337680
rect 449900 337628 449952 337680
rect 451004 337628 451056 337680
rect 518164 337628 518216 337680
rect 428372 337560 428424 337612
rect 431224 337560 431276 337612
rect 431316 337560 431368 337612
rect 449164 337560 449216 337612
rect 450452 337560 450504 337612
rect 451188 337560 451240 337612
rect 453304 337560 453356 337612
rect 453948 337560 454000 337612
rect 521016 337560 521068 337612
rect 375288 337492 375340 337544
rect 383752 337492 383804 337544
rect 405832 337492 405884 337544
rect 426440 337492 426492 337544
rect 442264 337492 442316 337544
rect 447508 337492 447560 337544
rect 448428 337492 448480 337544
rect 516784 337492 516836 337544
rect 374460 337424 374512 337476
rect 381820 337424 381872 337476
rect 387064 337424 387116 337476
rect 388720 337424 388772 337476
rect 397000 337424 397052 337476
rect 405924 337424 405976 337476
rect 409144 337424 409196 337476
rect 433524 337424 433576 337476
rect 437664 337424 437716 337476
rect 438676 337424 438728 337476
rect 443092 337424 443144 337476
rect 514024 337424 514076 337476
rect 369768 337356 369820 337408
rect 382188 337356 382240 337408
rect 386696 337356 386748 337408
rect 400956 337356 401008 337408
rect 402244 337356 402296 337408
rect 409236 337356 409288 337408
rect 433984 337356 434036 337408
rect 434260 337356 434312 337408
rect 439504 337356 439556 337408
rect 510620 337356 510672 337408
rect 333244 337220 333296 337272
rect 367008 337288 367060 337340
rect 380808 337288 380860 337340
rect 312544 337152 312596 337204
rect 341800 337152 341852 337204
rect 348976 337152 349028 337204
rect 359464 337152 359516 337204
rect 363696 337152 363748 337204
rect 372988 337220 373040 337272
rect 366640 337152 366692 337204
rect 401876 337152 401928 337204
rect 416964 337152 417016 337204
rect 420000 337288 420052 337340
rect 420736 337288 420788 337340
rect 421012 337288 421064 337340
rect 423496 337220 423548 337272
rect 460296 337220 460348 337272
rect 463884 337288 463936 337340
rect 465080 337288 465132 337340
rect 466368 337288 466420 337340
rect 470600 337288 470652 337340
rect 470692 337288 470744 337340
rect 529204 337288 529256 337340
rect 463608 337220 463660 337272
rect 469496 337220 469548 337272
rect 530584 337220 530636 337272
rect 424324 337152 424376 337204
rect 427912 337152 427964 337204
rect 432788 337152 432840 337204
rect 492680 337152 492732 337204
rect 314200 337084 314252 337136
rect 316684 337084 316736 337136
rect 342904 337084 342956 337136
rect 355968 337084 356020 337136
rect 369124 337084 369176 337136
rect 371056 337084 371108 337136
rect 415124 337084 415176 337136
rect 421564 337084 421616 337136
rect 429844 337084 429896 337136
rect 485780 337084 485832 337136
rect 95884 337016 95936 337068
rect 265256 337016 265308 337068
rect 335268 337016 335320 337068
rect 367652 337016 367704 337068
rect 397460 337016 397512 337068
rect 403624 337016 403676 337068
rect 407764 337016 407816 337068
rect 409144 337016 409196 337068
rect 426900 337016 426952 337068
rect 477592 337016 477644 337068
rect 107568 336948 107620 337000
rect 274088 336948 274140 337000
rect 319444 336948 319496 337000
rect 353392 336948 353444 337000
rect 378048 336948 378100 337000
rect 385224 336948 385276 337000
rect 401416 336948 401468 337000
rect 405004 336948 405056 337000
rect 475384 336948 475436 337000
rect 102784 336880 102836 336932
rect 268200 336880 268252 336932
rect 118608 336812 118660 336864
rect 278504 336812 278556 336864
rect 125508 336744 125560 336796
rect 281172 336744 281224 336796
rect 327724 336744 327776 336796
rect 345480 336880 345532 336932
rect 345940 336880 345992 336932
rect 360292 336880 360344 336932
rect 380808 336880 380860 336932
rect 386236 336880 386288 336932
rect 392124 336880 392176 336932
rect 393596 336880 393648 336932
rect 393872 336880 393924 336932
rect 397460 336880 397512 336932
rect 423956 336880 424008 336932
rect 466552 336880 466604 336932
rect 470508 336880 470560 336932
rect 344284 336812 344336 336864
rect 357348 336812 357400 336864
rect 362224 336812 362276 336864
rect 365168 336812 365220 336864
rect 381636 336812 381688 336864
rect 384764 336812 384816 336864
rect 396080 336812 396132 336864
rect 398196 336812 398248 336864
rect 424968 336812 425020 336864
rect 439596 336812 439648 336864
rect 441620 336812 441672 336864
rect 443644 336812 443696 336864
rect 456800 336812 456852 336864
rect 458088 336812 458140 336864
rect 459192 336812 459244 336864
rect 460204 336812 460256 336864
rect 469220 336812 469272 336864
rect 343088 336744 343140 336796
rect 251824 336676 251876 336728
rect 256424 336676 256476 336728
rect 330576 336676 330628 336728
rect 351460 336744 351512 336796
rect 352564 336744 352616 336796
rect 357808 336744 357860 336796
rect 363604 336744 363656 336796
rect 364708 336744 364760 336796
rect 370504 336744 370556 336796
rect 372528 336744 372580 336796
rect 376024 336744 376076 336796
rect 376944 336744 376996 336796
rect 377680 336744 377732 336796
rect 378416 336744 378468 336796
rect 394056 336744 394108 336796
rect 394608 336744 394660 336796
rect 395068 336744 395120 336796
rect 395896 336744 395948 336796
rect 396540 336744 396592 336796
rect 398104 336744 398156 336796
rect 424600 336744 424652 336796
rect 457260 336744 457312 336796
rect 457996 336744 458048 336796
rect 458272 336744 458324 336796
rect 459468 336744 459520 336796
rect 459744 336744 459796 336796
rect 460848 336744 460900 336796
rect 461216 336744 461268 336796
rect 462136 336744 462188 336796
rect 462688 336744 462740 336796
rect 463516 336744 463568 336796
rect 464160 336744 464212 336796
rect 464988 336744 465040 336796
rect 465080 336744 465132 336796
rect 509884 336812 509936 336864
rect 374552 336676 374604 336728
rect 375840 336719 375892 336728
rect 375840 336685 375849 336719
rect 375849 336685 375883 336719
rect 375883 336685 375892 336719
rect 375840 336676 375892 336685
rect 424968 336676 425020 336728
rect 505744 336744 505796 336796
rect 247684 336472 247736 336524
rect 248604 336472 248656 336524
rect 249064 336200 249116 336252
rect 250536 336200 250588 336252
rect 331404 336107 331456 336116
rect 331404 336073 331413 336107
rect 331413 336073 331447 336107
rect 331447 336073 331456 336107
rect 331404 336064 331456 336073
rect 331220 335860 331272 335912
rect 331496 335860 331548 335912
rect 236184 335656 236236 335708
rect 237012 335656 237064 335708
rect 302240 335656 302292 335708
rect 302700 335656 302752 335708
rect 316040 335656 316092 335708
rect 316868 335656 316920 335708
rect 318800 335656 318852 335708
rect 319812 335656 319864 335708
rect 332692 335656 332744 335708
rect 333428 335656 333480 335708
rect 334072 335656 334124 335708
rect 334900 335656 334952 335708
rect 236092 335588 236144 335640
rect 236552 335588 236604 335640
rect 241612 335588 241664 335640
rect 242348 335588 242400 335640
rect 260932 335588 260984 335640
rect 261484 335588 261536 335640
rect 263692 335588 263744 335640
rect 264428 335588 264480 335640
rect 265072 335588 265124 335640
rect 265900 335588 265952 335640
rect 266452 335588 266504 335640
rect 267372 335588 267424 335640
rect 280252 335588 280304 335640
rect 280620 335588 280672 335640
rect 281540 335588 281592 335640
rect 282092 335588 282144 335640
rect 283012 335588 283064 335640
rect 283564 335588 283616 335640
rect 285680 335588 285732 335640
rect 285956 335588 286008 335640
rect 286048 335588 286100 335640
rect 286600 335588 286652 335640
rect 287060 335588 287112 335640
rect 287980 335588 288032 335640
rect 288440 335588 288492 335640
rect 289452 335588 289504 335640
rect 292764 335588 292816 335640
rect 293316 335588 293368 335640
rect 298284 335588 298336 335640
rect 298652 335588 298704 335640
rect 300860 335588 300912 335640
rect 301228 335588 301280 335640
rect 303620 335588 303672 335640
rect 304172 335588 304224 335640
rect 307760 335588 307812 335640
rect 308588 335588 308640 335640
rect 309140 335588 309192 335640
rect 310060 335588 310112 335640
rect 310520 335588 310572 335640
rect 311532 335588 311584 335640
rect 314660 335588 314712 335640
rect 315396 335588 315448 335640
rect 316132 335588 316184 335640
rect 316316 335588 316368 335640
rect 317420 335588 317472 335640
rect 318340 335588 318392 335640
rect 318892 335588 318944 335640
rect 319260 335588 319312 335640
rect 320180 335588 320232 335640
rect 320732 335588 320784 335640
rect 321652 335588 321704 335640
rect 322204 335588 322256 335640
rect 329840 335588 329892 335640
rect 330116 335588 330168 335640
rect 332600 335588 332652 335640
rect 333060 335588 333112 335640
rect 333980 335588 334032 335640
rect 334532 335588 334584 335640
rect 338120 335588 338172 335640
rect 338948 335588 339000 335640
rect 356152 335588 356204 335640
rect 356612 335588 356664 335640
rect 359004 335588 359056 335640
rect 359372 335588 359424 335640
rect 363052 335588 363104 335640
rect 363788 335588 363840 335640
rect 367284 335588 367336 335640
rect 367928 335588 367980 335640
rect 458916 335588 458968 335640
rect 459376 335588 459428 335640
rect 341708 335563 341760 335572
rect 341708 335529 341717 335563
rect 341717 335529 341751 335563
rect 341751 335529 341760 335563
rect 341708 335520 341760 335529
rect 235080 335452 235132 335504
rect 235632 335452 235684 335504
rect 245844 335452 245896 335504
rect 246672 335452 246724 335504
rect 331312 335452 331364 335504
rect 331956 335452 332008 335504
rect 580080 335384 580132 335436
rect 581000 335384 581052 335436
rect 580080 335248 580132 335300
rect 581000 335248 581052 335300
rect 284484 335180 284536 335232
rect 278780 334772 278832 334824
rect 278964 334772 279016 334824
rect 303068 334704 303120 334756
rect 258172 334568 258224 334620
rect 258540 334568 258592 334620
rect 328552 334500 328604 334552
rect 329012 334500 329064 334552
rect 250628 334432 250680 334484
rect 270776 334296 270828 334348
rect 271236 334296 271288 334348
rect 272248 334296 272300 334348
rect 272708 334296 272760 334348
rect 247132 334160 247184 334212
rect 248144 334160 248196 334212
rect 335360 334160 335412 334212
rect 336004 334160 336056 334212
rect 305000 333752 305052 333804
rect 305644 333752 305696 333804
rect 301044 333276 301096 333328
rect 301688 333276 301740 333328
rect 325884 333276 325936 333328
rect 326620 333276 326672 333328
rect 361672 333276 361724 333328
rect 362316 333276 362368 333328
rect 306472 333072 306524 333124
rect 306656 333072 306708 333124
rect 262588 333004 262640 333056
rect 263048 333004 263100 333056
rect 284668 332528 284720 332580
rect 285128 332528 285180 332580
rect 242992 332052 243044 332104
rect 243452 332052 243504 332104
rect 336740 331984 336792 332036
rect 336924 331984 336976 332036
rect 284300 331916 284352 331968
rect 284576 331916 284628 331968
rect 357348 331848 357400 331900
rect 357992 331848 358044 331900
rect 299572 331304 299624 331356
rect 336832 331304 336884 331356
rect 259644 331168 259696 331220
rect 259828 331168 259880 331220
rect 262588 331168 262640 331220
rect 262772 331168 262824 331220
rect 389732 331236 389784 331288
rect 336832 331168 336884 331220
rect 389640 331168 389692 331220
rect 299572 331032 299624 331084
rect 299480 330964 299532 331016
rect 299848 330964 299900 331016
rect 321468 329128 321520 329180
rect 347504 328516 347556 328568
rect 250168 328491 250220 328500
rect 250168 328457 250177 328491
rect 250177 328457 250211 328491
rect 250211 328457 250220 328491
rect 250168 328448 250220 328457
rect 278872 328448 278924 328500
rect 279056 328448 279108 328500
rect 288808 328448 288860 328500
rect 289084 328448 289136 328500
rect 302516 328491 302568 328500
rect 302516 328457 302525 328491
rect 302525 328457 302559 328491
rect 302559 328457 302568 328491
rect 302516 328448 302568 328457
rect 303896 328448 303948 328500
rect 304632 328448 304684 328500
rect 323308 328448 323360 328500
rect 323676 328448 323728 328500
rect 324688 328448 324740 328500
rect 325056 328448 325108 328500
rect 338856 328448 338908 328500
rect 339776 328448 339828 328500
rect 340328 328448 340380 328500
rect 341432 328448 341484 328500
rect 372712 328448 372764 328500
rect 373264 328448 373316 328500
rect 259828 328423 259880 328432
rect 259828 328389 259837 328423
rect 259837 328389 259871 328423
rect 259871 328389 259880 328423
rect 259828 328380 259880 328389
rect 295524 328380 295576 328432
rect 295708 328380 295760 328432
rect 296812 328380 296864 328432
rect 296996 328380 297048 328432
rect 389640 328380 389692 328432
rect 470600 328423 470652 328432
rect 470600 328389 470609 328423
rect 470609 328389 470643 328423
rect 470643 328389 470652 328423
rect 470600 328380 470652 328389
rect 330208 327199 330260 327208
rect 330208 327165 330217 327199
rect 330217 327165 330251 327199
rect 330251 327165 330260 327199
rect 330208 327156 330260 327165
rect 327264 327088 327316 327140
rect 327448 327088 327500 327140
rect 331404 327131 331456 327140
rect 331404 327097 331413 327131
rect 331413 327097 331447 327131
rect 331447 327097 331456 327131
rect 331404 327088 331456 327097
rect 374460 327131 374512 327140
rect 374460 327097 374469 327131
rect 374469 327097 374503 327131
rect 374503 327097 374512 327131
rect 374460 327088 374512 327097
rect 375932 327088 375984 327140
rect 302516 327020 302568 327072
rect 302608 327020 302660 327072
rect 357440 327063 357492 327072
rect 357440 327029 357449 327063
rect 357449 327029 357483 327063
rect 357483 327029 357492 327063
rect 357440 327020 357492 327029
rect 360476 327020 360528 327072
rect 463700 325660 463752 325712
rect 463884 325660 463936 325712
rect 580080 325660 580132 325712
rect 580908 325660 580960 325712
rect 3332 324232 3384 324284
rect 14464 324232 14516 324284
rect 376852 323552 376904 323604
rect 377128 323552 377180 323604
rect 470048 322872 470100 322924
rect 580080 322872 580132 322924
rect 239128 321648 239180 321700
rect 235080 321580 235132 321632
rect 230756 321512 230808 321564
rect 230940 321512 230992 321564
rect 232228 321512 232280 321564
rect 232412 321512 232464 321564
rect 251456 321580 251508 321632
rect 239128 321512 239180 321564
rect 235080 321444 235132 321496
rect 286048 321580 286100 321632
rect 310796 321580 310848 321632
rect 337200 321623 337252 321632
rect 337200 321589 337209 321623
rect 337209 321589 337243 321623
rect 337243 321589 337252 321623
rect 337200 321580 337252 321589
rect 341432 321623 341484 321632
rect 341432 321589 341441 321623
rect 341441 321589 341475 321623
rect 341475 321589 341484 321623
rect 341432 321580 341484 321589
rect 285956 321512 286008 321564
rect 310888 321444 310940 321496
rect 251548 321376 251600 321428
rect 337200 320875 337252 320884
rect 337200 320841 337209 320875
rect 337209 320841 337243 320875
rect 337243 320841 337252 320875
rect 337200 320832 337252 320841
rect 259920 318792 259972 318844
rect 294236 318792 294288 318844
rect 294328 318792 294380 318844
rect 306748 318792 306800 318844
rect 306840 318792 306892 318844
rect 341432 318835 341484 318844
rect 341432 318801 341441 318835
rect 341441 318801 341475 318835
rect 341475 318801 341484 318835
rect 341432 318792 341484 318801
rect 374368 318792 374420 318844
rect 374460 318792 374512 318844
rect 375840 318792 375892 318844
rect 375932 318792 375984 318844
rect 389548 318835 389600 318844
rect 389548 318801 389557 318835
rect 389557 318801 389591 318835
rect 389591 318801 389600 318835
rect 389548 318792 389600 318801
rect 470600 318835 470652 318844
rect 470600 318801 470609 318835
rect 470609 318801 470643 318835
rect 470643 318801 470652 318835
rect 470600 318792 470652 318801
rect 230940 318724 230992 318776
rect 236276 318767 236328 318776
rect 236276 318733 236285 318767
rect 236285 318733 236319 318767
rect 236319 318733 236328 318767
rect 236276 318724 236328 318733
rect 239220 318767 239272 318776
rect 239220 318733 239229 318767
rect 239229 318733 239263 318767
rect 239263 318733 239272 318767
rect 239220 318724 239272 318733
rect 284760 318724 284812 318776
rect 285956 318724 286008 318776
rect 286140 318724 286192 318776
rect 357532 317432 357584 317484
rect 360384 317475 360436 317484
rect 360384 317441 360393 317475
rect 360393 317441 360427 317475
rect 360427 317441 360436 317475
rect 360384 317432 360436 317441
rect 291568 317364 291620 317416
rect 299848 317364 299900 317416
rect 325976 317364 326028 317416
rect 337200 317407 337252 317416
rect 337200 317373 337209 317407
rect 337209 317373 337243 317407
rect 337243 317373 337252 317407
rect 337200 317364 337252 317373
rect 375840 317407 375892 317416
rect 375840 317373 375849 317407
rect 375849 317373 375883 317407
rect 375883 317373 375892 317407
rect 375840 317364 375892 317373
rect 377128 317364 377180 317416
rect 377312 317364 377364 317416
rect 291660 317296 291712 317348
rect 579988 316072 580040 316124
rect 581000 316072 581052 316124
rect 262680 315936 262732 315988
rect 580080 315936 580132 315988
rect 581000 315936 581052 315988
rect 284944 314168 284996 314220
rect 250168 313964 250220 314016
rect 288624 313896 288676 313948
rect 288808 313896 288860 313948
rect 250168 313828 250220 313880
rect 273628 313420 273680 313472
rect 272248 311924 272300 311976
rect 259736 311856 259788 311908
rect 259920 311856 259972 311908
rect 273444 311899 273496 311908
rect 273444 311865 273453 311899
rect 273453 311865 273487 311899
rect 273487 311865 273496 311899
rect 273444 311856 273496 311865
rect 306840 311924 306892 311976
rect 310888 311967 310940 311976
rect 310888 311933 310897 311967
rect 310897 311933 310931 311967
rect 310931 311933 310940 311967
rect 310888 311924 310940 311933
rect 323308 311924 323360 311976
rect 374368 311924 374420 311976
rect 323216 311856 323268 311908
rect 341248 311856 341300 311908
rect 341432 311856 341484 311908
rect 244464 311831 244516 311840
rect 244464 311797 244473 311831
rect 244473 311797 244507 311831
rect 244507 311797 244516 311831
rect 244464 311788 244516 311797
rect 272248 311788 272300 311840
rect 306748 311788 306800 311840
rect 337200 311763 337252 311772
rect 337200 311729 337209 311763
rect 337209 311729 337243 311763
rect 337243 311729 337252 311763
rect 337200 311720 337252 311729
rect 374460 311720 374512 311772
rect 236276 309247 236328 309256
rect 236276 309213 236285 309247
rect 236285 309213 236319 309247
rect 236319 309213 236328 309247
rect 236276 309204 236328 309213
rect 230848 309179 230900 309188
rect 230848 309145 230857 309179
rect 230857 309145 230891 309179
rect 230891 309145 230900 309179
rect 230848 309136 230900 309145
rect 239220 309179 239272 309188
rect 239220 309145 239229 309179
rect 239229 309145 239263 309179
rect 239263 309145 239272 309179
rect 239220 309136 239272 309145
rect 244464 309179 244516 309188
rect 244464 309145 244473 309179
rect 244473 309145 244507 309179
rect 244507 309145 244516 309179
rect 244464 309136 244516 309145
rect 267740 309136 267792 309188
rect 267832 309136 267884 309188
rect 295616 309204 295668 309256
rect 296904 309204 296956 309256
rect 389364 309136 389416 309188
rect 389548 309136 389600 309188
rect 236276 309111 236328 309120
rect 236276 309077 236285 309111
rect 236285 309077 236319 309111
rect 236319 309077 236328 309111
rect 236276 309068 236328 309077
rect 259736 309068 259788 309120
rect 295524 309068 295576 309120
rect 296812 309068 296864 309120
rect 327172 309068 327224 309120
rect 327264 309068 327316 309120
rect 341248 309068 341300 309120
rect 357808 309111 357860 309120
rect 357808 309077 357817 309111
rect 357817 309077 357851 309111
rect 357851 309077 357860 309111
rect 357808 309068 357860 309077
rect 358728 309111 358780 309120
rect 358728 309077 358737 309111
rect 358737 309077 358771 309111
rect 358771 309077 358780 309111
rect 358728 309068 358780 309077
rect 470600 309111 470652 309120
rect 470600 309077 470609 309111
rect 470609 309077 470643 309111
rect 470643 309077 470652 309111
rect 470600 309068 470652 309077
rect 389364 309000 389416 309052
rect 2780 308796 2832 308848
rect 5448 308796 5500 308848
rect 310704 307844 310756 307896
rect 325884 307819 325936 307828
rect 325884 307785 325893 307819
rect 325893 307785 325927 307819
rect 325927 307785 325936 307819
rect 325884 307776 325936 307785
rect 375840 307819 375892 307828
rect 375840 307785 375849 307819
rect 375849 307785 375883 307819
rect 375883 307785 375892 307819
rect 375840 307776 375892 307785
rect 310704 307751 310756 307760
rect 310704 307717 310713 307751
rect 310713 307717 310747 307751
rect 310747 307717 310756 307751
rect 310704 307708 310756 307717
rect 327172 307751 327224 307760
rect 327172 307717 327181 307751
rect 327181 307717 327215 307751
rect 327215 307717 327224 307751
rect 327172 307708 327224 307717
rect 337200 307751 337252 307760
rect 337200 307717 337209 307751
rect 337209 307717 337243 307751
rect 337243 307717 337252 307751
rect 337200 307708 337252 307717
rect 374460 307708 374512 307760
rect 301044 306348 301096 306400
rect 301228 306348 301280 306400
rect 317512 306348 317564 306400
rect 317696 306348 317748 306400
rect 463700 306348 463752 306400
rect 463884 306348 463936 306400
rect 580080 306348 580132 306400
rect 580908 306348 580960 306400
rect 294236 304240 294288 304292
rect 294420 304240 294472 304292
rect 338856 302200 338908 302252
rect 338948 302064 339000 302116
rect 377128 302064 377180 302116
rect 377312 302064 377364 302116
rect 236276 299591 236328 299600
rect 236276 299557 236285 299591
rect 236285 299557 236319 299591
rect 236319 299557 236328 299591
rect 236276 299548 236328 299557
rect 259644 299591 259696 299600
rect 259644 299557 259653 299591
rect 259653 299557 259687 299591
rect 259687 299557 259696 299591
rect 259644 299548 259696 299557
rect 267832 299548 267884 299600
rect 288624 299480 288676 299532
rect 288808 299480 288860 299532
rect 299848 299480 299900 299532
rect 306748 299480 306800 299532
rect 306840 299480 306892 299532
rect 341156 299523 341208 299532
rect 341156 299489 341165 299523
rect 341165 299489 341199 299523
rect 341199 299489 341208 299523
rect 341156 299480 341208 299489
rect 357900 299480 357952 299532
rect 358728 299523 358780 299532
rect 358728 299489 358737 299523
rect 358737 299489 358771 299523
rect 358771 299489 358780 299523
rect 358728 299480 358780 299489
rect 389272 299523 389324 299532
rect 389272 299489 389281 299523
rect 389281 299489 389315 299523
rect 389315 299489 389324 299523
rect 389272 299480 389324 299489
rect 470600 299523 470652 299532
rect 470600 299489 470609 299523
rect 470609 299489 470643 299523
rect 470643 299489 470652 299523
rect 470600 299480 470652 299489
rect 235080 299412 235132 299464
rect 235172 299412 235224 299464
rect 236276 299455 236328 299464
rect 236276 299421 236285 299455
rect 236285 299421 236319 299455
rect 236319 299421 236328 299455
rect 236276 299412 236328 299421
rect 259644 299412 259696 299464
rect 259828 299412 259880 299464
rect 267740 299412 267792 299464
rect 323308 299455 323360 299464
rect 323308 299421 323317 299455
rect 323317 299421 323351 299455
rect 323351 299421 323360 299455
rect 323308 299412 323360 299421
rect 324688 299455 324740 299464
rect 324688 299421 324697 299455
rect 324697 299421 324731 299455
rect 324731 299421 324740 299455
rect 324688 299412 324740 299421
rect 325884 299412 325936 299464
rect 338948 299412 339000 299464
rect 372712 299455 372764 299464
rect 372712 299421 372721 299455
rect 372721 299421 372755 299455
rect 372755 299421 372764 299455
rect 372712 299412 372764 299421
rect 375932 299412 375984 299464
rect 469956 299412 470008 299464
rect 580172 299412 580224 299464
rect 325976 299344 326028 299396
rect 338856 299344 338908 299396
rect 262588 298231 262640 298240
rect 262588 298197 262597 298231
rect 262597 298197 262631 298231
rect 262631 298197 262640 298231
rect 262588 298188 262640 298197
rect 310888 298120 310940 298172
rect 327264 298120 327316 298172
rect 330116 298120 330168 298172
rect 330208 298120 330260 298172
rect 337292 298120 337344 298172
rect 262588 298052 262640 298104
rect 266728 298095 266780 298104
rect 266728 298061 266737 298095
rect 266737 298061 266771 298095
rect 266771 298061 266780 298095
rect 266728 298052 266780 298061
rect 267740 298095 267792 298104
rect 267740 298061 267749 298095
rect 267749 298061 267783 298095
rect 267783 298061 267792 298095
rect 267740 298052 267792 298061
rect 285956 298095 286008 298104
rect 285956 298061 285965 298095
rect 285965 298061 285999 298095
rect 285999 298061 286008 298095
rect 285956 298052 286008 298061
rect 325976 298052 326028 298104
rect 326068 298052 326120 298104
rect 358728 298095 358780 298104
rect 358728 298061 358737 298095
rect 358737 298061 358771 298095
rect 358771 298061 358780 298095
rect 358728 298052 358780 298061
rect 262588 297916 262640 297968
rect 301044 296760 301096 296812
rect 301412 296760 301464 296812
rect 580080 296760 580132 296812
rect 581000 296760 581052 296812
rect 284760 296692 284812 296744
rect 284852 296692 284904 296744
rect 299848 296624 299900 296676
rect 299940 296624 299992 296676
rect 301044 296624 301096 296676
rect 301136 296624 301188 296676
rect 306840 296624 306892 296676
rect 306932 296624 306984 296676
rect 580172 296624 580224 296676
rect 581000 296624 581052 296676
rect 272340 295400 272392 295452
rect 272248 295264 272300 295316
rect 302516 295264 302568 295316
rect 302700 295264 302752 295316
rect 251548 294652 251600 294704
rect 290004 294584 290056 294636
rect 290188 294584 290240 294636
rect 310888 293063 310940 293072
rect 310888 293029 310897 293063
rect 310897 293029 310931 293063
rect 310931 293029 310940 293063
rect 310888 293020 310940 293029
rect 377128 292612 377180 292664
rect 239220 292587 239272 292596
rect 239220 292553 239229 292587
rect 239229 292553 239263 292587
rect 239263 292553 239272 292587
rect 239220 292544 239272 292553
rect 288716 292544 288768 292596
rect 295524 292544 295576 292596
rect 296812 292544 296864 292596
rect 337108 292544 337160 292596
rect 337292 292544 337344 292596
rect 357440 292544 357492 292596
rect 357900 292544 357952 292596
rect 270776 292519 270828 292528
rect 270776 292485 270785 292519
rect 270785 292485 270819 292519
rect 270819 292485 270828 292519
rect 270776 292476 270828 292485
rect 288808 292476 288860 292528
rect 295616 292476 295668 292528
rect 296904 292476 296956 292528
rect 377128 292408 377180 292460
rect 236276 289867 236328 289876
rect 236276 289833 236285 289867
rect 236285 289833 236319 289867
rect 236319 289833 236328 289867
rect 236276 289824 236328 289833
rect 239220 289867 239272 289876
rect 239220 289833 239229 289867
rect 239229 289833 239263 289867
rect 239263 289833 239272 289867
rect 239220 289824 239272 289833
rect 251456 289867 251508 289876
rect 251456 289833 251465 289867
rect 251465 289833 251499 289867
rect 251499 289833 251508 289867
rect 251456 289824 251508 289833
rect 294328 289824 294380 289876
rect 324688 289867 324740 289876
rect 324688 289833 324697 289867
rect 324697 289833 324731 289867
rect 324731 289833 324740 289867
rect 324688 289824 324740 289833
rect 372712 289867 372764 289876
rect 372712 289833 372721 289867
rect 372721 289833 372755 289867
rect 372755 289833 372764 289867
rect 372712 289824 372764 289833
rect 374368 289867 374420 289876
rect 374368 289833 374377 289867
rect 374377 289833 374411 289867
rect 374411 289833 374420 289867
rect 374368 289824 374420 289833
rect 375840 289867 375892 289876
rect 375840 289833 375849 289867
rect 375849 289833 375883 289867
rect 375883 289833 375892 289867
rect 375840 289824 375892 289833
rect 244464 289799 244516 289808
rect 244464 289765 244473 289799
rect 244473 289765 244507 289799
rect 244507 289765 244516 289799
rect 244464 289756 244516 289765
rect 250076 289756 250128 289808
rect 250352 289756 250404 289808
rect 259736 289756 259788 289808
rect 259920 289756 259972 289808
rect 290004 289756 290056 289808
rect 290188 289756 290240 289808
rect 327264 289756 327316 289808
rect 357440 289799 357492 289808
rect 357440 289765 357449 289799
rect 357449 289765 357483 289799
rect 357483 289765 357492 289799
rect 357440 289756 357492 289765
rect 389456 289756 389508 289808
rect 470600 289799 470652 289808
rect 470600 289765 470609 289799
rect 470609 289765 470643 289799
rect 470643 289765 470652 289799
rect 470600 289756 470652 289765
rect 236276 289731 236328 289740
rect 236276 289697 236285 289731
rect 236285 289697 236319 289731
rect 236319 289697 236328 289731
rect 236276 289688 236328 289697
rect 266728 288439 266780 288448
rect 266728 288405 266737 288439
rect 266737 288405 266771 288439
rect 266771 288405 266780 288439
rect 266728 288396 266780 288405
rect 267740 288439 267792 288448
rect 267740 288405 267749 288439
rect 267749 288405 267783 288439
rect 267783 288405 267792 288439
rect 267740 288396 267792 288405
rect 285956 288439 286008 288448
rect 285956 288405 285965 288439
rect 285965 288405 285999 288439
rect 285999 288405 286008 288439
rect 285956 288396 286008 288405
rect 323308 288439 323360 288448
rect 323308 288405 323317 288439
rect 323317 288405 323351 288439
rect 323351 288405 323360 288439
rect 323308 288396 323360 288405
rect 358728 288439 358780 288448
rect 358728 288405 358737 288439
rect 358737 288405 358771 288439
rect 358771 288405 358780 288439
rect 358728 288396 358780 288405
rect 291568 287036 291620 287088
rect 291660 287036 291712 287088
rect 294236 287079 294288 287088
rect 294236 287045 294245 287079
rect 294245 287045 294279 287079
rect 294279 287045 294288 287079
rect 294236 287036 294288 287045
rect 330484 287036 330536 287088
rect 330668 287036 330720 287088
rect 463700 287036 463752 287088
rect 463884 287036 463936 287088
rect 580172 287036 580224 287088
rect 580908 287036 580960 287088
rect 270776 285651 270828 285660
rect 270776 285617 270785 285651
rect 270785 285617 270819 285651
rect 270819 285617 270828 285651
rect 270776 285608 270828 285617
rect 337292 285608 337344 285660
rect 284392 283568 284444 283620
rect 284852 283568 284904 283620
rect 323400 283568 323452 283620
rect 327264 283568 327316 283620
rect 296904 282956 296956 283008
rect 341156 282931 341208 282940
rect 341156 282897 341165 282931
rect 341165 282897 341199 282931
rect 341199 282897 341208 282931
rect 341156 282888 341208 282897
rect 360292 282888 360344 282940
rect 360476 282888 360528 282940
rect 296812 282820 296864 282872
rect 310888 282795 310940 282804
rect 310888 282761 310897 282795
rect 310897 282761 310931 282795
rect 310931 282761 310940 282795
rect 310888 282752 310940 282761
rect 358728 280304 358780 280356
rect 236276 280279 236328 280288
rect 236276 280245 236285 280279
rect 236285 280245 236319 280279
rect 236319 280245 236328 280279
rect 236276 280236 236328 280245
rect 244464 280211 244516 280220
rect 244464 280177 244473 280211
rect 244473 280177 244507 280211
rect 244507 280177 244516 280211
rect 244464 280168 244516 280177
rect 265256 280168 265308 280220
rect 295524 280168 295576 280220
rect 295616 280168 295668 280220
rect 341156 280211 341208 280220
rect 341156 280177 341165 280211
rect 341165 280177 341199 280211
rect 341199 280177 341208 280211
rect 341156 280168 341208 280177
rect 357716 280168 357768 280220
rect 358728 280168 358780 280220
rect 389364 280211 389416 280220
rect 389364 280177 389373 280211
rect 389373 280177 389407 280211
rect 389407 280177 389416 280211
rect 389364 280168 389416 280177
rect 470600 280211 470652 280220
rect 470600 280177 470609 280211
rect 470609 280177 470643 280211
rect 470643 280177 470652 280211
rect 470600 280168 470652 280177
rect 235080 280100 235132 280152
rect 235172 280100 235224 280152
rect 236276 280143 236328 280152
rect 236276 280109 236285 280143
rect 236285 280109 236319 280143
rect 236319 280109 236328 280143
rect 236276 280100 236328 280109
rect 239128 280143 239180 280152
rect 239128 280109 239137 280143
rect 239137 280109 239171 280143
rect 239171 280109 239180 280143
rect 239128 280100 239180 280109
rect 251456 280143 251508 280152
rect 251456 280109 251465 280143
rect 251465 280109 251499 280143
rect 251499 280109 251508 280143
rect 251456 280100 251508 280109
rect 259552 280143 259604 280152
rect 259552 280109 259561 280143
rect 259561 280109 259595 280143
rect 259595 280109 259604 280143
rect 259552 280100 259604 280109
rect 273536 280100 273588 280152
rect 273628 280100 273680 280152
rect 285956 280100 286008 280152
rect 286140 280100 286192 280152
rect 288624 280100 288676 280152
rect 288808 280100 288860 280152
rect 331404 280143 331456 280152
rect 331404 280109 331413 280143
rect 331413 280109 331447 280143
rect 331447 280109 331456 280143
rect 331404 280100 331456 280109
rect 338856 280143 338908 280152
rect 338856 280109 338865 280143
rect 338865 280109 338899 280143
rect 338899 280109 338908 280143
rect 338856 280100 338908 280109
rect 372712 280143 372764 280152
rect 372712 280109 372721 280143
rect 372721 280109 372755 280143
rect 372755 280109 372764 280143
rect 372712 280100 372764 280109
rect 377128 280143 377180 280152
rect 377128 280109 377137 280143
rect 377137 280109 377171 280143
rect 377171 280109 377180 280143
rect 377128 280100 377180 280109
rect 265256 280032 265308 280084
rect 291568 278808 291620 278860
rect 291752 278808 291804 278860
rect 250076 278740 250128 278792
rect 250168 278740 250220 278792
rect 301044 278740 301096 278792
rect 301228 278740 301280 278792
rect 302516 278740 302568 278792
rect 323492 278783 323544 278792
rect 323492 278749 323501 278783
rect 323501 278749 323535 278783
rect 323535 278749 323544 278783
rect 323492 278740 323544 278749
rect 330208 278740 330260 278792
rect 330484 278740 330536 278792
rect 302608 278672 302660 278724
rect 310888 278715 310940 278724
rect 310888 278681 310897 278715
rect 310897 278681 310931 278715
rect 310931 278681 310940 278715
rect 310888 278672 310940 278681
rect 294236 277380 294288 277432
rect 294328 277380 294380 277432
rect 580172 277312 580224 277364
rect 580908 277312 580960 277364
rect 337200 276063 337252 276072
rect 337200 276029 337209 276063
rect 337209 276029 337243 276063
rect 337243 276029 337252 276063
rect 337200 276020 337252 276029
rect 302608 275952 302660 276004
rect 302792 275952 302844 276004
rect 306656 275952 306708 276004
rect 306932 275952 306984 276004
rect 284392 273912 284444 273964
rect 284760 273912 284812 273964
rect 330116 273887 330168 273896
rect 330116 273853 330125 273887
rect 330125 273853 330159 273887
rect 330159 273853 330168 273887
rect 330116 273844 330168 273853
rect 250168 273300 250220 273352
rect 301044 273232 301096 273284
rect 357440 273232 357492 273284
rect 357716 273232 357768 273284
rect 250076 273164 250128 273216
rect 301136 273164 301188 273216
rect 374368 273164 374420 273216
rect 375840 273164 375892 273216
rect 259552 273071 259604 273080
rect 259552 273037 259561 273071
rect 259561 273037 259595 273071
rect 259595 273037 259604 273071
rect 259552 273028 259604 273037
rect 374368 273028 374420 273080
rect 375840 273028 375892 273080
rect 299940 270580 299992 270632
rect 236276 270555 236328 270564
rect 236276 270521 236285 270555
rect 236285 270521 236319 270555
rect 236319 270521 236328 270555
rect 236276 270512 236328 270521
rect 239220 270512 239272 270564
rect 251456 270555 251508 270564
rect 251456 270521 251465 270555
rect 251465 270521 251499 270555
rect 251499 270521 251508 270555
rect 251456 270512 251508 270521
rect 262496 270512 262548 270564
rect 262680 270512 262732 270564
rect 267740 270512 267792 270564
rect 267832 270512 267884 270564
rect 299756 270512 299808 270564
rect 331404 270555 331456 270564
rect 331404 270521 331413 270555
rect 331413 270521 331447 270555
rect 331447 270521 331456 270555
rect 331404 270512 331456 270521
rect 338856 270555 338908 270564
rect 338856 270521 338865 270555
rect 338865 270521 338899 270555
rect 338899 270521 338908 270555
rect 338856 270512 338908 270521
rect 372712 270555 372764 270564
rect 372712 270521 372721 270555
rect 372721 270521 372755 270555
rect 372755 270521 372764 270555
rect 372712 270512 372764 270521
rect 377128 270555 377180 270564
rect 377128 270521 377137 270555
rect 377137 270521 377171 270555
rect 377171 270521 377180 270555
rect 377128 270512 377180 270521
rect 325976 270444 326028 270496
rect 326068 270444 326120 270496
rect 341248 270444 341300 270496
rect 341432 270444 341484 270496
rect 389456 270444 389508 270496
rect 470600 270487 470652 270496
rect 470600 270453 470609 270487
rect 470609 270453 470643 270487
rect 470643 270453 470652 270487
rect 470600 270444 470652 270453
rect 236276 270419 236328 270428
rect 236276 270385 236285 270419
rect 236285 270385 236319 270419
rect 236319 270385 236328 270419
rect 236276 270376 236328 270385
rect 290096 269084 290148 269136
rect 290188 269084 290240 269136
rect 291752 269152 291804 269204
rect 296812 269084 296864 269136
rect 297088 269084 297140 269136
rect 324596 269084 324648 269136
rect 324780 269084 324832 269136
rect 330208 269084 330260 269136
rect 358544 269084 358596 269136
rect 358728 269084 358780 269136
rect 250076 269059 250128 269068
rect 250076 269025 250085 269059
rect 250085 269025 250119 269059
rect 250119 269025 250128 269059
rect 250076 269016 250128 269025
rect 291568 269016 291620 269068
rect 265256 267724 265308 267776
rect 265440 267724 265492 267776
rect 294144 267724 294196 267776
rect 294328 267724 294380 267776
rect 295524 267724 295576 267776
rect 295800 267724 295852 267776
rect 463700 267724 463752 267776
rect 463884 267724 463936 267776
rect 337016 266296 337068 266348
rect 337200 266296 337252 266348
rect 270684 263576 270736 263628
rect 327264 263644 327316 263696
rect 360292 263576 360344 263628
rect 360476 263576 360528 263628
rect 327172 263508 327224 263560
rect 270684 263440 270736 263492
rect 310888 263483 310940 263492
rect 310888 263449 310897 263483
rect 310897 263449 310931 263483
rect 310931 263449 310940 263483
rect 310888 263440 310940 263449
rect 296812 262896 296864 262948
rect 296996 262896 297048 262948
rect 236276 260967 236328 260976
rect 236276 260933 236285 260967
rect 236285 260933 236319 260967
rect 236319 260933 236328 260967
rect 236276 260924 236328 260933
rect 323400 260924 323452 260976
rect 323492 260924 323544 260976
rect 262588 260899 262640 260908
rect 262588 260865 262597 260899
rect 262597 260865 262631 260899
rect 262631 260865 262640 260899
rect 262588 260856 262640 260865
rect 266636 260856 266688 260908
rect 266728 260856 266780 260908
rect 288624 260856 288676 260908
rect 288808 260856 288860 260908
rect 295708 260856 295760 260908
rect 389364 260899 389416 260908
rect 389364 260865 389373 260899
rect 389373 260865 389407 260899
rect 389407 260865 389416 260899
rect 389364 260856 389416 260865
rect 470600 260899 470652 260908
rect 470600 260865 470609 260899
rect 470609 260865 470643 260899
rect 470643 260865 470652 260899
rect 470600 260856 470652 260865
rect 235080 260788 235132 260840
rect 235172 260788 235224 260840
rect 236276 260831 236328 260840
rect 236276 260797 236285 260831
rect 236285 260797 236319 260831
rect 236319 260797 236328 260831
rect 236276 260788 236328 260797
rect 239128 260831 239180 260840
rect 239128 260797 239137 260831
rect 239137 260797 239171 260831
rect 239171 260797 239180 260831
rect 239128 260788 239180 260797
rect 251456 260831 251508 260840
rect 251456 260797 251465 260831
rect 251465 260797 251499 260831
rect 251499 260797 251508 260831
rect 251456 260788 251508 260797
rect 259552 260831 259604 260840
rect 259552 260797 259561 260831
rect 259561 260797 259595 260831
rect 259595 260797 259604 260831
rect 259552 260788 259604 260797
rect 270684 260831 270736 260840
rect 270684 260797 270693 260831
rect 270693 260797 270727 260831
rect 270727 260797 270736 260831
rect 270684 260788 270736 260797
rect 272156 260788 272208 260840
rect 273536 260788 273588 260840
rect 273628 260788 273680 260840
rect 295800 260788 295852 260840
rect 324596 260788 324648 260840
rect 338856 260831 338908 260840
rect 338856 260797 338865 260831
rect 338865 260797 338899 260831
rect 338899 260797 338908 260831
rect 338856 260788 338908 260797
rect 341064 260831 341116 260840
rect 341064 260797 341073 260831
rect 341073 260797 341107 260831
rect 341107 260797 341116 260831
rect 341064 260788 341116 260797
rect 372712 260831 372764 260840
rect 372712 260797 372721 260831
rect 372721 260797 372755 260831
rect 372755 260797 372764 260831
rect 372712 260788 372764 260797
rect 377128 260831 377180 260840
rect 377128 260797 377137 260831
rect 377137 260797 377171 260831
rect 377171 260797 377180 260831
rect 377128 260788 377180 260797
rect 463792 260788 463844 260840
rect 324688 260720 324740 260772
rect 272156 260652 272208 260704
rect 250168 259428 250220 259480
rect 262588 259471 262640 259480
rect 262588 259437 262597 259471
rect 262597 259437 262631 259471
rect 262631 259437 262640 259471
rect 262588 259428 262640 259437
rect 267740 259428 267792 259480
rect 267832 259428 267884 259480
rect 284576 259428 284628 259480
rect 284760 259428 284812 259480
rect 330116 259428 330168 259480
rect 330392 259428 330444 259480
rect 324688 259360 324740 259412
rect 324780 259360 324832 259412
rect 357532 259403 357584 259412
rect 357532 259369 357541 259403
rect 357541 259369 357575 259403
rect 357575 259369 357584 259403
rect 357532 259360 357584 259369
rect 250168 259335 250220 259344
rect 250168 259301 250177 259335
rect 250177 259301 250211 259335
rect 250211 259301 250220 259335
rect 250168 259292 250220 259301
rect 264980 258000 265032 258052
rect 265348 258000 265400 258052
rect 267924 258000 267976 258052
rect 268108 258000 268160 258052
rect 301228 258000 301280 258052
rect 301412 258000 301464 258052
rect 306840 258000 306892 258052
rect 330116 258000 330168 258052
rect 330300 258000 330352 258052
rect 310888 256071 310940 256080
rect 310888 256037 310897 256071
rect 310897 256037 310931 256071
rect 310931 256037 310940 256071
rect 310888 256028 310940 256037
rect 337200 253988 337252 254040
rect 374368 253852 374420 253904
rect 375840 253852 375892 253904
rect 259552 253759 259604 253768
rect 259552 253725 259561 253759
rect 259561 253725 259595 253759
rect 259595 253725 259604 253759
rect 259552 253716 259604 253725
rect 341064 253759 341116 253768
rect 341064 253725 341073 253759
rect 341073 253725 341107 253759
rect 341107 253725 341116 253759
rect 341064 253716 341116 253725
rect 374368 253716 374420 253768
rect 375840 253716 375892 253768
rect 295248 253172 295300 253224
rect 295616 253172 295668 253224
rect 469864 252492 469916 252544
rect 579620 252492 579672 252544
rect 2780 252016 2832 252068
rect 5356 252016 5408 252068
rect 310704 251268 310756 251320
rect 236276 251243 236328 251252
rect 236276 251209 236285 251243
rect 236285 251209 236319 251243
rect 236319 251209 236328 251243
rect 236276 251200 236328 251209
rect 239220 251200 239272 251252
rect 251456 251243 251508 251252
rect 251456 251209 251465 251243
rect 251465 251209 251499 251243
rect 251499 251209 251508 251243
rect 251456 251200 251508 251209
rect 290004 251200 290056 251252
rect 290096 251200 290148 251252
rect 327172 251200 327224 251252
rect 327264 251200 327316 251252
rect 338856 251243 338908 251252
rect 338856 251209 338865 251243
rect 338865 251209 338899 251243
rect 338899 251209 338908 251243
rect 338856 251200 338908 251209
rect 372712 251243 372764 251252
rect 372712 251209 372721 251243
rect 372721 251209 372755 251243
rect 372755 251209 372764 251243
rect 372712 251200 372764 251209
rect 377128 251243 377180 251252
rect 377128 251209 377137 251243
rect 377137 251209 377171 251243
rect 377171 251209 377180 251243
rect 377128 251200 377180 251209
rect 389180 251200 389232 251252
rect 389364 251200 389416 251252
rect 463700 251243 463752 251252
rect 463700 251209 463709 251243
rect 463709 251209 463743 251243
rect 463743 251209 463752 251243
rect 463700 251200 463752 251209
rect 259552 251175 259604 251184
rect 259552 251141 259561 251175
rect 259561 251141 259595 251175
rect 259595 251141 259604 251175
rect 259552 251132 259604 251141
rect 310704 251175 310756 251184
rect 310704 251141 310713 251175
rect 310713 251141 310747 251175
rect 310747 251141 310756 251175
rect 310704 251132 310756 251141
rect 325976 251132 326028 251184
rect 326068 251132 326120 251184
rect 470600 251175 470652 251184
rect 470600 251141 470609 251175
rect 470609 251141 470643 251175
rect 470643 251141 470652 251175
rect 470600 251132 470652 251141
rect 250352 251064 250404 251116
rect 270776 251064 270828 251116
rect 284668 249840 284720 249892
rect 284760 249840 284812 249892
rect 285956 249772 286008 249824
rect 286048 249772 286100 249824
rect 302700 249772 302752 249824
rect 302792 249772 302844 249824
rect 323216 249772 323268 249824
rect 323492 249772 323544 249824
rect 357716 249772 357768 249824
rect 358544 249772 358596 249824
rect 358728 249772 358780 249824
rect 290004 249704 290056 249756
rect 290188 249704 290240 249756
rect 296904 248412 296956 248464
rect 296996 248412 297048 248464
rect 295524 248344 295576 248396
rect 295800 248344 295852 248396
rect 306748 248387 306800 248396
rect 306748 248353 306757 248387
rect 306757 248353 306791 248387
rect 306791 248353 306800 248387
rect 306748 248344 306800 248353
rect 337108 247163 337160 247172
rect 337108 247129 337117 247163
rect 337117 247129 337151 247163
rect 337151 247129 337160 247163
rect 337108 247120 337160 247129
rect 337108 247027 337160 247036
rect 337108 246993 337117 247027
rect 337117 246993 337151 247027
rect 337151 246993 337160 247027
rect 337108 246984 337160 246993
rect 285956 244987 286008 244996
rect 285956 244953 285965 244987
rect 285965 244953 285999 244987
rect 285999 244953 286008 244987
rect 285956 244944 286008 244953
rect 272156 244443 272208 244452
rect 272156 244409 272165 244443
rect 272165 244409 272199 244443
rect 272199 244409 272208 244443
rect 272156 244400 272208 244409
rect 360292 244264 360344 244316
rect 360476 244264 360528 244316
rect 329932 244196 329984 244248
rect 330208 244196 330260 244248
rect 337108 244239 337160 244248
rect 337108 244205 337117 244239
rect 337117 244205 337151 244239
rect 337151 244205 337160 244239
rect 337108 244196 337160 244205
rect 259644 244128 259696 244180
rect 262680 241544 262732 241596
rect 236276 241476 236328 241528
rect 236460 241476 236512 241528
rect 262588 241476 262640 241528
rect 266636 241476 266688 241528
rect 266728 241476 266780 241528
rect 270776 241544 270828 241596
rect 272156 241587 272208 241596
rect 272156 241553 272165 241587
rect 272165 241553 272199 241587
rect 272199 241553 272208 241587
rect 272156 241544 272208 241553
rect 323492 241544 323544 241596
rect 388996 241544 389048 241596
rect 389272 241544 389324 241596
rect 310888 241476 310940 241528
rect 323400 241476 323452 241528
rect 470600 241519 470652 241528
rect 470600 241485 470609 241519
rect 470609 241485 470643 241519
rect 470643 241485 470652 241519
rect 470600 241476 470652 241485
rect 270684 241408 270736 241460
rect 299480 241451 299532 241460
rect 299480 241417 299489 241451
rect 299489 241417 299523 241451
rect 299523 241417 299532 241451
rect 331404 241451 331456 241460
rect 299480 241408 299532 241417
rect 331404 241417 331413 241451
rect 331413 241417 331447 241451
rect 331447 241417 331456 241451
rect 331404 241408 331456 241417
rect 389272 241451 389324 241460
rect 389272 241417 389281 241451
rect 389281 241417 389315 241451
rect 389315 241417 389324 241451
rect 389272 241408 389324 241417
rect 259644 241340 259696 241392
rect 259828 241340 259880 241392
rect 284760 240116 284812 240168
rect 284944 240116 284996 240168
rect 301320 240184 301372 240236
rect 267740 240091 267792 240100
rect 267740 240057 267749 240091
rect 267749 240057 267783 240091
rect 267783 240057 267792 240091
rect 267740 240048 267792 240057
rect 272156 240091 272208 240100
rect 272156 240057 272165 240091
rect 272165 240057 272199 240091
rect 272199 240057 272208 240091
rect 272156 240048 272208 240057
rect 273536 240048 273588 240100
rect 273628 240048 273680 240100
rect 294328 240048 294380 240100
rect 294420 240048 294472 240100
rect 301044 240048 301096 240100
rect 306748 238756 306800 238808
rect 290372 238731 290424 238740
rect 290372 238697 290381 238731
rect 290381 238697 290415 238731
rect 290415 238697 290424 238731
rect 290372 238688 290424 238697
rect 295616 238731 295668 238740
rect 295616 238697 295625 238731
rect 295625 238697 295659 238731
rect 295659 238697 295668 238731
rect 295616 238688 295668 238697
rect 3056 237328 3108 237380
rect 15844 237328 15896 237380
rect 266728 234855 266780 234864
rect 266728 234821 266737 234855
rect 266737 234821 266771 234855
rect 266771 234821 266780 234855
rect 266728 234812 266780 234821
rect 265164 234608 265216 234660
rect 310888 234676 310940 234728
rect 389456 234608 389508 234660
rect 310796 234540 310848 234592
rect 374368 234540 374420 234592
rect 375840 234540 375892 234592
rect 265256 234472 265308 234524
rect 272248 234472 272300 234524
rect 285956 234515 286008 234524
rect 285956 234481 285965 234515
rect 285965 234481 285999 234515
rect 285999 234481 286008 234515
rect 285956 234472 286008 234481
rect 374368 234404 374420 234456
rect 375840 234404 375892 234456
rect 235080 231820 235132 231872
rect 235172 231820 235224 231872
rect 244280 231820 244332 231872
rect 244464 231820 244516 231872
rect 250076 231820 250128 231872
rect 250352 231820 250404 231872
rect 251456 231820 251508 231872
rect 251640 231820 251692 231872
rect 299480 231863 299532 231872
rect 299480 231829 299489 231863
rect 299489 231829 299523 231863
rect 299523 231829 299532 231863
rect 299480 231820 299532 231829
rect 323308 231820 323360 231872
rect 323492 231820 323544 231872
rect 324688 231820 324740 231872
rect 324780 231820 324832 231872
rect 331404 231863 331456 231872
rect 331404 231829 331413 231863
rect 331413 231829 331447 231863
rect 331447 231829 331456 231863
rect 331404 231820 331456 231829
rect 338672 231820 338724 231872
rect 338856 231820 338908 231872
rect 341064 231820 341116 231872
rect 341156 231820 341208 231872
rect 372528 231820 372580 231872
rect 372712 231820 372764 231872
rect 376944 231820 376996 231872
rect 377128 231820 377180 231872
rect 267924 231752 267976 231804
rect 310796 231795 310848 231804
rect 310796 231761 310805 231795
rect 310805 231761 310839 231795
rect 310839 231761 310848 231795
rect 310796 231752 310848 231761
rect 337200 231616 337252 231668
rect 266728 230503 266780 230512
rect 266728 230469 266737 230503
rect 266737 230469 266771 230503
rect 266771 230469 266780 230503
rect 266728 230460 266780 230469
rect 301044 230460 301096 230512
rect 301228 230460 301280 230512
rect 306840 230460 306892 230512
rect 327172 230460 327224 230512
rect 327356 230460 327408 230512
rect 358544 230460 358596 230512
rect 358728 230460 358780 230512
rect 290372 230435 290424 230444
rect 290372 230401 290381 230435
rect 290381 230401 290415 230435
rect 290415 230401 290424 230435
rect 290372 230392 290424 230401
rect 295616 229143 295668 229152
rect 295616 229109 295625 229143
rect 295625 229109 295659 229143
rect 295659 229109 295668 229143
rect 295616 229100 295668 229109
rect 270684 224995 270736 225004
rect 270684 224961 270693 224995
rect 270693 224961 270727 224995
rect 270727 224961 270736 224995
rect 270684 224952 270736 224961
rect 341156 224952 341208 225004
rect 360292 224952 360344 225004
rect 360476 224952 360528 225004
rect 236276 222164 236328 222216
rect 236460 222164 236512 222216
rect 259644 222164 259696 222216
rect 259828 222164 259880 222216
rect 262680 222164 262732 222216
rect 262772 222164 262824 222216
rect 265164 222164 265216 222216
rect 265348 222164 265400 222216
rect 284760 222164 284812 222216
rect 295524 222164 295576 222216
rect 295616 222164 295668 222216
rect 301228 222232 301280 222284
rect 302516 222164 302568 222216
rect 302700 222164 302752 222216
rect 310888 222164 310940 222216
rect 324688 222164 324740 222216
rect 324780 222164 324832 222216
rect 341064 222207 341116 222216
rect 341064 222173 341073 222207
rect 341073 222173 341107 222207
rect 341107 222173 341116 222207
rect 341064 222164 341116 222173
rect 389272 222164 389324 222216
rect 389548 222164 389600 222216
rect 463792 222164 463844 222216
rect 464068 222164 464120 222216
rect 470416 222164 470468 222216
rect 470600 222164 470652 222216
rect 299480 222139 299532 222148
rect 299480 222105 299489 222139
rect 299489 222105 299523 222139
rect 299523 222105 299532 222139
rect 299480 222096 299532 222105
rect 301044 222096 301096 222148
rect 259644 222028 259696 222080
rect 259828 222028 259880 222080
rect 284760 222028 284812 222080
rect 270684 220847 270736 220856
rect 270684 220813 270693 220847
rect 270693 220813 270727 220847
rect 270727 220813 270736 220847
rect 270684 220804 270736 220813
rect 288900 220804 288952 220856
rect 289084 220804 289136 220856
rect 290188 220804 290240 220856
rect 290372 220804 290424 220856
rect 291660 220804 291712 220856
rect 291936 220804 291988 220856
rect 294328 220804 294380 220856
rect 294420 220804 294472 220856
rect 337292 220804 337344 220856
rect 290188 219419 290240 219428
rect 290188 219385 290197 219419
rect 290197 219385 290231 219419
rect 290231 219385 290240 219419
rect 290188 219376 290240 219385
rect 291660 219419 291712 219428
rect 291660 219385 291669 219419
rect 291669 219385 291703 219419
rect 291703 219385 291712 219419
rect 291660 219376 291712 219385
rect 317512 219376 317564 219428
rect 317696 219376 317748 219428
rect 310888 215364 310940 215416
rect 389548 215364 389600 215416
rect 464068 215364 464120 215416
rect 273444 215228 273496 215280
rect 273628 215228 273680 215280
rect 310796 215228 310848 215280
rect 374368 215228 374420 215280
rect 375840 215228 375892 215280
rect 389456 215228 389508 215280
rect 463976 215228 464028 215280
rect 374368 215092 374420 215144
rect 375840 215092 375892 215144
rect 235080 212508 235132 212560
rect 235172 212508 235224 212560
rect 244280 212508 244332 212560
rect 244464 212508 244516 212560
rect 250076 212508 250128 212560
rect 250352 212508 250404 212560
rect 251456 212508 251508 212560
rect 251640 212508 251692 212560
rect 265164 212508 265216 212560
rect 265256 212508 265308 212560
rect 266636 212508 266688 212560
rect 266820 212508 266872 212560
rect 267832 212508 267884 212560
rect 267924 212508 267976 212560
rect 284760 212508 284812 212560
rect 299480 212551 299532 212560
rect 299480 212517 299489 212551
rect 299489 212517 299523 212551
rect 299523 212517 299532 212551
rect 299480 212508 299532 212517
rect 323308 212508 323360 212560
rect 323492 212508 323544 212560
rect 324688 212508 324740 212560
rect 324780 212508 324832 212560
rect 331404 212508 331456 212560
rect 331588 212508 331640 212560
rect 337292 212576 337344 212628
rect 338672 212508 338724 212560
rect 338856 212508 338908 212560
rect 372528 212508 372580 212560
rect 372712 212508 372764 212560
rect 376944 212508 376996 212560
rect 377128 212508 377180 212560
rect 284944 212440 284996 212492
rect 290188 212483 290240 212492
rect 290188 212449 290197 212483
rect 290197 212449 290231 212483
rect 290231 212449 290240 212483
rect 290188 212440 290240 212449
rect 291660 212483 291712 212492
rect 291660 212449 291669 212483
rect 291669 212449 291703 212483
rect 291703 212449 291712 212483
rect 291660 212440 291712 212449
rect 310796 212483 310848 212492
rect 310796 212449 310805 212483
rect 310805 212449 310839 212483
rect 310839 212449 310848 212483
rect 310796 212440 310848 212449
rect 337200 212440 337252 212492
rect 299848 211148 299900 211200
rect 299940 211148 299992 211200
rect 250076 211080 250128 211132
rect 250260 211080 250312 211132
rect 267832 211080 267884 211132
rect 267924 211080 267976 211132
rect 294236 211080 294288 211132
rect 294328 211080 294380 211132
rect 306656 211080 306708 211132
rect 306840 211080 306892 211132
rect 337200 211080 337252 211132
rect 337384 211080 337436 211132
rect 317512 209788 317564 209840
rect 317696 209788 317748 209840
rect 306656 209720 306708 209772
rect 306932 209720 306984 209772
rect 341248 209720 341300 209772
rect 341340 209720 341392 209772
rect 262588 207884 262640 207936
rect 262772 207884 262824 207936
rect 302608 207791 302660 207800
rect 302608 207757 302617 207791
rect 302617 207757 302651 207791
rect 302651 207757 302660 207791
rect 302608 207748 302660 207757
rect 266636 205640 266688 205692
rect 270684 205683 270736 205692
rect 270684 205649 270693 205683
rect 270693 205649 270727 205683
rect 270727 205649 270736 205683
rect 270684 205640 270736 205649
rect 323308 205640 323360 205692
rect 360292 205640 360344 205692
rect 360476 205640 360528 205692
rect 266728 205572 266780 205624
rect 323400 205504 323452 205556
rect 236276 202852 236328 202904
rect 236460 202852 236512 202904
rect 270684 202895 270736 202904
rect 270684 202861 270693 202895
rect 270693 202861 270727 202895
rect 270727 202861 270736 202895
rect 270684 202852 270736 202861
rect 285956 202852 286008 202904
rect 286140 202852 286192 202904
rect 295524 202852 295576 202904
rect 295616 202852 295668 202904
rect 296812 202852 296864 202904
rect 296904 202852 296956 202904
rect 302608 202895 302660 202904
rect 302608 202861 302617 202895
rect 302617 202861 302651 202895
rect 302651 202861 302660 202895
rect 302608 202852 302660 202861
rect 310888 202852 310940 202904
rect 324596 202852 324648 202904
rect 324688 202852 324740 202904
rect 329932 202852 329984 202904
rect 330116 202852 330168 202904
rect 389272 202852 389324 202904
rect 389548 202852 389600 202904
rect 463792 202852 463844 202904
rect 464068 202852 464120 202904
rect 470416 202852 470468 202904
rect 470600 202852 470652 202904
rect 273536 202784 273588 202836
rect 273628 202784 273680 202836
rect 250076 201424 250128 201476
rect 250352 201424 250404 201476
rect 301044 201424 301096 201476
rect 301136 201356 301188 201408
rect 250076 200107 250128 200116
rect 250076 200073 250085 200107
rect 250085 200073 250119 200107
rect 250119 200073 250128 200107
rect 250076 200064 250128 200073
rect 289912 200064 289964 200116
rect 290188 200064 290240 200116
rect 291384 200064 291436 200116
rect 291660 200064 291712 200116
rect 299756 200064 299808 200116
rect 299848 200064 299900 200116
rect 306748 200064 306800 200116
rect 306840 200064 306892 200116
rect 317512 200064 317564 200116
rect 317696 200064 317748 200116
rect 341248 198704 341300 198756
rect 341340 198704 341392 198756
rect 266728 198092 266780 198144
rect 266636 198024 266688 198076
rect 285772 198024 285824 198076
rect 285956 198024 286008 198076
rect 294236 198024 294288 198076
rect 294420 198024 294472 198076
rect 329932 198024 329984 198076
rect 330116 198024 330168 198076
rect 310888 196052 310940 196104
rect 389548 196052 389600 196104
rect 464068 196052 464120 196104
rect 310796 195916 310848 195968
rect 357532 195916 357584 195968
rect 357716 195916 357768 195968
rect 374368 195916 374420 195968
rect 375840 195916 375892 195968
rect 389456 195916 389508 195968
rect 463976 195916 464028 195968
rect 374368 195780 374420 195832
rect 375840 195780 375892 195832
rect 288716 193332 288768 193384
rect 337108 193332 337160 193384
rect 230848 193196 230900 193248
rect 231032 193196 231084 193248
rect 235080 193196 235132 193248
rect 235172 193196 235224 193248
rect 239128 193196 239180 193248
rect 239220 193196 239272 193248
rect 244280 193196 244332 193248
rect 244464 193196 244516 193248
rect 251456 193196 251508 193248
rect 251640 193196 251692 193248
rect 259736 193196 259788 193248
rect 259920 193196 259972 193248
rect 265256 193196 265308 193248
rect 265348 193196 265400 193248
rect 267832 193196 267884 193248
rect 267924 193196 267976 193248
rect 288716 193196 288768 193248
rect 323308 193196 323360 193248
rect 323492 193196 323544 193248
rect 324596 193196 324648 193248
rect 324688 193196 324740 193248
rect 331404 193196 331456 193248
rect 331588 193196 331640 193248
rect 337108 193196 337160 193248
rect 338672 193196 338724 193248
rect 338856 193196 338908 193248
rect 372528 193196 372580 193248
rect 372712 193196 372764 193248
rect 376944 193196 376996 193248
rect 377128 193196 377180 193248
rect 367008 193171 367060 193180
rect 367008 193137 367017 193171
rect 367017 193137 367051 193171
rect 367051 193137 367060 193171
rect 367008 193128 367060 193137
rect 324688 191768 324740 191820
rect 324872 191768 324924 191820
rect 358544 191768 358596 191820
rect 358820 191768 358872 191820
rect 317512 190476 317564 190528
rect 317696 190476 317748 190528
rect 264980 190408 265032 190460
rect 265256 190408 265308 190460
rect 299848 190451 299900 190460
rect 299848 190417 299857 190451
rect 299857 190417 299891 190451
rect 299891 190417 299900 190451
rect 299848 190408 299900 190417
rect 302792 190408 302844 190460
rect 306840 190451 306892 190460
rect 306840 190417 306849 190451
rect 306849 190417 306883 190451
rect 306883 190417 306892 190451
rect 306840 190408 306892 190417
rect 288716 189023 288768 189032
rect 288716 188989 288725 189023
rect 288725 188989 288759 189023
rect 288759 188989 288768 189023
rect 288716 188980 288768 188989
rect 341248 188980 341300 189032
rect 341432 188980 341484 189032
rect 339776 188411 339828 188420
rect 339776 188377 339785 188411
rect 339785 188377 339819 188411
rect 339819 188377 339828 188411
rect 339776 188368 339828 188377
rect 330116 186940 330168 186992
rect 330300 186940 330352 186992
rect 266636 186328 266688 186380
rect 267740 186371 267792 186380
rect 267740 186337 267749 186371
rect 267749 186337 267783 186371
rect 267783 186337 267792 186371
rect 267740 186328 267792 186337
rect 270684 186371 270736 186380
rect 270684 186337 270693 186371
rect 270693 186337 270727 186371
rect 270727 186337 270736 186371
rect 270684 186328 270736 186337
rect 250076 186303 250128 186312
rect 250076 186269 250085 186303
rect 250085 186269 250119 186303
rect 250119 186269 250128 186303
rect 250076 186260 250128 186269
rect 295616 186328 295668 186380
rect 296904 186396 296956 186448
rect 327264 186396 327316 186448
rect 295524 186260 295576 186312
rect 296812 186260 296864 186312
rect 327172 186260 327224 186312
rect 266728 186192 266780 186244
rect 236276 183540 236328 183592
rect 236460 183540 236512 183592
rect 267740 183583 267792 183592
rect 267740 183549 267749 183583
rect 267749 183549 267783 183583
rect 267783 183549 267792 183583
rect 267740 183540 267792 183549
rect 270684 183583 270736 183592
rect 270684 183549 270693 183583
rect 270693 183549 270727 183583
rect 270727 183549 270736 183583
rect 270684 183540 270736 183549
rect 284760 183540 284812 183592
rect 294236 183540 294288 183592
rect 294420 183540 294472 183592
rect 310888 183540 310940 183592
rect 311072 183540 311124 183592
rect 339868 183540 339920 183592
rect 367008 183583 367060 183592
rect 367008 183549 367017 183583
rect 367017 183549 367051 183583
rect 367051 183549 367060 183583
rect 367008 183540 367060 183549
rect 389272 183540 389324 183592
rect 389548 183540 389600 183592
rect 463792 183540 463844 183592
rect 464068 183540 464120 183592
rect 470416 183540 470468 183592
rect 470600 183540 470652 183592
rect 273536 183472 273588 183524
rect 273628 183472 273680 183524
rect 284760 183404 284812 183456
rect 232320 182155 232372 182164
rect 232320 182121 232329 182155
rect 232329 182121 232363 182155
rect 232363 182121 232372 182155
rect 232320 182112 232372 182121
rect 301044 182112 301096 182164
rect 301228 182112 301280 182164
rect 324504 182112 324556 182164
rect 326068 182112 326120 182164
rect 326252 182112 326304 182164
rect 324688 182044 324740 182096
rect 358728 182019 358780 182028
rect 358728 181985 358737 182019
rect 358737 181985 358771 182019
rect 358771 181985 358780 182019
rect 358728 181976 358780 181985
rect 299848 180863 299900 180872
rect 299848 180829 299857 180863
rect 299857 180829 299891 180863
rect 299891 180829 299900 180863
rect 299848 180820 299900 180829
rect 302516 180863 302568 180872
rect 302516 180829 302525 180863
rect 302525 180829 302559 180863
rect 302559 180829 302568 180863
rect 302516 180820 302568 180829
rect 306840 180863 306892 180872
rect 306840 180829 306849 180863
rect 306849 180829 306883 180863
rect 306883 180829 306892 180863
rect 306840 180820 306892 180829
rect 265164 180752 265216 180804
rect 265256 180752 265308 180804
rect 272248 180752 272300 180804
rect 272432 180752 272484 180804
rect 284760 180795 284812 180804
rect 284760 180761 284769 180795
rect 284769 180761 284803 180795
rect 284803 180761 284812 180795
rect 284760 180752 284812 180761
rect 317512 180752 317564 180804
rect 317696 180752 317748 180804
rect 259644 179571 259696 179580
rect 259644 179537 259653 179571
rect 259653 179537 259687 179571
rect 259687 179537 259696 179571
rect 259644 179528 259696 179537
rect 288900 179392 288952 179444
rect 265256 179367 265308 179376
rect 265256 179333 265265 179367
rect 265265 179333 265299 179367
rect 265299 179333 265308 179367
rect 265256 179324 265308 179333
rect 341248 179367 341300 179376
rect 341248 179333 341257 179367
rect 341257 179333 341291 179367
rect 341291 179333 341300 179367
rect 341248 179324 341300 179333
rect 294236 178712 294288 178764
rect 294420 178712 294472 178764
rect 295524 178712 295576 178764
rect 295708 178712 295760 178764
rect 296812 178712 296864 178764
rect 296996 178712 297048 178764
rect 250076 177284 250128 177336
rect 250352 177284 250404 177336
rect 310888 176740 310940 176792
rect 389548 176740 389600 176792
rect 463884 176672 463936 176724
rect 464068 176672 464120 176724
rect 310796 176604 310848 176656
rect 338856 176604 338908 176656
rect 374368 176604 374420 176656
rect 375840 176604 375892 176656
rect 389456 176604 389508 176656
rect 338856 176468 338908 176520
rect 374368 176468 374420 176520
rect 375840 176468 375892 176520
rect 366916 174063 366968 174072
rect 366916 174029 366925 174063
rect 366925 174029 366959 174063
rect 366959 174029 366968 174063
rect 366916 174020 366968 174029
rect 259736 173952 259788 174004
rect 366824 173952 366876 174004
rect 367008 173952 367060 174004
rect 230848 173884 230900 173936
rect 231032 173884 231084 173936
rect 235080 173884 235132 173936
rect 235172 173884 235224 173936
rect 236368 173884 236420 173936
rect 236460 173884 236512 173936
rect 239128 173884 239180 173936
rect 239220 173884 239272 173936
rect 251456 173884 251508 173936
rect 251640 173884 251692 173936
rect 266636 173884 266688 173936
rect 266820 173884 266872 173936
rect 323308 173884 323360 173936
rect 323492 173884 323544 173936
rect 327172 173884 327224 173936
rect 327264 173884 327316 173936
rect 331404 173884 331456 173936
rect 331588 173884 331640 173936
rect 337108 173884 337160 173936
rect 337384 173884 337436 173936
rect 339684 173884 339736 173936
rect 339868 173884 339920 173936
rect 357624 173884 357676 173936
rect 357900 173884 357952 173936
rect 360476 173884 360528 173936
rect 360568 173884 360620 173936
rect 366916 173927 366968 173936
rect 366916 173893 366925 173927
rect 366925 173893 366959 173927
rect 366959 173893 366968 173927
rect 366916 173884 366968 173893
rect 372528 173884 372580 173936
rect 372804 173884 372856 173936
rect 376944 173884 376996 173936
rect 377128 173884 377180 173936
rect 358820 173816 358872 173868
rect 232320 172567 232372 172576
rect 232320 172533 232329 172567
rect 232329 172533 232363 172567
rect 232363 172533 232372 172567
rect 232320 172524 232372 172533
rect 232228 172499 232280 172508
rect 232228 172465 232237 172499
rect 232237 172465 232271 172499
rect 232271 172465 232280 172499
rect 232228 172456 232280 172465
rect 270500 172456 270552 172508
rect 270776 172456 270828 172508
rect 301044 172456 301096 172508
rect 301136 172456 301188 172508
rect 330116 172456 330168 172508
rect 330300 172456 330352 172508
rect 337108 172499 337160 172508
rect 337108 172465 337117 172499
rect 337117 172465 337151 172499
rect 337151 172465 337160 172499
rect 337108 172456 337160 172465
rect 284944 171096 284996 171148
rect 267832 171071 267884 171080
rect 267832 171037 267841 171071
rect 267841 171037 267875 171071
rect 267875 171037 267884 171071
rect 267832 171028 267884 171037
rect 294420 171071 294472 171080
rect 294420 171037 294429 171071
rect 294429 171037 294463 171071
rect 294463 171037 294472 171071
rect 294420 171028 294472 171037
rect 306840 171028 306892 171080
rect 307024 171028 307076 171080
rect 341248 169779 341300 169788
rect 341248 169745 341257 169779
rect 341257 169745 341291 169779
rect 341291 169745 341300 169779
rect 341248 169736 341300 169745
rect 259736 169056 259788 169108
rect 259920 169056 259972 169108
rect 310796 167016 310848 167068
rect 310888 166880 310940 166932
rect 2780 165452 2832 165504
rect 5264 165452 5316 165504
rect 358728 164228 358780 164280
rect 358820 164228 358872 164280
rect 232228 164203 232280 164212
rect 232228 164169 232237 164203
rect 232237 164169 232271 164203
rect 232271 164169 232280 164203
rect 232228 164160 232280 164169
rect 244280 164160 244332 164212
rect 244464 164160 244516 164212
rect 251456 164160 251508 164212
rect 251640 164160 251692 164212
rect 259644 164160 259696 164212
rect 259828 164160 259880 164212
rect 295524 164160 295576 164212
rect 295708 164160 295760 164212
rect 337108 164203 337160 164212
rect 337108 164169 337117 164203
rect 337117 164169 337151 164203
rect 337151 164169 337160 164203
rect 337108 164160 337160 164169
rect 372804 164203 372856 164212
rect 372804 164169 372813 164203
rect 372813 164169 372847 164203
rect 372847 164169 372856 164203
rect 372804 164160 372856 164169
rect 376944 164160 376996 164212
rect 377128 164160 377180 164212
rect 463792 164160 463844 164212
rect 464068 164160 464120 164212
rect 284760 162868 284812 162920
rect 284944 162868 284996 162920
rect 285772 162800 285824 162852
rect 285956 162800 286008 162852
rect 325884 162800 325936 162852
rect 326160 162800 326212 162852
rect 329932 162800 329984 162852
rect 330116 162800 330168 162852
rect 357532 162800 357584 162852
rect 357808 162800 357860 162852
rect 358728 162843 358780 162852
rect 358728 162809 358737 162843
rect 358737 162809 358771 162843
rect 358771 162809 358780 162843
rect 358728 162800 358780 162809
rect 267832 162775 267884 162784
rect 267832 162741 267841 162775
rect 267841 162741 267875 162775
rect 267875 162741 267884 162775
rect 267832 162732 267884 162741
rect 262588 161440 262640 161492
rect 262680 161440 262732 161492
rect 265348 161440 265400 161492
rect 288900 161508 288952 161560
rect 290004 161508 290056 161560
rect 290096 161440 290148 161492
rect 294420 161483 294472 161492
rect 294420 161449 294429 161483
rect 294429 161449 294463 161483
rect 294463 161449 294472 161483
rect 294420 161440 294472 161449
rect 296996 161440 297048 161492
rect 297088 161440 297140 161492
rect 302516 161440 302568 161492
rect 302608 161440 302660 161492
rect 267832 161415 267884 161424
rect 267832 161381 267841 161415
rect 267841 161381 267875 161415
rect 267875 161381 267884 161415
rect 267832 161372 267884 161381
rect 288808 161372 288860 161424
rect 306840 161415 306892 161424
rect 306840 161381 306849 161415
rect 306849 161381 306883 161415
rect 306883 161381 306892 161415
rect 306840 161372 306892 161381
rect 291384 161304 291436 161356
rect 291568 161304 291620 161356
rect 288716 160012 288768 160064
rect 288808 160012 288860 160064
rect 291568 160012 291620 160064
rect 294420 160055 294472 160064
rect 294420 160021 294429 160055
rect 294429 160021 294463 160055
rect 294463 160021 294472 160055
rect 294420 160012 294472 160021
rect 341248 160055 341300 160064
rect 341248 160021 341257 160055
rect 341257 160021 341291 160055
rect 341291 160021 341300 160055
rect 341248 160012 341300 160021
rect 372804 159307 372856 159316
rect 372804 159273 372813 159307
rect 372813 159273 372847 159307
rect 372847 159273 372856 159307
rect 372804 159264 372856 159273
rect 417884 157496 417936 157548
rect 418160 157496 418212 157548
rect 437204 157496 437256 157548
rect 437480 157496 437532 157548
rect 456524 157496 456576 157548
rect 456892 157496 456944 157548
rect 306288 157428 306340 157480
rect 314568 157428 314620 157480
rect 230756 157360 230808 157412
rect 282644 157360 282696 157412
rect 288900 157360 288952 157412
rect 327172 157360 327224 157412
rect 230848 157292 230900 157344
rect 374368 157292 374420 157344
rect 375840 157292 375892 157344
rect 327264 157224 327316 157276
rect 374368 157156 374420 157208
rect 375840 157156 375892 157208
rect 339592 154640 339644 154692
rect 247224 154572 247276 154624
rect 247316 154572 247368 154624
rect 302516 154504 302568 154556
rect 302608 154504 302660 154556
rect 337200 154547 337252 154556
rect 337200 154513 337209 154547
rect 337209 154513 337243 154547
rect 337243 154513 337252 154547
rect 337200 154504 337252 154513
rect 339592 154504 339644 154556
rect 358728 154547 358780 154556
rect 358728 154513 358737 154547
rect 358737 154513 358771 154547
rect 358771 154513 358780 154547
rect 358728 154504 358780 154513
rect 367008 154547 367060 154556
rect 367008 154513 367017 154547
rect 367017 154513 367051 154547
rect 367051 154513 367060 154547
rect 367008 154504 367060 154513
rect 389456 154504 389508 154556
rect 389640 154504 389692 154556
rect 470416 154504 470468 154556
rect 470600 154504 470652 154556
rect 259828 154164 259880 154216
rect 272156 153212 272208 153264
rect 272248 153212 272300 153264
rect 285956 153144 286008 153196
rect 286048 153144 286100 153196
rect 302424 153144 302476 153196
rect 302516 153144 302568 153196
rect 310796 153187 310848 153196
rect 310796 153153 310805 153187
rect 310805 153153 310839 153187
rect 310839 153153 310848 153187
rect 310796 153144 310848 153153
rect 375840 153187 375892 153196
rect 375840 153153 375849 153187
rect 375849 153153 375883 153187
rect 375883 153153 375892 153187
rect 375840 153144 375892 153153
rect 264980 153076 265032 153128
rect 265348 153076 265400 153128
rect 337292 152328 337344 152380
rect 267832 151827 267884 151836
rect 267832 151793 267841 151827
rect 267841 151793 267875 151827
rect 267875 151793 267884 151827
rect 267832 151784 267884 151793
rect 296904 151784 296956 151836
rect 297088 151784 297140 151836
rect 306932 151784 306984 151836
rect 3332 151716 3384 151768
rect 17224 151716 17276 151768
rect 264980 151759 265032 151768
rect 264980 151725 264989 151759
rect 264989 151725 265023 151759
rect 265023 151725 265032 151759
rect 264980 151716 265032 151725
rect 339868 151716 339920 151768
rect 294512 150424 294564 150476
rect 294512 150288 294564 150340
rect 291476 149107 291528 149116
rect 291476 149073 291485 149107
rect 291485 149073 291519 149107
rect 291519 149073 291528 149107
rect 291476 149064 291528 149073
rect 338856 147636 338908 147688
rect 310796 147611 310848 147620
rect 310796 147577 310805 147611
rect 310805 147577 310839 147611
rect 310839 147577 310848 147611
rect 310796 147568 310848 147577
rect 338948 147568 339000 147620
rect 259644 145027 259696 145036
rect 259644 144993 259653 145027
rect 259653 144993 259687 145027
rect 259687 144993 259696 145027
rect 259644 144984 259696 144993
rect 357532 144916 357584 144968
rect 357808 144916 357860 144968
rect 358728 144916 358780 144968
rect 358820 144916 358872 144968
rect 367008 144959 367060 144968
rect 367008 144925 367017 144959
rect 367017 144925 367051 144959
rect 367051 144925 367060 144959
rect 367008 144916 367060 144925
rect 236000 144848 236052 144900
rect 236276 144848 236328 144900
rect 244280 144848 244332 144900
rect 244464 144848 244516 144900
rect 247132 144848 247184 144900
rect 247224 144848 247276 144900
rect 270684 144891 270736 144900
rect 270684 144857 270693 144891
rect 270693 144857 270727 144891
rect 270727 144857 270736 144891
rect 270684 144848 270736 144857
rect 272156 144848 272208 144900
rect 272248 144848 272300 144900
rect 323308 144848 323360 144900
rect 323400 144848 323452 144900
rect 324596 144848 324648 144900
rect 324780 144848 324832 144900
rect 325884 144848 325936 144900
rect 327172 144848 327224 144900
rect 327356 144848 327408 144900
rect 376944 144848 376996 144900
rect 377128 144848 377180 144900
rect 325976 144780 326028 144832
rect 265072 143556 265124 143608
rect 375840 143599 375892 143608
rect 375840 143565 375849 143599
rect 375849 143565 375883 143599
rect 375883 143565 375892 143599
rect 375840 143556 375892 143565
rect 250260 143531 250312 143540
rect 250260 143497 250269 143531
rect 250269 143497 250303 143531
rect 250303 143497 250312 143531
rect 250260 143488 250312 143497
rect 262588 143488 262640 143540
rect 262864 143488 262916 143540
rect 323308 143488 323360 143540
rect 323492 143488 323544 143540
rect 325976 143531 326028 143540
rect 325976 143497 325985 143531
rect 325985 143497 326019 143531
rect 326019 143497 326028 143531
rect 325976 143488 326028 143497
rect 330116 143531 330168 143540
rect 330116 143497 330125 143531
rect 330125 143497 330159 143531
rect 330159 143497 330168 143531
rect 330116 143488 330168 143497
rect 357256 143488 357308 143540
rect 357532 143488 357584 143540
rect 358728 143531 358780 143540
rect 358728 143497 358737 143531
rect 358737 143497 358771 143531
rect 358771 143497 358780 143531
rect 358728 143488 358780 143497
rect 360292 143531 360344 143540
rect 360292 143497 360301 143531
rect 360301 143497 360335 143531
rect 360335 143497 360344 143531
rect 360292 143488 360344 143497
rect 265072 143420 265124 143472
rect 341248 143395 341300 143404
rect 341248 143361 341257 143395
rect 341257 143361 341291 143395
rect 341291 143361 341300 143395
rect 341248 143352 341300 143361
rect 265256 142128 265308 142180
rect 288624 142128 288676 142180
rect 288808 142128 288860 142180
rect 290096 142128 290148 142180
rect 290188 142128 290240 142180
rect 317512 142128 317564 142180
rect 317696 142128 317748 142180
rect 339776 142171 339828 142180
rect 339776 142137 339785 142171
rect 339785 142137 339819 142171
rect 339819 142137 339828 142171
rect 339776 142128 339828 142137
rect 296812 142103 296864 142112
rect 296812 142069 296821 142103
rect 296821 142069 296855 142103
rect 296855 142069 296864 142103
rect 296812 142060 296864 142069
rect 301228 142060 301280 142112
rect 294236 140811 294288 140820
rect 294236 140777 294245 140811
rect 294245 140777 294279 140811
rect 294279 140777 294288 140811
rect 294236 140768 294288 140777
rect 270684 139995 270736 140004
rect 270684 139961 270693 139995
rect 270693 139961 270727 139995
rect 270727 139961 270736 139995
rect 270684 139952 270736 139961
rect 291476 139383 291528 139392
rect 291476 139349 291485 139383
rect 291485 139349 291519 139383
rect 291519 139349 291528 139383
rect 291476 139340 291528 139349
rect 310888 138660 310940 138712
rect 330208 138660 330260 138712
rect 372804 138116 372856 138168
rect 239128 137980 239180 138032
rect 338764 137980 338816 138032
rect 338948 137980 339000 138032
rect 389364 137980 389416 138032
rect 239220 137912 239272 137964
rect 317512 137912 317564 137964
rect 317788 137912 317840 137964
rect 360384 137912 360436 137964
rect 389456 137912 389508 137964
rect 299756 137368 299808 137420
rect 299940 137368 299992 137420
rect 306748 137368 306800 137420
rect 306932 137368 306984 137420
rect 2780 136348 2832 136400
rect 5172 136348 5224 136400
rect 372712 135303 372764 135312
rect 372712 135269 372721 135303
rect 372721 135269 372755 135303
rect 372755 135269 372764 135303
rect 372712 135260 372764 135269
rect 302516 135192 302568 135244
rect 302608 135192 302660 135244
rect 327264 135192 327316 135244
rect 358728 135235 358780 135244
rect 358728 135201 358737 135235
rect 358737 135201 358771 135235
rect 358771 135201 358780 135235
rect 358728 135192 358780 135201
rect 470416 135192 470468 135244
rect 470600 135192 470652 135244
rect 250352 133900 250404 133952
rect 302516 133875 302568 133884
rect 302516 133841 302525 133875
rect 302525 133841 302559 133875
rect 302559 133841 302568 133875
rect 302516 133832 302568 133841
rect 306748 133875 306800 133884
rect 306748 133841 306757 133875
rect 306757 133841 306791 133875
rect 306791 133841 306800 133875
rect 306748 133832 306800 133841
rect 337108 133875 337160 133884
rect 337108 133841 337117 133875
rect 337117 133841 337151 133875
rect 337151 133841 337160 133875
rect 337108 133832 337160 133841
rect 375840 133875 375892 133884
rect 375840 133841 375849 133875
rect 375849 133841 375883 133875
rect 375883 133841 375892 133875
rect 375840 133832 375892 133841
rect 389456 133875 389508 133884
rect 389456 133841 389465 133875
rect 389465 133841 389499 133875
rect 389499 133841 389508 133875
rect 389456 133832 389508 133841
rect 290004 132472 290056 132524
rect 290096 132472 290148 132524
rect 295524 132472 295576 132524
rect 295616 132472 295668 132524
rect 296904 132472 296956 132524
rect 301136 132515 301188 132524
rect 301136 132481 301145 132515
rect 301145 132481 301179 132515
rect 301179 132481 301188 132515
rect 301136 132472 301188 132481
rect 325976 132515 326028 132524
rect 325976 132481 325985 132515
rect 325985 132481 326019 132515
rect 326019 132481 326028 132515
rect 325976 132472 326028 132481
rect 284668 132447 284720 132456
rect 284668 132413 284677 132447
rect 284677 132413 284711 132447
rect 284711 132413 284720 132447
rect 284668 132404 284720 132413
rect 270500 130364 270552 130416
rect 270684 130364 270736 130416
rect 272156 130364 272208 130416
rect 272340 130364 272392 130416
rect 463884 130364 463936 130416
rect 464068 130364 464120 130416
rect 327172 129727 327224 129736
rect 327172 129693 327181 129727
rect 327181 129693 327215 129727
rect 327215 129693 327224 129727
rect 327172 129684 327224 129693
rect 259736 128324 259788 128376
rect 259828 128256 259880 128308
rect 310796 128299 310848 128308
rect 310796 128265 310805 128299
rect 310805 128265 310839 128299
rect 310839 128265 310848 128299
rect 310796 128256 310848 128265
rect 284668 126939 284720 126948
rect 284668 126905 284677 126939
rect 284677 126905 284711 126939
rect 284711 126905 284720 126939
rect 284668 126896 284720 126905
rect 358728 125604 358780 125656
rect 358820 125604 358872 125656
rect 251456 125579 251508 125588
rect 251456 125545 251465 125579
rect 251465 125545 251499 125579
rect 251499 125545 251508 125579
rect 251456 125536 251508 125545
rect 265164 125536 265216 125588
rect 265348 125536 265400 125588
rect 266544 125536 266596 125588
rect 266728 125536 266780 125588
rect 267740 125536 267792 125588
rect 267924 125536 267976 125588
rect 270684 125579 270736 125588
rect 270684 125545 270693 125579
rect 270693 125545 270727 125579
rect 270727 125545 270736 125579
rect 270684 125536 270736 125545
rect 272156 125579 272208 125588
rect 272156 125545 272165 125579
rect 272165 125545 272199 125579
rect 272199 125545 272208 125579
rect 272156 125536 272208 125545
rect 323216 125536 323268 125588
rect 323400 125536 323452 125588
rect 324596 125536 324648 125588
rect 324780 125536 324832 125588
rect 327172 125536 327224 125588
rect 327356 125536 327408 125588
rect 367008 125579 367060 125588
rect 367008 125545 367017 125579
rect 367017 125545 367051 125579
rect 367051 125545 367060 125579
rect 367008 125536 367060 125545
rect 372712 125579 372764 125588
rect 372712 125545 372721 125579
rect 372721 125545 372755 125579
rect 372755 125545 372764 125579
rect 372712 125536 372764 125545
rect 259736 125468 259788 125520
rect 259828 125468 259880 125520
rect 310888 125468 310940 125520
rect 302608 124176 302660 124228
rect 306840 124176 306892 124228
rect 330116 124176 330168 124228
rect 330300 124176 330352 124228
rect 337200 124176 337252 124228
rect 375840 124219 375892 124228
rect 375840 124185 375849 124219
rect 375849 124185 375883 124219
rect 375883 124185 375892 124219
rect 375840 124176 375892 124185
rect 300952 124108 301004 124160
rect 358728 124151 358780 124160
rect 358728 124117 358737 124151
rect 358737 124117 358771 124151
rect 358771 124117 358780 124151
rect 358728 124108 358780 124117
rect 300952 123972 301004 124024
rect 288808 122859 288860 122868
rect 288808 122825 288817 122859
rect 288817 122825 288851 122859
rect 288851 122825 288860 122859
rect 288808 122816 288860 122825
rect 389180 122816 389232 122868
rect 235172 122748 235224 122800
rect 239220 122748 239272 122800
rect 284668 122748 284720 122800
rect 284852 122748 284904 122800
rect 290004 122791 290056 122800
rect 290004 122757 290013 122791
rect 290013 122757 290047 122791
rect 290047 122757 290056 122791
rect 290004 122748 290056 122757
rect 301136 122791 301188 122800
rect 301136 122757 301145 122791
rect 301145 122757 301179 122791
rect 301179 122757 301188 122791
rect 301136 122748 301188 122757
rect 306840 122748 306892 122800
rect 330116 122791 330168 122800
rect 330116 122757 330125 122791
rect 330125 122757 330159 122791
rect 330159 122757 330168 122791
rect 330116 122748 330168 122757
rect 337200 122791 337252 122800
rect 337200 122757 337209 122791
rect 337209 122757 337243 122791
rect 337243 122757 337252 122791
rect 337200 122748 337252 122757
rect 296904 122723 296956 122732
rect 296904 122689 296913 122723
rect 296913 122689 296947 122723
rect 296947 122689 296956 122723
rect 296904 122680 296956 122689
rect 2780 122340 2832 122392
rect 5080 122340 5132 122392
rect 288808 121499 288860 121508
rect 288808 121465 288817 121499
rect 288817 121465 288851 121499
rect 288851 121465 288860 121499
rect 288808 121456 288860 121465
rect 291660 121456 291712 121508
rect 295800 121431 295852 121440
rect 295800 121397 295809 121431
rect 295809 121397 295843 121431
rect 295843 121397 295852 121431
rect 295800 121388 295852 121397
rect 244464 120708 244516 120760
rect 244648 120708 244700 120760
rect 267832 120640 267884 120692
rect 267924 120640 267976 120692
rect 270684 120683 270736 120692
rect 270684 120649 270693 120683
rect 270693 120649 270727 120683
rect 270727 120649 270736 120683
rect 270684 120640 270736 120649
rect 272156 120683 272208 120692
rect 272156 120649 272165 120683
rect 272165 120649 272199 120683
rect 272199 120649 272208 120683
rect 272156 120640 272208 120649
rect 273536 118736 273588 118788
rect 357532 118736 357584 118788
rect 360384 118668 360436 118720
rect 377128 118668 377180 118720
rect 463884 118668 463936 118720
rect 273536 118600 273588 118652
rect 357440 118600 357492 118652
rect 360476 118600 360528 118652
rect 463976 118600 464028 118652
rect 377128 118532 377180 118584
rect 239128 118031 239180 118040
rect 239128 117997 239137 118031
rect 239137 117997 239171 118031
rect 239171 117997 239180 118031
rect 239128 117988 239180 117997
rect 325976 117988 326028 118040
rect 337200 118031 337252 118040
rect 337200 117997 337209 118031
rect 337209 117997 337243 118031
rect 337243 117997 337252 118031
rect 337200 117988 337252 117997
rect 310796 116059 310848 116068
rect 310796 116025 310805 116059
rect 310805 116025 310839 116059
rect 310839 116025 310848 116059
rect 310796 116016 310848 116025
rect 367008 116059 367060 116068
rect 367008 116025 367017 116059
rect 367017 116025 367051 116059
rect 367051 116025 367060 116059
rect 367008 116016 367060 116025
rect 251456 115991 251508 116000
rect 251456 115957 251465 115991
rect 251465 115957 251499 115991
rect 251499 115957 251508 115991
rect 251456 115948 251508 115957
rect 372712 115991 372764 116000
rect 372712 115957 372721 115991
rect 372721 115957 372755 115991
rect 372755 115957 372764 115991
rect 372712 115948 372764 115957
rect 310796 115923 310848 115932
rect 310796 115889 310805 115923
rect 310805 115889 310839 115923
rect 310839 115889 310848 115923
rect 310796 115880 310848 115889
rect 367008 115923 367060 115932
rect 367008 115889 367017 115923
rect 367017 115889 367051 115923
rect 367051 115889 367060 115923
rect 367008 115880 367060 115889
rect 377128 115880 377180 115932
rect 358728 114563 358780 114572
rect 358728 114529 358737 114563
rect 358737 114529 358771 114563
rect 358771 114529 358780 114563
rect 358728 114520 358780 114529
rect 267832 114495 267884 114504
rect 267832 114461 267841 114495
rect 267841 114461 267875 114495
rect 267875 114461 267884 114495
rect 267832 114452 267884 114461
rect 374368 114495 374420 114504
rect 374368 114461 374377 114495
rect 374377 114461 374411 114495
rect 374411 114461 374420 114495
rect 374368 114452 374420 114461
rect 375840 114495 375892 114504
rect 375840 114461 375849 114495
rect 375849 114461 375883 114495
rect 375883 114461 375892 114495
rect 375840 114452 375892 114461
rect 301136 114427 301188 114436
rect 301136 114393 301145 114427
rect 301145 114393 301179 114427
rect 301179 114393 301188 114427
rect 301136 114384 301188 114393
rect 235080 113203 235132 113212
rect 235080 113169 235089 113203
rect 235089 113169 235123 113203
rect 235123 113169 235132 113203
rect 235080 113160 235132 113169
rect 290004 113203 290056 113212
rect 290004 113169 290013 113203
rect 290013 113169 290047 113203
rect 290047 113169 290056 113203
rect 290004 113160 290056 113169
rect 296904 113203 296956 113212
rect 296904 113169 296913 113203
rect 296913 113169 296947 113203
rect 296947 113169 296956 113203
rect 296904 113160 296956 113169
rect 302424 113160 302476 113212
rect 302608 113160 302660 113212
rect 306656 113203 306708 113212
rect 306656 113169 306665 113203
rect 306665 113169 306699 113203
rect 306699 113169 306708 113203
rect 306656 113160 306708 113169
rect 330116 113203 330168 113212
rect 330116 113169 330125 113203
rect 330125 113169 330159 113203
rect 330159 113169 330168 113203
rect 330116 113160 330168 113169
rect 327264 113092 327316 113144
rect 295524 111800 295576 111852
rect 456524 110644 456576 110696
rect 458824 110644 458876 110696
rect 307668 110576 307720 110628
rect 315948 110576 316000 110628
rect 417884 110576 417936 110628
rect 418160 110576 418212 110628
rect 437204 110576 437256 110628
rect 437480 110576 437532 110628
rect 270408 110440 270460 110492
rect 278688 110440 278740 110492
rect 272156 109012 272208 109064
rect 463792 109012 463844 109064
rect 463976 109012 464028 109064
rect 278780 108944 278832 108996
rect 279056 108944 279108 108996
rect 310796 108987 310848 108996
rect 310796 108953 310805 108987
rect 310805 108953 310839 108987
rect 310839 108953 310848 108987
rect 310796 108944 310848 108953
rect 272156 108876 272208 108928
rect 265164 106292 265216 106344
rect 265256 106292 265308 106344
rect 367008 106335 367060 106344
rect 367008 106301 367017 106335
rect 367017 106301 367051 106335
rect 367051 106301 367060 106335
rect 367008 106292 367060 106301
rect 377036 106335 377088 106344
rect 377036 106301 377045 106335
rect 377045 106301 377079 106335
rect 377079 106301 377088 106335
rect 377036 106292 377088 106301
rect 251456 106267 251508 106276
rect 251456 106233 251465 106267
rect 251465 106233 251499 106267
rect 251499 106233 251508 106267
rect 251456 106224 251508 106233
rect 259552 106224 259604 106276
rect 259828 106224 259880 106276
rect 266728 106224 266780 106276
rect 270684 106224 270736 106276
rect 272156 106224 272208 106276
rect 272248 106224 272300 106276
rect 317696 106224 317748 106276
rect 317880 106224 317932 106276
rect 357532 106224 357584 106276
rect 357624 106224 357676 106276
rect 377128 106267 377180 106276
rect 377128 106233 377137 106267
rect 377137 106233 377171 106267
rect 377171 106233 377180 106267
rect 377128 106224 377180 106233
rect 267832 106199 267884 106208
rect 267832 106165 267841 106199
rect 267841 106165 267875 106199
rect 267875 106165 267884 106199
rect 267832 106156 267884 106165
rect 270684 106088 270736 106140
rect 374368 104975 374420 104984
rect 374368 104941 374377 104975
rect 374377 104941 374411 104975
rect 374411 104941 374420 104975
rect 374368 104932 374420 104941
rect 375840 104975 375892 104984
rect 375840 104941 375849 104975
rect 375849 104941 375883 104975
rect 375883 104941 375892 104975
rect 375840 104932 375892 104941
rect 288716 104864 288768 104916
rect 288900 104864 288952 104916
rect 291568 104864 291620 104916
rect 291660 104864 291712 104916
rect 296812 104864 296864 104916
rect 296904 104864 296956 104916
rect 302424 104864 302476 104916
rect 302516 104864 302568 104916
rect 306656 104864 306708 104916
rect 306840 104864 306892 104916
rect 325884 104907 325936 104916
rect 325884 104873 325893 104907
rect 325893 104873 325927 104907
rect 325927 104873 325936 104907
rect 325884 104864 325936 104873
rect 230848 104839 230900 104848
rect 230848 104805 230857 104839
rect 230857 104805 230891 104839
rect 230891 104805 230900 104839
rect 230848 104796 230900 104805
rect 265164 104839 265216 104848
rect 265164 104805 265173 104839
rect 265173 104805 265207 104839
rect 265207 104805 265216 104839
rect 265164 104796 265216 104805
rect 267832 104839 267884 104848
rect 267832 104805 267841 104839
rect 267841 104805 267875 104839
rect 267875 104805 267884 104839
rect 267832 104796 267884 104805
rect 272248 104839 272300 104848
rect 272248 104805 272257 104839
rect 272257 104805 272291 104839
rect 272291 104805 272300 104839
rect 272248 104796 272300 104805
rect 273536 104839 273588 104848
rect 273536 104805 273545 104839
rect 273545 104805 273579 104839
rect 273579 104805 273588 104839
rect 273536 104796 273588 104805
rect 301136 104796 301188 104848
rect 301320 104796 301372 104848
rect 357624 104839 357676 104848
rect 357624 104805 357633 104839
rect 357633 104805 357667 104839
rect 357667 104805 357676 104839
rect 357624 104796 357676 104805
rect 358728 104839 358780 104848
rect 358728 104805 358737 104839
rect 358737 104805 358771 104839
rect 358771 104805 358780 104839
rect 358728 104796 358780 104805
rect 374368 104839 374420 104848
rect 374368 104805 374377 104839
rect 374377 104805 374411 104839
rect 374411 104805 374420 104839
rect 374368 104796 374420 104805
rect 375840 104839 375892 104848
rect 375840 104805 375849 104839
rect 375849 104805 375883 104839
rect 375883 104805 375892 104839
rect 375840 104796 375892 104805
rect 327172 103547 327224 103556
rect 327172 103513 327181 103547
rect 327181 103513 327215 103547
rect 327215 103513 327224 103547
rect 327172 103504 327224 103513
rect 285956 103479 286008 103488
rect 285956 103445 285965 103479
rect 285965 103445 285999 103479
rect 285999 103445 286008 103479
rect 285956 103436 286008 103445
rect 288716 103436 288768 103488
rect 337108 103436 337160 103488
rect 341156 103436 341208 103488
rect 288808 103368 288860 103420
rect 295524 101983 295576 101992
rect 295524 101949 295533 101983
rect 295533 101949 295567 101983
rect 295567 101949 295576 101983
rect 295524 101940 295576 101949
rect 235080 101396 235132 101448
rect 235264 101396 235316 101448
rect 232228 100036 232280 100088
rect 270684 100036 270736 100088
rect 270868 100036 270920 100088
rect 294236 100036 294288 100088
rect 294420 100036 294472 100088
rect 323400 99424 323452 99476
rect 239128 99356 239180 99408
rect 244372 99356 244424 99408
rect 278872 99356 278924 99408
rect 279056 99356 279108 99408
rect 244464 99288 244516 99340
rect 323400 99288 323452 99340
rect 374368 99331 374420 99340
rect 374368 99297 374377 99331
rect 374377 99297 374411 99331
rect 374411 99297 374420 99331
rect 374368 99288 374420 99297
rect 377128 99331 377180 99340
rect 377128 99297 377137 99331
rect 377137 99297 377171 99331
rect 377171 99297 377180 99331
rect 377128 99288 377180 99297
rect 239128 99220 239180 99272
rect 389456 99152 389508 99204
rect 306840 98676 306892 98728
rect 307024 98676 307076 98728
rect 330208 98719 330260 98728
rect 330208 98685 330217 98719
rect 330217 98685 330251 98719
rect 330251 98685 330260 98719
rect 330208 98676 330260 98685
rect 310888 96772 310940 96824
rect 250076 96636 250128 96688
rect 250168 96636 250220 96688
rect 251456 96679 251508 96688
rect 251456 96645 251465 96679
rect 251465 96645 251499 96679
rect 251499 96645 251508 96679
rect 251456 96636 251508 96645
rect 266636 96679 266688 96688
rect 266636 96645 266645 96679
rect 266645 96645 266679 96679
rect 266679 96645 266688 96679
rect 266636 96636 266688 96645
rect 302516 96636 302568 96688
rect 310796 96636 310848 96688
rect 236276 96611 236328 96620
rect 236276 96577 236285 96611
rect 236285 96577 236319 96611
rect 236319 96577 236328 96611
rect 236276 96568 236328 96577
rect 247132 96611 247184 96620
rect 247132 96577 247141 96611
rect 247141 96577 247175 96611
rect 247175 96577 247184 96611
rect 247132 96568 247184 96577
rect 265164 96611 265216 96620
rect 265164 96577 265173 96611
rect 265173 96577 265207 96611
rect 265207 96577 265216 96611
rect 265164 96568 265216 96577
rect 272340 96500 272392 96552
rect 317788 96611 317840 96620
rect 317788 96577 317797 96611
rect 317797 96577 317831 96611
rect 317831 96577 317840 96611
rect 317788 96568 317840 96577
rect 360292 96568 360344 96620
rect 360384 96568 360436 96620
rect 367008 96611 367060 96620
rect 367008 96577 367017 96611
rect 367017 96577 367051 96611
rect 367051 96577 367060 96611
rect 367008 96568 367060 96577
rect 302608 96500 302660 96552
rect 325976 95276 326028 95328
rect 230848 95251 230900 95260
rect 230848 95217 230857 95251
rect 230857 95217 230891 95251
rect 230891 95217 230900 95251
rect 230848 95208 230900 95217
rect 267924 95208 267976 95260
rect 273628 95208 273680 95260
rect 296812 95208 296864 95260
rect 326068 95208 326120 95260
rect 357624 95251 357676 95260
rect 357624 95217 357633 95251
rect 357633 95217 357667 95251
rect 357667 95217 357676 95251
rect 357624 95208 357676 95217
rect 358820 95208 358872 95260
rect 375840 95251 375892 95260
rect 375840 95217 375849 95251
rect 375849 95217 375883 95251
rect 375883 95217 375892 95251
rect 375840 95208 375892 95217
rect 290004 95140 290056 95192
rect 290096 95140 290148 95192
rect 324596 95140 324648 95192
rect 324780 95140 324832 95192
rect 339684 95140 339736 95192
rect 296996 95072 297048 95124
rect 291660 93916 291712 93968
rect 286140 93848 286192 93900
rect 291752 93848 291804 93900
rect 337200 93891 337252 93900
rect 337200 93857 337209 93891
rect 337209 93857 337243 93891
rect 337243 93857 337252 93891
rect 337200 93848 337252 93857
rect 463700 93848 463752 93900
rect 463884 93848 463936 93900
rect 301136 93823 301188 93832
rect 301136 93789 301145 93823
rect 301145 93789 301179 93823
rect 301179 93789 301188 93823
rect 301136 93780 301188 93789
rect 306748 93823 306800 93832
rect 306748 93789 306757 93823
rect 306757 93789 306791 93823
rect 306791 93789 306800 93823
rect 306748 93780 306800 93789
rect 295708 92488 295760 92540
rect 267924 92420 267976 92472
rect 268108 92420 268160 92472
rect 327264 90380 327316 90432
rect 327448 90380 327500 90432
rect 337016 90380 337068 90432
rect 337200 90380 337252 90432
rect 284760 90219 284812 90228
rect 284760 90185 284769 90219
rect 284769 90185 284803 90219
rect 284803 90185 284812 90219
rect 284760 90176 284812 90185
rect 247132 89675 247184 89684
rect 247132 89641 247141 89675
rect 247141 89641 247175 89675
rect 247175 89641 247184 89675
rect 247132 89632 247184 89641
rect 317788 89675 317840 89684
rect 317788 89641 317797 89675
rect 317797 89641 317831 89675
rect 317831 89641 317840 89675
rect 317788 89632 317840 89641
rect 389364 87907 389416 87916
rect 389364 87873 389373 87907
rect 389373 87873 389407 87907
rect 389407 87873 389416 87907
rect 389364 87864 389416 87873
rect 336924 87184 336976 87236
rect 395896 87184 395948 87236
rect 395988 87184 396040 87236
rect 251180 87048 251232 87100
rect 260656 87048 260708 87100
rect 376760 87048 376812 87100
rect 386236 87048 386288 87100
rect 386420 87048 386472 87100
rect 395804 87048 395856 87100
rect 437204 87116 437256 87168
rect 437480 87116 437532 87168
rect 456524 87116 456576 87168
rect 456984 87116 457036 87168
rect 494612 87116 494664 87168
rect 502248 87116 502300 87168
rect 417884 87048 417936 87100
rect 418160 87048 418212 87100
rect 232320 87023 232372 87032
rect 232320 86989 232329 87023
rect 232329 86989 232363 87023
rect 232363 86989 232372 87023
rect 232320 86980 232372 86989
rect 236276 87023 236328 87032
rect 236276 86989 236285 87023
rect 236285 86989 236319 87023
rect 236319 86989 236328 87023
rect 236276 86980 236328 86989
rect 295708 86980 295760 87032
rect 251456 86955 251508 86964
rect 251456 86921 251465 86955
rect 251465 86921 251499 86955
rect 251499 86921 251508 86955
rect 251456 86912 251508 86921
rect 326068 86980 326120 87032
rect 336924 86980 336976 87032
rect 367008 87023 367060 87032
rect 367008 86989 367017 87023
rect 367017 86989 367051 87023
rect 367051 86989 367060 87023
rect 367008 86980 367060 86989
rect 395896 86980 395948 87032
rect 395988 86980 396040 87032
rect 325976 86912 326028 86964
rect 330208 86955 330260 86964
rect 330208 86921 330217 86955
rect 330217 86921 330251 86955
rect 330251 86921 330260 86955
rect 330208 86912 330260 86921
rect 331312 86912 331364 86964
rect 331404 86912 331456 86964
rect 360384 86912 360436 86964
rect 295708 86844 295760 86896
rect 301228 86844 301280 86896
rect 317696 86844 317748 86896
rect 317880 86844 317932 86896
rect 331312 86776 331364 86828
rect 331404 86776 331456 86828
rect 286140 85620 286192 85672
rect 284760 85595 284812 85604
rect 284760 85561 284769 85595
rect 284769 85561 284803 85595
rect 284803 85561 284812 85595
rect 284760 85552 284812 85561
rect 286048 85552 286100 85604
rect 291660 85552 291712 85604
rect 294236 85552 294288 85604
rect 294420 85552 294472 85604
rect 358544 85552 358596 85604
rect 358636 85552 358688 85604
rect 232320 85527 232372 85536
rect 232320 85493 232329 85527
rect 232329 85493 232363 85527
rect 232363 85493 232372 85527
rect 232320 85484 232372 85493
rect 236276 85527 236328 85536
rect 236276 85493 236285 85527
rect 236285 85493 236319 85527
rect 236319 85493 236328 85527
rect 236276 85484 236328 85493
rect 324688 85484 324740 85536
rect 357532 85527 357584 85536
rect 357532 85493 357541 85527
rect 357541 85493 357575 85527
rect 357575 85493 357584 85527
rect 357532 85484 357584 85493
rect 291568 84235 291620 84244
rect 291568 84201 291577 84235
rect 291577 84201 291611 84235
rect 291611 84201 291620 84235
rect 291568 84192 291620 84201
rect 306840 84192 306892 84244
rect 270776 84167 270828 84176
rect 270776 84133 270785 84167
rect 270785 84133 270819 84167
rect 270819 84133 270828 84167
rect 270776 84124 270828 84133
rect 284760 84167 284812 84176
rect 284760 84133 284769 84167
rect 284769 84133 284803 84167
rect 284803 84133 284812 84167
rect 284760 84124 284812 84133
rect 337016 84124 337068 84176
rect 265256 82807 265308 82816
rect 265256 82773 265265 82807
rect 265265 82773 265299 82807
rect 265299 82773 265308 82807
rect 265256 82764 265308 82773
rect 267832 82764 267884 82816
rect 268016 82764 268068 82816
rect 301228 82807 301280 82816
rect 301228 82773 301237 82807
rect 301237 82773 301271 82807
rect 301271 82773 301280 82807
rect 301228 82764 301280 82773
rect 302608 82807 302660 82816
rect 302608 82773 302617 82807
rect 302617 82773 302651 82807
rect 302651 82773 302660 82807
rect 302608 82764 302660 82773
rect 249800 80724 249852 80776
rect 250076 80724 250128 80776
rect 247224 80223 247276 80232
rect 247224 80189 247233 80223
rect 247233 80189 247267 80223
rect 247267 80189 247276 80223
rect 247224 80180 247276 80189
rect 234988 80044 235040 80096
rect 235172 80044 235224 80096
rect 303896 80044 303948 80096
rect 338856 80044 338908 80096
rect 389364 80044 389416 80096
rect 463792 80044 463844 80096
rect 303896 79908 303948 79960
rect 338856 79908 338908 79960
rect 372436 79908 372488 79960
rect 372804 79908 372856 79960
rect 389456 79908 389508 79960
rect 463792 79908 463844 79960
rect 2780 79840 2832 79892
rect 4988 79840 5040 79892
rect 286048 78480 286100 78532
rect 367008 77392 367060 77444
rect 336832 77324 336884 77376
rect 336924 77324 336976 77376
rect 247224 77299 247276 77308
rect 247224 77265 247233 77299
rect 247233 77265 247267 77299
rect 247267 77265 247276 77299
rect 247224 77256 247276 77265
rect 251456 77299 251508 77308
rect 251456 77265 251465 77299
rect 251465 77265 251499 77299
rect 251499 77265 251508 77299
rect 251456 77256 251508 77265
rect 266636 77256 266688 77308
rect 266728 77256 266780 77308
rect 299756 77256 299808 77308
rect 299848 77256 299900 77308
rect 323400 77299 323452 77308
rect 323400 77265 323409 77299
rect 323409 77265 323443 77299
rect 323443 77265 323452 77299
rect 323400 77256 323452 77265
rect 339776 77299 339828 77308
rect 339776 77265 339785 77299
rect 339785 77265 339819 77299
rect 339819 77265 339828 77299
rect 339776 77256 339828 77265
rect 341064 77299 341116 77308
rect 341064 77265 341073 77299
rect 341073 77265 341107 77299
rect 341107 77265 341116 77299
rect 341064 77256 341116 77265
rect 360200 77299 360252 77308
rect 360200 77265 360209 77299
rect 360209 77265 360243 77299
rect 360243 77265 360252 77299
rect 360200 77256 360252 77265
rect 367008 77256 367060 77308
rect 272248 77188 272300 77240
rect 272340 77188 272392 77240
rect 303896 77188 303948 77240
rect 303988 77188 304040 77240
rect 336832 77188 336884 77240
rect 336924 77188 336976 77240
rect 389456 77188 389508 77240
rect 341064 77163 341116 77172
rect 341064 77129 341073 77163
rect 341073 77129 341107 77163
rect 341107 77129 341116 77163
rect 341064 77120 341116 77129
rect 309048 76236 309100 76288
rect 317328 76236 317380 76288
rect 417884 76100 417936 76152
rect 420368 76100 420420 76152
rect 253848 76032 253900 76084
rect 259276 76032 259328 76084
rect 437204 76032 437256 76084
rect 437480 76032 437532 76084
rect 456524 76032 456576 76084
rect 456800 76032 456852 76084
rect 232320 75939 232372 75948
rect 232320 75905 232329 75939
rect 232329 75905 232363 75939
rect 232363 75905 232372 75939
rect 232320 75896 232372 75905
rect 236276 75939 236328 75948
rect 236276 75905 236285 75939
rect 236285 75905 236319 75939
rect 236319 75905 236328 75939
rect 236276 75896 236328 75905
rect 288716 75896 288768 75948
rect 288808 75896 288860 75948
rect 289912 75896 289964 75948
rect 290096 75896 290148 75948
rect 291384 75896 291436 75948
rect 291568 75896 291620 75948
rect 295524 75896 295576 75948
rect 295708 75896 295760 75948
rect 296812 75896 296864 75948
rect 296996 75896 297048 75948
rect 323400 75939 323452 75948
rect 323400 75905 323409 75939
rect 323409 75905 323443 75939
rect 323443 75905 323452 75939
rect 323400 75896 323452 75905
rect 324596 75939 324648 75948
rect 324596 75905 324605 75939
rect 324605 75905 324639 75939
rect 324639 75905 324648 75939
rect 324596 75896 324648 75905
rect 357624 75896 357676 75948
rect 358544 75896 358596 75948
rect 358728 75896 358780 75948
rect 250076 75871 250128 75880
rect 250076 75837 250085 75871
rect 250085 75837 250119 75871
rect 250119 75837 250128 75871
rect 250076 75828 250128 75837
rect 272248 75828 272300 75880
rect 372804 75828 372856 75880
rect 284852 75760 284904 75812
rect 270776 74579 270828 74588
rect 270776 74545 270785 74579
rect 270785 74545 270819 74579
rect 270819 74545 270828 74579
rect 270776 74536 270828 74545
rect 306748 74536 306800 74588
rect 306840 74536 306892 74588
rect 266728 74511 266780 74520
rect 266728 74477 266737 74511
rect 266737 74477 266771 74511
rect 266771 74477 266780 74511
rect 266728 74468 266780 74477
rect 288716 74468 288768 74520
rect 288992 74468 289044 74520
rect 265256 73219 265308 73228
rect 265256 73185 265265 73219
rect 265265 73185 265299 73219
rect 265299 73185 265308 73219
rect 265256 73176 265308 73185
rect 301228 73219 301280 73228
rect 301228 73185 301237 73219
rect 301237 73185 301271 73219
rect 301271 73185 301280 73219
rect 301228 73176 301280 73185
rect 302700 73176 302752 73228
rect 324596 72428 324648 72480
rect 324780 72428 324832 72480
rect 267832 71748 267884 71800
rect 268016 71748 268068 71800
rect 239128 70456 239180 70508
rect 244464 70499 244516 70508
rect 244464 70465 244473 70499
rect 244473 70465 244507 70499
rect 244507 70465 244516 70499
rect 244464 70456 244516 70465
rect 273628 70456 273680 70508
rect 325976 70456 326028 70508
rect 239128 70320 239180 70372
rect 325884 70320 325936 70372
rect 341156 70252 341208 70304
rect 301228 69640 301280 69692
rect 236276 67600 236328 67652
rect 273536 67643 273588 67652
rect 273536 67609 273545 67643
rect 273545 67609 273579 67643
rect 273579 67609 273588 67643
rect 273536 67600 273588 67609
rect 323308 67600 323360 67652
rect 323400 67600 323452 67652
rect 330116 67600 330168 67652
rect 330300 67600 330352 67652
rect 389364 67643 389416 67652
rect 389364 67609 389373 67643
rect 389373 67609 389407 67643
rect 389407 67609 389416 67643
rect 389364 67600 389416 67609
rect 236368 67532 236420 67584
rect 247132 67532 247184 67584
rect 247224 67532 247276 67584
rect 244464 66283 244516 66292
rect 244464 66249 244473 66283
rect 244473 66249 244507 66283
rect 244507 66249 244516 66283
rect 244464 66240 244516 66249
rect 250076 66283 250128 66292
rect 250076 66249 250085 66283
rect 250085 66249 250119 66283
rect 250119 66249 250128 66283
rect 250076 66240 250128 66249
rect 259644 66240 259696 66292
rect 259736 66240 259788 66292
rect 272156 66283 272208 66292
rect 272156 66249 272165 66283
rect 272165 66249 272199 66283
rect 272199 66249 272208 66283
rect 272156 66240 272208 66249
rect 285956 66283 286008 66292
rect 285956 66249 285965 66283
rect 285965 66249 285999 66283
rect 285999 66249 286008 66283
rect 285956 66240 286008 66249
rect 337200 66283 337252 66292
rect 337200 66249 337209 66283
rect 337209 66249 337243 66283
rect 337243 66249 337252 66283
rect 337200 66240 337252 66249
rect 372712 66283 372764 66292
rect 372712 66249 372721 66283
rect 372721 66249 372755 66283
rect 372755 66249 372764 66283
rect 372712 66240 372764 66249
rect 232320 66215 232372 66224
rect 232320 66181 232329 66215
rect 232329 66181 232363 66215
rect 232363 66181 232372 66215
rect 232320 66172 232372 66181
rect 270684 66215 270736 66224
rect 270684 66181 270693 66215
rect 270693 66181 270727 66215
rect 270727 66181 270736 66215
rect 270684 66172 270736 66181
rect 296812 66215 296864 66224
rect 296812 66181 296821 66215
rect 296821 66181 296855 66215
rect 296855 66181 296864 66215
rect 296812 66172 296864 66181
rect 310796 66215 310848 66224
rect 310796 66181 310805 66215
rect 310805 66181 310839 66215
rect 310839 66181 310848 66215
rect 310796 66172 310848 66181
rect 323308 66215 323360 66224
rect 323308 66181 323317 66215
rect 323317 66181 323351 66215
rect 323351 66181 323360 66215
rect 323308 66172 323360 66181
rect 324780 66172 324832 66224
rect 330116 66172 330168 66224
rect 266912 64880 266964 64932
rect 3332 64812 3384 64864
rect 24124 64812 24176 64864
rect 294236 64855 294288 64864
rect 294236 64821 294245 64855
rect 294245 64821 294279 64855
rect 294279 64821 294288 64855
rect 294236 64812 294288 64821
rect 273168 63656 273220 63708
rect 278688 63656 278740 63708
rect 417884 63656 417936 63708
rect 418160 63656 418212 63708
rect 437204 63656 437256 63708
rect 437480 63656 437532 63708
rect 456524 63656 456576 63708
rect 456892 63656 456944 63708
rect 265348 63452 265400 63504
rect 230848 61412 230900 61464
rect 236368 61412 236420 61464
rect 272156 60732 272208 60784
rect 273444 60664 273496 60716
rect 273628 60664 273680 60716
rect 310796 60707 310848 60716
rect 310796 60673 310805 60707
rect 310805 60673 310839 60707
rect 310839 60673 310848 60707
rect 310796 60664 310848 60673
rect 341156 60664 341208 60716
rect 341340 60664 341392 60716
rect 360292 60664 360344 60716
rect 360476 60664 360528 60716
rect 272156 60596 272208 60648
rect 262680 60367 262732 60376
rect 262680 60333 262689 60367
rect 262689 60333 262723 60367
rect 262723 60333 262732 60367
rect 262680 60324 262732 60333
rect 302700 59508 302752 59560
rect 325884 58012 325936 58064
rect 284760 57944 284812 57996
rect 284852 57944 284904 57996
rect 285956 57944 286008 57996
rect 286048 57944 286100 57996
rect 327172 57944 327224 57996
rect 325884 57876 325936 57928
rect 341340 57919 341392 57928
rect 341340 57885 341349 57919
rect 341349 57885 341383 57919
rect 341383 57885 341392 57919
rect 341340 57876 341392 57885
rect 360384 57876 360436 57928
rect 360476 57876 360528 57928
rect 367008 57919 367060 57928
rect 367008 57885 367017 57919
rect 367017 57885 367051 57919
rect 367051 57885 367060 57919
rect 367008 57876 367060 57885
rect 389180 57919 389232 57928
rect 389180 57885 389189 57919
rect 389189 57885 389223 57919
rect 389223 57885 389232 57919
rect 389180 57876 389232 57885
rect 470600 57919 470652 57928
rect 470600 57885 470609 57919
rect 470609 57885 470643 57919
rect 470643 57885 470652 57919
rect 470600 57876 470652 57885
rect 327264 57808 327316 57860
rect 295524 57035 295576 57044
rect 295524 57001 295533 57035
rect 295533 57001 295567 57035
rect 295567 57001 295576 57035
rect 295524 56992 295576 57001
rect 232320 56627 232372 56636
rect 232320 56593 232329 56627
rect 232329 56593 232363 56627
rect 232363 56593 232372 56627
rect 232320 56584 232372 56593
rect 259644 56584 259696 56636
rect 324688 56627 324740 56636
rect 324688 56593 324697 56627
rect 324697 56593 324731 56627
rect 324731 56593 324740 56627
rect 324688 56584 324740 56593
rect 329932 56627 329984 56636
rect 329932 56593 329941 56627
rect 329941 56593 329975 56627
rect 329975 56593 329984 56627
rect 329932 56584 329984 56593
rect 358728 56584 358780 56636
rect 358820 56584 358872 56636
rect 250076 56559 250128 56568
rect 250076 56525 250085 56559
rect 250085 56525 250119 56559
rect 250119 56525 250128 56559
rect 250076 56516 250128 56525
rect 259552 56516 259604 56568
rect 286048 56516 286100 56568
rect 310796 56516 310848 56568
rect 310888 56516 310940 56568
rect 339684 56559 339736 56568
rect 339684 56525 339693 56559
rect 339693 56525 339727 56559
rect 339727 56525 339736 56559
rect 339684 56516 339736 56525
rect 296812 56219 296864 56228
rect 296812 56185 296821 56219
rect 296821 56185 296855 56219
rect 296855 56185 296864 56219
rect 296812 56176 296864 56185
rect 262772 55224 262824 55276
rect 294236 55267 294288 55276
rect 294236 55233 294245 55267
rect 294245 55233 294279 55267
rect 294279 55233 294288 55267
rect 294236 55224 294288 55233
rect 317512 55224 317564 55276
rect 317696 55224 317748 55276
rect 301228 55088 301280 55140
rect 244372 53796 244424 53848
rect 244464 53796 244516 53848
rect 265256 53839 265308 53848
rect 265256 53805 265265 53839
rect 265265 53805 265299 53839
rect 265299 53805 265308 53839
rect 265256 53796 265308 53805
rect 232320 53048 232372 53100
rect 267832 52436 267884 52488
rect 268016 52436 268068 52488
rect 273628 51076 273680 51128
rect 250076 51051 250128 51060
rect 250076 51017 250085 51051
rect 250085 51017 250119 51051
rect 250119 51017 250128 51051
rect 250076 51008 250128 51017
rect 273536 51008 273588 51060
rect 341432 50872 341484 50924
rect 2780 50124 2832 50176
rect 4896 50124 4948 50176
rect 236276 48399 236328 48408
rect 236276 48365 236285 48399
rect 236285 48365 236319 48399
rect 236319 48365 236328 48399
rect 236276 48356 236328 48365
rect 303896 48356 303948 48408
rect 230756 48331 230808 48340
rect 230756 48297 230765 48331
rect 230765 48297 230799 48331
rect 230799 48297 230808 48331
rect 230756 48288 230808 48297
rect 288716 48288 288768 48340
rect 288992 48288 289044 48340
rect 295524 48331 295576 48340
rect 295524 48297 295533 48331
rect 295533 48297 295567 48331
rect 295567 48297 295576 48331
rect 295524 48288 295576 48297
rect 323308 48331 323360 48340
rect 323308 48297 323317 48331
rect 323317 48297 323351 48331
rect 323351 48297 323360 48331
rect 323308 48288 323360 48297
rect 324688 48288 324740 48340
rect 324780 48288 324832 48340
rect 358728 48331 358780 48340
rect 358728 48297 358737 48331
rect 358737 48297 358771 48331
rect 358771 48297 358780 48331
rect 358728 48288 358780 48297
rect 367008 48331 367060 48340
rect 367008 48297 367017 48331
rect 367017 48297 367051 48331
rect 367051 48297 367060 48331
rect 367008 48288 367060 48297
rect 389272 48288 389324 48340
rect 470600 48331 470652 48340
rect 470600 48297 470609 48331
rect 470609 48297 470643 48331
rect 470643 48297 470652 48331
rect 470600 48288 470652 48297
rect 273536 48263 273588 48272
rect 273536 48229 273545 48263
rect 273545 48229 273579 48263
rect 273579 48229 273588 48263
rect 273536 48220 273588 48229
rect 303896 48220 303948 48272
rect 325884 48220 325936 48272
rect 327172 48220 327224 48272
rect 327356 48220 327408 48272
rect 325976 48152 326028 48204
rect 262772 46996 262824 47048
rect 268016 46928 268068 46980
rect 285956 46971 286008 46980
rect 285956 46937 285965 46971
rect 285965 46937 285999 46971
rect 285999 46937 286008 46971
rect 285956 46928 286008 46937
rect 302516 46971 302568 46980
rect 302516 46937 302525 46971
rect 302525 46937 302559 46971
rect 302559 46937 302568 46971
rect 302516 46928 302568 46937
rect 339960 46928 340012 46980
rect 358728 46971 358780 46980
rect 358728 46937 358737 46971
rect 358737 46937 358771 46971
rect 358771 46937 358780 46971
rect 358728 46928 358780 46937
rect 236276 46903 236328 46912
rect 236276 46869 236285 46903
rect 236285 46869 236319 46903
rect 236319 46869 236328 46903
rect 236276 46860 236328 46869
rect 247132 46903 247184 46912
rect 247132 46869 247141 46903
rect 247141 46869 247175 46903
rect 247175 46869 247184 46903
rect 247132 46860 247184 46869
rect 250168 46860 250220 46912
rect 251364 46903 251416 46912
rect 251364 46869 251373 46903
rect 251373 46869 251407 46903
rect 251407 46869 251416 46903
rect 251364 46860 251416 46869
rect 262680 46860 262732 46912
rect 267740 46860 267792 46912
rect 306748 46860 306800 46912
rect 323308 46903 323360 46912
rect 323308 46869 323317 46903
rect 323317 46869 323351 46903
rect 323351 46869 323360 46903
rect 323308 46860 323360 46869
rect 324780 46860 324832 46912
rect 325976 46860 326028 46912
rect 326068 46860 326120 46912
rect 327356 46903 327408 46912
rect 327356 46869 327365 46903
rect 327365 46869 327399 46903
rect 327399 46869 327408 46903
rect 327356 46860 327408 46869
rect 330116 46903 330168 46912
rect 330116 46869 330125 46903
rect 330125 46869 330159 46903
rect 330159 46869 330168 46903
rect 330116 46860 330168 46869
rect 338488 46860 338540 46912
rect 338948 46860 339000 46912
rect 296812 46835 296864 46844
rect 296812 46801 296821 46835
rect 296821 46801 296855 46835
rect 296855 46801 296864 46835
rect 296812 46792 296864 46801
rect 306840 46792 306892 46844
rect 294236 45500 294288 45552
rect 294420 45500 294472 45552
rect 310888 45500 310940 45552
rect 311072 45500 311124 45552
rect 317512 45500 317564 45552
rect 317696 45500 317748 45552
rect 338488 45543 338540 45552
rect 338488 45509 338497 45543
rect 338497 45509 338531 45543
rect 338531 45509 338540 45543
rect 338488 45500 338540 45509
rect 284668 44684 284720 44736
rect 266636 44140 266688 44192
rect 266912 44140 266964 44192
rect 272156 44140 272208 44192
rect 272432 44140 272484 44192
rect 296904 43936 296956 43988
rect 270684 42848 270736 42900
rect 303896 42032 303948 42084
rect 265256 41463 265308 41472
rect 265256 41429 265265 41463
rect 265265 41429 265299 41463
rect 265299 41429 265308 41463
rect 265256 41420 265308 41429
rect 341432 41463 341484 41472
rect 341432 41429 341441 41463
rect 341441 41429 341475 41463
rect 341475 41429 341484 41463
rect 341432 41420 341484 41429
rect 266636 41395 266688 41404
rect 266636 41361 266645 41395
rect 266645 41361 266679 41395
rect 266679 41361 266688 41395
rect 266636 41352 266688 41361
rect 360292 41352 360344 41404
rect 360476 41352 360528 41404
rect 377128 41327 377180 41336
rect 377128 41293 377137 41327
rect 377137 41293 377171 41327
rect 377171 41293 377180 41327
rect 377128 41284 377180 41293
rect 241428 40264 241480 40316
rect 245016 40264 245068 40316
rect 417884 40196 417936 40248
rect 420368 40196 420420 40248
rect 437204 40196 437256 40248
rect 437480 40196 437532 40248
rect 456524 40128 456576 40180
rect 456892 40128 456944 40180
rect 253848 40060 253900 40112
rect 262864 40060 262916 40112
rect 230756 38743 230808 38752
rect 230756 38709 230765 38743
rect 230765 38709 230799 38743
rect 230799 38709 230808 38743
rect 230756 38700 230808 38709
rect 232228 38743 232280 38752
rect 232228 38709 232237 38743
rect 232237 38709 232271 38743
rect 232271 38709 232280 38743
rect 232228 38700 232280 38709
rect 377036 38700 377088 38752
rect 273536 38675 273588 38684
rect 273536 38641 273545 38675
rect 273545 38641 273579 38675
rect 273579 38641 273588 38675
rect 273536 38632 273588 38641
rect 295524 38632 295576 38684
rect 341432 38607 341484 38616
rect 341432 38573 341441 38607
rect 341441 38573 341475 38607
rect 341475 38573 341484 38607
rect 341432 38564 341484 38573
rect 367008 38607 367060 38616
rect 367008 38573 367017 38607
rect 367017 38573 367051 38607
rect 367051 38573 367060 38607
rect 367008 38564 367060 38573
rect 377128 38564 377180 38616
rect 377312 38564 377364 38616
rect 295616 38496 295668 38548
rect 327356 38539 327408 38548
rect 327356 38505 327365 38539
rect 327365 38505 327399 38539
rect 327399 38505 327408 38539
rect 327356 38496 327408 38505
rect 286048 37340 286100 37392
rect 300032 37340 300084 37392
rect 230756 37315 230808 37324
rect 230756 37281 230765 37315
rect 230765 37281 230799 37315
rect 230799 37281 230808 37315
rect 230756 37272 230808 37281
rect 236460 37272 236512 37324
rect 250076 37315 250128 37324
rect 250076 37281 250085 37315
rect 250085 37281 250119 37315
rect 250119 37281 250128 37315
rect 250076 37272 250128 37281
rect 251456 37272 251508 37324
rect 285956 37272 286008 37324
rect 323308 37315 323360 37324
rect 323308 37281 323317 37315
rect 323317 37281 323351 37315
rect 323351 37281 323360 37315
rect 323308 37272 323360 37281
rect 324688 37315 324740 37324
rect 324688 37281 324697 37315
rect 324697 37281 324731 37315
rect 324731 37281 324740 37315
rect 324688 37272 324740 37281
rect 330116 37315 330168 37324
rect 330116 37281 330125 37315
rect 330125 37281 330159 37315
rect 330159 37281 330168 37315
rect 330116 37272 330168 37281
rect 339776 37272 339828 37324
rect 339960 37272 340012 37324
rect 358728 37272 358780 37324
rect 358820 37272 358872 37324
rect 288716 37247 288768 37256
rect 288716 37213 288725 37247
rect 288725 37213 288759 37247
rect 288759 37213 288768 37247
rect 288716 37204 288768 37213
rect 265256 35955 265308 35964
rect 265256 35921 265265 35955
rect 265265 35921 265299 35955
rect 265299 35921 265308 35955
rect 265256 35912 265308 35921
rect 3148 35844 3200 35896
rect 6184 35844 6236 35896
rect 251456 35887 251508 35896
rect 251456 35853 251465 35887
rect 251465 35853 251499 35887
rect 251499 35853 251508 35887
rect 251456 35844 251508 35853
rect 244372 34484 244424 34536
rect 244556 34484 244608 34536
rect 247132 34527 247184 34536
rect 247132 34493 247141 34527
rect 247141 34493 247175 34527
rect 247175 34493 247184 34527
rect 247132 34484 247184 34493
rect 272248 34484 272300 34536
rect 272432 34484 272484 34536
rect 266636 34459 266688 34468
rect 266636 34425 266645 34459
rect 266645 34425 266679 34459
rect 266679 34425 266688 34459
rect 266636 34416 266688 34425
rect 303896 32376 303948 32428
rect 372712 31875 372764 31884
rect 372712 31841 372721 31875
rect 372721 31841 372755 31875
rect 372755 31841 372764 31875
rect 372712 31832 372764 31841
rect 239128 31764 239180 31816
rect 317512 31764 317564 31816
rect 317696 31764 317748 31816
rect 360476 31764 360528 31816
rect 389364 31764 389416 31816
rect 239036 31696 239088 31748
rect 360292 31696 360344 31748
rect 389456 31628 389508 31680
rect 248420 29180 248472 29232
rect 257896 29180 257948 29232
rect 417884 29180 417936 29232
rect 418804 29180 418856 29232
rect 456524 29180 456576 29232
rect 456984 29180 457036 29232
rect 437204 29112 437256 29164
rect 437480 29112 437532 29164
rect 284760 29019 284812 29028
rect 284760 28985 284769 29019
rect 284769 28985 284803 29019
rect 284803 28985 284812 29019
rect 284760 28976 284812 28985
rect 285956 28976 286008 29028
rect 286048 28976 286100 29028
rect 295524 28976 295576 29028
rect 295616 28976 295668 29028
rect 301320 29044 301372 29096
rect 367008 29087 367060 29096
rect 367008 29053 367017 29087
rect 367017 29053 367051 29087
rect 367051 29053 367060 29087
rect 367008 29044 367060 29053
rect 367100 29044 367152 29096
rect 376668 29044 376720 29096
rect 492772 29044 492824 29096
rect 502248 29044 502300 29096
rect 327172 28976 327224 29028
rect 327356 28976 327408 29028
rect 341156 28976 341208 29028
rect 341432 28976 341484 29028
rect 372712 29019 372764 29028
rect 372712 28985 372721 29019
rect 372721 28985 372755 29019
rect 372755 28985 372764 29019
rect 372712 28976 372764 28985
rect 232228 28908 232280 28960
rect 232320 28908 232372 28960
rect 236368 28951 236420 28960
rect 236368 28917 236377 28951
rect 236377 28917 236411 28951
rect 236411 28917 236420 28951
rect 236368 28908 236420 28917
rect 301228 28908 301280 28960
rect 323216 28908 323268 28960
rect 323400 28908 323452 28960
rect 357624 28908 357676 28960
rect 357808 28908 357860 28960
rect 367008 28951 367060 28960
rect 367008 28917 367017 28951
rect 367017 28917 367051 28951
rect 367051 28917 367060 28951
rect 367008 28908 367060 28917
rect 375840 28951 375892 28960
rect 375840 28917 375849 28951
rect 375849 28917 375883 28951
rect 375883 28917 375892 28951
rect 375840 28908 375892 28917
rect 377128 28951 377180 28960
rect 377128 28917 377137 28951
rect 377137 28917 377171 28951
rect 377171 28917 377180 28951
rect 377128 28908 377180 28917
rect 307668 28840 307720 28892
rect 315948 28840 316000 28892
rect 259736 27616 259788 27668
rect 259828 27616 259880 27668
rect 288808 27616 288860 27668
rect 338672 27616 338724 27668
rect 265256 27548 265308 27600
rect 286048 27548 286100 27600
rect 295524 27591 295576 27600
rect 295524 27557 295533 27591
rect 295533 27557 295567 27591
rect 295567 27557 295576 27591
rect 295524 27548 295576 27557
rect 330208 27548 330260 27600
rect 358636 27548 358688 27600
rect 301228 27480 301280 27532
rect 247040 26324 247092 26376
rect 247132 26324 247184 26376
rect 251456 26299 251508 26308
rect 251456 26265 251465 26299
rect 251465 26265 251499 26299
rect 251499 26265 251508 26299
rect 251456 26256 251508 26265
rect 249984 26188 250036 26240
rect 250168 26188 250220 26240
rect 288808 26231 288860 26240
rect 288808 26197 288817 26231
rect 288817 26197 288851 26231
rect 288851 26197 288860 26231
rect 288808 26188 288860 26197
rect 310888 26231 310940 26240
rect 310888 26197 310897 26231
rect 310897 26197 310931 26231
rect 310931 26197 310940 26231
rect 310888 26188 310940 26197
rect 266728 24896 266780 24948
rect 244464 24760 244516 24812
rect 266636 24760 266688 24812
rect 337200 24284 337252 24336
rect 270500 22176 270552 22228
rect 270776 22176 270828 22228
rect 247224 22108 247276 22160
rect 268016 22108 268068 22160
rect 272248 22108 272300 22160
rect 374368 22108 374420 22160
rect 247132 22040 247184 22092
rect 372712 22040 372764 22092
rect 377128 22083 377180 22092
rect 377128 22049 377137 22083
rect 377137 22049 377171 22083
rect 377171 22049 377180 22083
rect 377128 22040 377180 22049
rect 372804 21972 372856 22024
rect 374368 21972 374420 22024
rect 239036 19388 239088 19440
rect 236368 19363 236420 19372
rect 236368 19329 236377 19363
rect 236377 19329 236411 19363
rect 236411 19329 236420 19363
rect 236368 19320 236420 19329
rect 302516 19320 302568 19372
rect 302608 19320 302660 19372
rect 306748 19320 306800 19372
rect 306840 19320 306892 19372
rect 337108 19363 337160 19372
rect 337108 19329 337117 19363
rect 337117 19329 337151 19363
rect 337151 19329 337160 19363
rect 337108 19320 337160 19329
rect 338672 19320 338724 19372
rect 338856 19320 338908 19372
rect 367008 19363 367060 19372
rect 367008 19329 367017 19363
rect 367017 19329 367051 19363
rect 367051 19329 367060 19363
rect 367008 19320 367060 19329
rect 375840 19363 375892 19372
rect 375840 19329 375849 19363
rect 375849 19329 375883 19363
rect 375883 19329 375892 19363
rect 375840 19320 375892 19329
rect 239036 19252 239088 19304
rect 366916 19295 366968 19304
rect 366916 19261 366925 19295
rect 366925 19261 366959 19295
rect 366959 19261 366968 19295
rect 366916 19252 366968 19261
rect 366824 19184 366876 19236
rect 367008 19184 367060 19236
rect 267832 18028 267884 18080
rect 284852 18028 284904 18080
rect 265164 18003 265216 18012
rect 265164 17969 265173 18003
rect 265173 17969 265207 18003
rect 265207 17969 265216 18003
rect 265164 17960 265216 17969
rect 267740 17960 267792 18012
rect 284668 17960 284720 18012
rect 285956 18003 286008 18012
rect 285956 17969 285965 18003
rect 285965 17969 285999 18003
rect 285999 17969 286008 18003
rect 285956 17960 286008 17969
rect 299848 18003 299900 18012
rect 299848 17969 299857 18003
rect 299857 17969 299891 18003
rect 299891 17969 299900 18003
rect 299848 17960 299900 17969
rect 301136 18003 301188 18012
rect 301136 17969 301145 18003
rect 301145 17969 301179 18003
rect 301179 17969 301188 18003
rect 301136 17960 301188 17969
rect 324504 17960 324556 18012
rect 324688 17960 324740 18012
rect 327264 17935 327316 17944
rect 327264 17901 327273 17935
rect 327273 17901 327307 17935
rect 327307 17901 327316 17935
rect 327264 17892 327316 17901
rect 389364 17935 389416 17944
rect 389364 17901 389373 17935
rect 389373 17901 389407 17935
rect 389407 17901 389416 17935
rect 389364 17892 389416 17901
rect 456524 16804 456576 16856
rect 458824 16804 458876 16856
rect 417884 16736 417936 16788
rect 418160 16736 418212 16788
rect 437204 16736 437256 16788
rect 437480 16736 437532 16788
rect 336740 16668 336792 16720
rect 338212 16668 338264 16720
rect 251088 16600 251140 16652
rect 259368 16600 259420 16652
rect 270592 16600 270644 16652
rect 288808 16643 288860 16652
rect 288808 16609 288817 16643
rect 288817 16609 288851 16643
rect 288851 16609 288860 16643
rect 310888 16643 310940 16652
rect 288808 16600 288860 16609
rect 310888 16609 310897 16643
rect 310897 16609 310931 16643
rect 310931 16609 310940 16643
rect 310888 16600 310940 16609
rect 273444 16575 273496 16584
rect 273444 16541 273453 16575
rect 273453 16541 273487 16575
rect 273487 16541 273496 16575
rect 273444 16532 273496 16541
rect 270592 16464 270644 16516
rect 114468 15104 114520 15156
rect 276112 15104 276164 15156
rect 110328 15036 110380 15088
rect 274732 15036 274784 15088
rect 107476 14968 107528 15020
rect 273352 14968 273404 15020
rect 103428 14900 103480 14952
rect 271972 14900 272024 14952
rect 99288 14832 99340 14884
rect 270592 14832 270644 14884
rect 96528 14764 96580 14816
rect 269212 14764 269264 14816
rect 92388 14696 92440 14748
rect 266452 14696 266504 14748
rect 89628 14628 89680 14680
rect 265072 14628 265124 14680
rect 85488 14560 85540 14612
rect 263692 14560 263744 14612
rect 82728 14492 82780 14544
rect 262588 14492 262640 14544
rect 78588 14424 78640 14476
rect 260932 14424 260984 14476
rect 117228 14356 117280 14408
rect 277676 14356 277728 14408
rect 121368 14288 121420 14340
rect 278872 14288 278924 14340
rect 125416 14220 125468 14272
rect 280252 14220 280304 14272
rect 186228 13744 186280 13796
rect 306564 13744 306616 13796
rect 183468 13676 183520 13728
rect 303896 13676 303948 13728
rect 179328 13608 179380 13660
rect 302516 13608 302568 13660
rect 176568 13540 176620 13592
rect 301136 13540 301188 13592
rect 172428 13472 172480 13524
rect 299848 13472 299900 13524
rect 168288 13404 168340 13456
rect 298284 13404 298336 13456
rect 165528 13336 165580 13388
rect 296904 13336 296956 13388
rect 160008 13268 160060 13320
rect 294236 13268 294288 13320
rect 74448 13200 74500 13252
rect 259644 13200 259696 13252
rect 71688 13132 71740 13184
rect 258172 13132 258224 13184
rect 31668 13064 31720 13116
rect 241612 13064 241664 13116
rect 190368 12996 190420 13048
rect 307944 12996 307996 13048
rect 206928 12928 206980 12980
rect 314844 12928 314896 12980
rect 211068 12860 211120 12912
rect 316224 12860 316276 12912
rect 213828 12792 213880 12844
rect 317604 12792 317656 12844
rect 217968 12724 218020 12776
rect 318984 12724 319036 12776
rect 220728 12656 220780 12708
rect 320272 12656 320324 12708
rect 224868 12588 224920 12640
rect 321744 12588 321796 12640
rect 229008 12520 229060 12572
rect 323124 12520 323176 12572
rect 230756 12452 230808 12504
rect 323308 12452 323360 12504
rect 325976 12452 326028 12504
rect 337108 12452 337160 12504
rect 169668 12384 169720 12436
rect 299572 12384 299624 12436
rect 323124 12384 323176 12436
rect 325884 12384 325936 12436
rect 337016 12384 337068 12436
rect 166908 12316 166960 12368
rect 298192 12316 298244 12368
rect 366916 12359 366968 12368
rect 366916 12325 366925 12359
rect 366925 12325 366959 12359
rect 366959 12325 366968 12359
rect 366916 12316 366968 12325
rect 162768 12248 162820 12300
rect 155868 12180 155920 12232
rect 292764 12180 292816 12232
rect 151728 12112 151780 12164
rect 291476 12112 291528 12164
rect 148968 12044 149020 12096
rect 290004 12044 290056 12096
rect 144828 11976 144880 12028
rect 288808 11976 288860 12028
rect 142068 11908 142120 11960
rect 287336 11908 287388 11960
rect 128268 11840 128320 11892
rect 281540 11840 281592 11892
rect 126888 11772 126940 11824
rect 281632 11772 281684 11824
rect 23388 11704 23440 11756
rect 238944 11704 238996 11756
rect 173808 11636 173860 11688
rect 300952 11636 301004 11688
rect 176476 11568 176528 11620
rect 302332 11568 302384 11620
rect 180708 11500 180760 11552
rect 303712 11500 303764 11552
rect 184848 11432 184900 11484
rect 305092 11432 305144 11484
rect 187608 11364 187660 11416
rect 306472 11364 306524 11416
rect 191748 11296 191800 11348
rect 308036 11296 308088 11348
rect 194508 11228 194560 11280
rect 309416 11228 309468 11280
rect 198648 11160 198700 11212
rect 310888 11160 310940 11212
rect 230664 11135 230716 11144
rect 230664 11101 230673 11135
rect 230673 11101 230707 11135
rect 230707 11101 230716 11135
rect 230664 11092 230716 11101
rect 113088 10956 113140 11008
rect 276020 10956 276072 11008
rect 108948 10888 109000 10940
rect 106188 10820 106240 10872
rect 268016 10820 268068 10872
rect 102048 10752 102100 10804
rect 270500 10752 270552 10804
rect 99196 10684 99248 10736
rect 269304 10684 269356 10736
rect 95148 10616 95200 10668
rect 267740 10616 267792 10668
rect 91008 10548 91060 10600
rect 266636 10548 266688 10600
rect 64788 10480 64840 10532
rect 255596 10480 255648 10532
rect 60648 10412 60700 10464
rect 254032 10412 254084 10464
rect 56508 10344 56560 10396
rect 252652 10344 252704 10396
rect 53748 10276 53800 10328
rect 251272 10276 251324 10328
rect 117136 10208 117188 10260
rect 277584 10208 277636 10260
rect 119988 10140 120040 10192
rect 278964 10140 279016 10192
rect 124128 10072 124180 10124
rect 280344 10072 280396 10124
rect 143448 10004 143500 10056
rect 288532 10004 288584 10056
rect 147588 9936 147640 9988
rect 289820 9936 289872 9988
rect 151636 9868 151688 9920
rect 291292 9868 291344 9920
rect 154488 9800 154540 9852
rect 292856 9800 292908 9852
rect 158628 9732 158680 9784
rect 294052 9732 294104 9784
rect 306748 9732 306800 9784
rect 161388 9664 161440 9716
rect 295432 9664 295484 9716
rect 306656 9664 306708 9716
rect 330116 9707 330168 9716
rect 330116 9673 330125 9707
rect 330125 9673 330159 9707
rect 330159 9673 330168 9707
rect 330116 9664 330168 9673
rect 358544 9707 358596 9716
rect 358544 9673 358553 9707
rect 358553 9673 358587 9707
rect 358587 9673 358596 9707
rect 358544 9664 358596 9673
rect 203892 9596 203944 9648
rect 313372 9596 313424 9648
rect 327264 9639 327316 9648
rect 327264 9605 327273 9639
rect 327273 9605 327307 9639
rect 327307 9605 327316 9639
rect 327264 9596 327316 9605
rect 200396 9528 200448 9580
rect 311992 9528 312044 9580
rect 196808 9460 196860 9512
rect 310612 9460 310664 9512
rect 193220 9392 193272 9444
rect 309232 9392 309284 9444
rect 139676 9324 139728 9376
rect 287152 9324 287204 9376
rect 136088 9256 136140 9308
rect 285864 9256 285916 9308
rect 49332 9188 49384 9240
rect 249892 9188 249944 9240
rect 253848 9188 253900 9240
rect 334164 9188 334216 9240
rect 44548 9120 44600 9172
rect 247132 9120 247184 9172
rect 250352 9120 250404 9172
rect 332784 9120 332836 9172
rect 27896 9052 27948 9104
rect 233884 9052 233936 9104
rect 243176 9052 243228 9104
rect 330024 9052 330076 9104
rect 18328 8984 18380 9036
rect 236184 8984 236236 9036
rect 239588 8984 239640 9036
rect 328644 8984 328696 9036
rect 13636 8916 13688 8968
rect 234804 8916 234856 8968
rect 236000 8916 236052 8968
rect 325884 8916 325936 8968
rect 207480 8848 207532 8900
rect 314936 8848 314988 8900
rect 210976 8780 211028 8832
rect 316132 8780 316184 8832
rect 214656 8712 214708 8764
rect 317512 8712 317564 8764
rect 218152 8644 218204 8696
rect 318892 8644 318944 8696
rect 221740 8576 221792 8628
rect 320180 8576 320232 8628
rect 225328 8508 225380 8560
rect 321652 8508 321704 8560
rect 228916 8440 228968 8492
rect 323124 8440 323176 8492
rect 232504 8372 232556 8424
rect 324504 8372 324556 8424
rect 244372 8347 244424 8356
rect 244372 8313 244381 8347
rect 244381 8313 244415 8347
rect 244415 8313 244424 8347
rect 244372 8304 244424 8313
rect 246764 8304 246816 8356
rect 331404 8304 331456 8356
rect 389456 8304 389508 8356
rect 468760 8304 468812 8356
rect 469036 8304 469088 8356
rect 87328 8236 87380 8288
rect 265164 8236 265216 8288
rect 270500 8236 270552 8288
rect 340972 8236 341024 8288
rect 445484 8236 445536 8288
rect 523868 8236 523920 8288
rect 83832 8168 83884 8220
rect 263876 8168 263928 8220
rect 267004 8168 267056 8220
rect 339592 8168 339644 8220
rect 446956 8168 447008 8220
rect 527456 8168 527508 8220
rect 2780 8100 2832 8152
rect 4804 8100 4856 8152
rect 80244 8100 80296 8152
rect 262404 8100 262456 8152
rect 263416 8100 263468 8152
rect 338304 8100 338356 8152
rect 448244 8100 448296 8152
rect 531044 8100 531096 8152
rect 40960 8032 41012 8084
rect 245844 8032 245896 8084
rect 259828 8032 259880 8084
rect 336924 8032 336976 8084
rect 451004 8032 451056 8084
rect 534540 8032 534592 8084
rect 37372 7964 37424 8016
rect 244372 7964 244424 8016
rect 256240 7964 256292 8016
rect 334072 7964 334124 8016
rect 452476 7964 452528 8016
rect 538128 7964 538180 8016
rect 33876 7896 33928 7948
rect 242992 7896 243044 7948
rect 252652 7896 252704 7948
rect 332692 7896 332744 7948
rect 453764 7896 453816 7948
rect 541716 7896 541768 7948
rect 30288 7828 30340 7880
rect 241796 7828 241848 7880
rect 249156 7828 249208 7880
rect 331312 7828 331364 7880
rect 455236 7828 455288 7880
rect 545304 7828 545356 7880
rect 26700 7760 26752 7812
rect 240416 7760 240468 7812
rect 245568 7760 245620 7812
rect 330116 7760 330168 7812
rect 456616 7760 456668 7812
rect 548892 7760 548944 7812
rect 21916 7692 21968 7744
rect 238852 7692 238904 7744
rect 241980 7692 242032 7744
rect 328552 7692 328604 7744
rect 457996 7692 458048 7744
rect 552388 7692 552440 7744
rect 8852 7624 8904 7676
rect 4068 7556 4120 7608
rect 230664 7624 230716 7676
rect 234804 7624 234856 7676
rect 325792 7624 325844 7676
rect 459376 7624 459428 7676
rect 555976 7624 556028 7676
rect 227720 7556 227772 7608
rect 229008 7556 229060 7608
rect 231308 7556 231360 7608
rect 324412 7556 324464 7608
rect 460756 7556 460808 7608
rect 559564 7556 559616 7608
rect 134892 7488 134944 7540
rect 284576 7488 284628 7540
rect 444196 7488 444248 7540
rect 520280 7488 520332 7540
rect 138480 7420 138532 7472
rect 285956 7420 286008 7472
rect 442816 7420 442868 7472
rect 516784 7420 516836 7472
rect 141976 7352 142028 7404
rect 287060 7352 287112 7404
rect 441436 7352 441488 7404
rect 513196 7352 513248 7404
rect 145656 7284 145708 7336
rect 288440 7284 288492 7336
rect 440056 7284 440108 7336
rect 509608 7284 509660 7336
rect 149244 7216 149296 7268
rect 291200 7216 291252 7268
rect 152740 7148 152792 7200
rect 292580 7148 292632 7200
rect 156328 7080 156380 7132
rect 293960 7080 294012 7132
rect 159916 7012 159968 7064
rect 295340 7012 295392 7064
rect 233424 6944 233476 6996
rect 238392 6944 238444 6996
rect 327172 6944 327224 6996
rect 516692 6876 516744 6928
rect 516876 6876 516928 6928
rect 170588 6808 170640 6860
rect 299480 6808 299532 6860
rect 431776 6808 431828 6860
rect 490564 6808 490616 6860
rect 167092 6740 167144 6792
rect 298376 6740 298428 6792
rect 433156 6740 433208 6792
rect 491760 6740 491812 6792
rect 163504 6672 163556 6724
rect 296720 6672 296772 6724
rect 297364 6672 297416 6724
rect 336832 6672 336884 6724
rect 434628 6672 434680 6724
rect 495348 6672 495400 6724
rect 131396 6604 131448 6656
rect 283012 6604 283064 6656
rect 295892 6604 295944 6656
rect 335452 6604 335504 6656
rect 433248 6604 433300 6656
rect 494152 6604 494204 6656
rect 76656 6536 76708 6588
rect 261024 6536 261076 6588
rect 298100 6536 298152 6588
rect 338396 6536 338448 6588
rect 435916 6536 435968 6588
rect 497740 6536 497792 6588
rect 73068 6468 73120 6520
rect 259460 6468 259512 6520
rect 289820 6468 289872 6520
rect 339684 6468 339736 6520
rect 436008 6468 436060 6520
rect 498936 6468 498988 6520
rect 69480 6400 69532 6452
rect 258264 6400 258316 6452
rect 288440 6400 288492 6452
rect 341248 6400 341300 6452
rect 437388 6400 437440 6452
rect 501236 6400 501288 6452
rect 65984 6332 66036 6384
rect 256792 6332 256844 6384
rect 288532 6332 288584 6384
rect 343640 6332 343692 6384
rect 438676 6332 438728 6384
rect 504824 6332 504876 6384
rect 62396 6264 62448 6316
rect 255504 6264 255556 6316
rect 294328 6264 294380 6316
rect 350632 6264 350684 6316
rect 437296 6264 437348 6316
rect 502432 6264 502484 6316
rect 58808 6196 58860 6248
rect 253940 6196 253992 6248
rect 280068 6196 280120 6248
rect 345204 6196 345256 6248
rect 438768 6196 438820 6248
rect 506020 6196 506072 6248
rect 55220 6128 55272 6180
rect 251364 6128 251416 6180
rect 274088 6128 274140 6180
rect 342352 6128 342404 6180
rect 440148 6128 440200 6180
rect 508412 6128 508464 6180
rect 174176 6060 174228 6112
rect 300860 6060 300912 6112
rect 430396 6060 430448 6112
rect 486976 6060 487028 6112
rect 177764 5992 177816 6044
rect 302240 5992 302292 6044
rect 431868 5992 431920 6044
rect 488172 5992 488224 6044
rect 181352 5924 181404 5976
rect 303620 5924 303672 5976
rect 430488 5924 430540 5976
rect 484584 5924 484636 5976
rect 184848 5856 184900 5908
rect 305000 5856 305052 5908
rect 429108 5856 429160 5908
rect 483480 5856 483532 5908
rect 188436 5788 188488 5840
rect 306656 5788 306708 5840
rect 427728 5788 427780 5840
rect 479892 5788 479944 5840
rect 192024 5720 192076 5772
rect 307760 5720 307812 5772
rect 426348 5720 426400 5772
rect 476304 5720 476356 5772
rect 195612 5652 195664 5704
rect 309140 5652 309192 5704
rect 199200 5584 199252 5636
rect 310520 5584 310572 5636
rect 470600 5584 470652 5636
rect 202696 5516 202748 5568
rect 313280 5516 313332 5568
rect 327080 5516 327132 5568
rect 468944 5516 468996 5568
rect 137284 5448 137336 5500
rect 285680 5448 285732 5500
rect 297824 5448 297876 5500
rect 352104 5448 352156 5500
rect 452568 5448 452620 5500
rect 540520 5448 540572 5500
rect 133788 5380 133840 5432
rect 284300 5380 284352 5432
rect 290740 5380 290792 5432
rect 349344 5380 349396 5432
rect 408408 5380 408460 5432
rect 433524 5380 433576 5432
rect 453856 5380 453908 5432
rect 544108 5380 544160 5432
rect 130200 5312 130252 5364
rect 283196 5312 283248 5364
rect 287152 5312 287204 5364
rect 347964 5312 348016 5364
rect 412364 5312 412416 5364
rect 440608 5312 440660 5364
rect 455328 5312 455380 5364
rect 547696 5312 547748 5364
rect 67180 5244 67232 5296
rect 256976 5244 257028 5296
rect 283656 5244 283708 5296
rect 346584 5244 346636 5296
rect 413836 5244 413888 5296
rect 444196 5244 444248 5296
rect 459468 5244 459520 5296
rect 48136 5176 48188 5228
rect 248512 5176 248564 5228
rect 251456 5176 251508 5228
rect 332600 5176 332652 5228
rect 415308 5176 415360 5228
rect 447784 5176 447836 5228
rect 460848 5176 460900 5228
rect 551192 5244 551244 5296
rect 17224 5108 17276 5160
rect 236092 5108 236144 5160
rect 247960 5108 248012 5160
rect 331220 5108 331272 5160
rect 416504 5108 416556 5160
rect 451280 5108 451332 5160
rect 12440 5040 12492 5092
rect 234712 5040 234764 5092
rect 244372 5040 244424 5092
rect 329840 5040 329892 5092
rect 337108 5040 337160 5092
rect 368572 5040 368624 5092
rect 417976 5040 418028 5092
rect 454868 5040 454920 5092
rect 7656 4972 7708 5024
rect 232136 4972 232188 5024
rect 240784 4972 240836 5024
rect 315948 4972 316000 5024
rect 325608 4972 325660 5024
rect 338120 4972 338172 5024
rect 419448 4972 419500 5024
rect 458456 4972 458508 5024
rect 463516 5108 463568 5160
rect 554780 5176 554832 5228
rect 464988 5040 465040 5092
rect 558368 5108 558420 5160
rect 465632 4972 465684 5024
rect 561956 5040 562008 5092
rect 2872 4904 2924 4956
rect 230572 4904 230624 4956
rect 237196 4904 237248 4956
rect 1676 4836 1728 4888
rect 572 4768 624 4820
rect 230480 4836 230532 4888
rect 233700 4836 233752 4888
rect 325700 4836 325752 4888
rect 230112 4768 230164 4820
rect 212264 4700 212316 4752
rect 316040 4700 316092 4752
rect 318708 4700 318760 4752
rect 328736 4904 328788 4956
rect 333612 4904 333664 4956
rect 367192 4904 367244 4956
rect 420736 4904 420788 4956
rect 458088 4904 458140 4956
rect 466184 4904 466236 4956
rect 565544 4972 565596 5024
rect 327080 4836 327132 4888
rect 361672 4836 361724 4888
rect 422208 4836 422260 4888
rect 328460 4768 328512 4820
rect 363052 4768 363104 4820
rect 423588 4768 423640 4820
rect 469128 4836 469180 4888
rect 569040 4904 569092 4956
rect 572628 4836 572680 4888
rect 462136 4768 462188 4820
rect 579804 4768 579856 4820
rect 324320 4700 324372 4752
rect 215852 4632 215904 4684
rect 317420 4632 317472 4684
rect 219348 4564 219400 4616
rect 318800 4564 318852 4616
rect 222936 4496 222988 4548
rect 321560 4632 321612 4684
rect 324228 4632 324280 4684
rect 359004 4700 359056 4752
rect 451096 4700 451148 4752
rect 536932 4700 536984 4752
rect 226524 4428 226576 4480
rect 322940 4564 322992 4616
rect 326528 4632 326580 4684
rect 360476 4632 360528 4684
rect 449808 4632 449860 4684
rect 533436 4632 533488 4684
rect 333980 4564 334032 4616
rect 448336 4564 448388 4616
rect 529848 4564 529900 4616
rect 322848 4496 322900 4548
rect 337016 4496 337068 4548
rect 353484 4496 353536 4548
rect 447048 4496 447100 4548
rect 526260 4496 526312 4548
rect 320364 4428 320416 4480
rect 335360 4428 335412 4480
rect 352564 4428 352616 4480
rect 445576 4428 445628 4480
rect 522672 4428 522724 4480
rect 201500 4360 201552 4412
rect 271144 4360 271196 4412
rect 301412 4360 301464 4412
rect 355324 4360 355376 4412
rect 380164 4360 380216 4412
rect 444288 4360 444340 4412
rect 519084 4360 519136 4412
rect 205088 4292 205140 4344
rect 272524 4292 272576 4344
rect 305000 4292 305052 4344
rect 354956 4292 355008 4344
rect 442908 4292 442960 4344
rect 515588 4292 515640 4344
rect 229100 4224 229152 4276
rect 308588 4224 308640 4276
rect 356152 4224 356204 4276
rect 441528 4224 441580 4276
rect 512000 4224 512052 4276
rect 124220 4156 124272 4208
rect 125416 4156 125468 4208
rect 140872 4156 140924 4208
rect 142068 4156 142120 4208
rect 150440 4156 150492 4208
rect 151636 4156 151688 4208
rect 158720 4156 158772 4208
rect 160008 4156 160060 4208
rect 175372 4156 175424 4208
rect 176568 4156 176620 4208
rect 209872 4156 209924 4208
rect 211068 4156 211120 4208
rect 34980 4088 35032 4140
rect 50344 4088 50396 4140
rect 57612 4088 57664 4140
rect 250444 4088 250496 4140
rect 268108 4088 268160 4140
rect 269028 4088 269080 4140
rect 284760 4088 284812 4140
rect 285588 4088 285640 4140
rect 312084 4156 312136 4208
rect 312176 4156 312228 4208
rect 357808 4156 357860 4208
rect 424968 4156 425020 4208
rect 472716 4156 472768 4208
rect 20720 4020 20772 4072
rect 28264 4020 28316 4072
rect 50528 4020 50580 4072
rect 249064 4020 249116 4072
rect 295892 4088 295944 4140
rect 296720 4088 296772 4140
rect 297916 4088 297968 4140
rect 300308 4088 300360 4140
rect 342904 4088 342956 4140
rect 343640 4088 343692 4140
rect 344284 4088 344336 4140
rect 347872 4088 347924 4140
rect 349068 4088 349120 4140
rect 351368 4088 351420 4140
rect 351828 4088 351880 4140
rect 352564 4088 352616 4140
rect 298100 4020 298152 4072
rect 302608 4020 302660 4072
rect 309784 4020 309836 4072
rect 314568 4020 314620 4072
rect 350632 4020 350684 4072
rect 46940 3952 46992 4004
rect 248696 3952 248748 4004
rect 257436 3952 257488 4004
rect 297364 3952 297416 4004
rect 313372 3952 313424 4004
rect 350540 3952 350592 4004
rect 360936 4088 360988 4140
rect 357440 4020 357492 4072
rect 358084 4020 358136 4072
rect 358176 4020 358228 4072
rect 362224 4020 362276 4072
rect 363328 4088 363380 4140
rect 364248 4088 364300 4140
rect 369216 4088 369268 4140
rect 369768 4088 369820 4140
rect 370412 4088 370464 4140
rect 371148 4088 371200 4140
rect 377588 4088 377640 4140
rect 378048 4088 378100 4140
rect 378784 4088 378836 4140
rect 385316 4088 385368 4140
rect 390836 4088 390888 4140
rect 391848 4088 391900 4140
rect 393136 4088 393188 4140
rect 395436 4088 395488 4140
rect 398104 4088 398156 4140
rect 404912 4088 404964 4140
rect 411076 4088 411128 4140
rect 438216 4088 438268 4140
rect 442264 4088 442316 4140
rect 445668 4088 445720 4140
rect 521476 4088 521528 4140
rect 529204 4088 529256 4140
rect 575020 4088 575072 4140
rect 377404 4020 377456 4072
rect 379980 4020 380032 4072
rect 380808 4020 380860 4072
rect 381176 4020 381228 4072
rect 382188 4020 382240 4072
rect 383568 4020 383620 4072
rect 384304 4020 384356 4072
rect 393228 4020 393280 4072
rect 396632 4020 396684 4072
rect 411168 4020 411220 4072
rect 439412 4020 439464 4072
rect 439504 4020 439556 4072
rect 448428 4020 448480 4072
rect 528652 4020 528704 4072
rect 530584 4020 530636 4072
rect 582196 4020 582248 4072
rect 377128 3952 377180 4004
rect 402796 3952 402848 4004
rect 419172 3952 419224 4004
rect 421564 3952 421616 4004
rect 450176 3952 450228 4004
rect 451188 3952 451240 4004
rect 535736 3952 535788 4004
rect 45744 3884 45796 3936
rect 247684 3884 247736 3936
rect 282460 3884 282512 3936
rect 325608 3884 325660 3936
rect 326436 3884 326488 3936
rect 328460 3884 328512 3936
rect 328828 3884 328880 3936
rect 354128 3884 354180 3936
rect 354220 3884 354272 3936
rect 359096 3884 359148 3936
rect 359740 3884 359792 3936
rect 374092 3884 374144 3936
rect 412456 3884 412508 3936
rect 441804 3884 441856 3936
rect 442356 3884 442408 3936
rect 446312 3884 446364 3936
rect 453672 3884 453724 3936
rect 453948 3884 454000 3936
rect 542912 3884 542964 3936
rect 39764 3816 39816 3868
rect 245936 3816 245988 3868
rect 264612 3816 264664 3868
rect 285956 3816 286008 3868
rect 332416 3816 332468 3868
rect 333244 3816 333296 3868
rect 334716 3816 334768 3868
rect 335268 3816 335320 3868
rect 338764 3816 338816 3868
rect 19524 3748 19576 3800
rect 32404 3748 32456 3800
rect 38568 3748 38620 3800
rect 245752 3748 245804 3800
rect 289544 3748 289596 3800
rect 341524 3816 341576 3868
rect 341892 3816 341944 3868
rect 370136 3816 370188 3868
rect 372804 3816 372856 3868
rect 373908 3816 373960 3868
rect 412548 3816 412600 3868
rect 443000 3816 443052 3868
rect 443644 3816 443696 3868
rect 446588 3816 446640 3868
rect 452476 3816 452528 3868
rect 343088 3748 343140 3800
rect 32680 3680 32732 3732
rect 243084 3680 243136 3732
rect 327632 3680 327684 3732
rect 24308 3612 24360 3664
rect 239036 3612 239088 3664
rect 265808 3612 265860 3664
rect 11244 3544 11296 3596
rect 19984 3544 20036 3596
rect 25504 3544 25556 3596
rect 240324 3544 240376 3596
rect 262220 3544 262272 3596
rect 322848 3612 322900 3664
rect 326528 3612 326580 3664
rect 327724 3544 327776 3596
rect 338304 3680 338356 3732
rect 368664 3748 368716 3800
rect 374000 3748 374052 3800
rect 375288 3748 375340 3800
rect 376392 3748 376444 3800
rect 381636 3748 381688 3800
rect 399484 3748 399536 3800
rect 408500 3748 408552 3800
rect 416688 3748 416740 3800
rect 372712 3680 372764 3732
rect 379704 3680 379756 3732
rect 400036 3680 400088 3732
rect 412088 3680 412140 3732
rect 420368 3680 420420 3732
rect 445392 3748 445444 3800
rect 456708 3748 456760 3800
rect 550088 3816 550140 3868
rect 460296 3748 460348 3800
rect 463240 3748 463292 3800
rect 449164 3680 449216 3732
rect 331312 3612 331364 3664
rect 365812 3612 365864 3664
rect 375196 3612 375248 3664
rect 383844 3612 383896 3664
rect 400128 3612 400180 3664
rect 413192 3612 413244 3664
rect 413928 3612 413980 3664
rect 363604 3544 363656 3596
rect 365720 3544 365772 3596
rect 366916 3544 366968 3596
rect 371608 3544 371660 3596
rect 381544 3544 381596 3596
rect 402888 3544 402940 3596
rect 14832 3476 14884 3528
rect 234896 3476 234948 3528
rect 258632 3476 258684 3528
rect 320364 3476 320416 3528
rect 320456 3476 320508 3528
rect 321468 3476 321520 3528
rect 324044 3476 324096 3528
rect 363144 3476 363196 3528
rect 5264 3408 5316 3460
rect 10324 3408 10376 3460
rect 16028 3408 16080 3460
rect 236276 3408 236328 3460
rect 255044 3408 255096 3460
rect 318708 3408 318760 3460
rect 321652 3408 321704 3460
rect 361856 3408 361908 3460
rect 369124 3476 369176 3528
rect 368020 3408 368072 3460
rect 388260 3476 388312 3528
rect 389088 3476 389140 3528
rect 394608 3476 394660 3528
rect 399024 3476 399076 3528
rect 402244 3476 402296 3528
rect 415676 3544 415728 3596
rect 420276 3612 420328 3664
rect 423956 3612 424008 3664
rect 424416 3612 424468 3664
rect 427084 3612 427136 3664
rect 431132 3612 431184 3664
rect 446496 3612 446548 3664
rect 460204 3680 460256 3732
rect 557172 3748 557224 3800
rect 420828 3544 420880 3596
rect 460848 3544 460900 3596
rect 462228 3544 462280 3596
rect 564348 3680 564400 3732
rect 463608 3612 463660 3664
rect 566740 3612 566792 3664
rect 466368 3544 466420 3596
rect 571432 3544 571484 3596
rect 413284 3476 413336 3528
rect 414480 3476 414532 3528
rect 418068 3476 418120 3528
rect 457260 3476 457312 3528
rect 466276 3476 466328 3528
rect 573824 3476 573876 3528
rect 382372 3408 382424 3460
rect 386604 3408 386656 3460
rect 403624 3408 403676 3460
rect 407304 3408 407356 3460
rect 29092 3340 29144 3392
rect 35164 3340 35216 3392
rect 36176 3340 36228 3392
rect 39304 3340 39356 3392
rect 10048 3272 10100 3324
rect 13084 3272 13136 3324
rect 42156 3272 42208 3324
rect 57244 3272 57296 3324
rect 60004 3340 60056 3392
rect 60648 3340 60700 3392
rect 63592 3340 63644 3392
rect 64788 3340 64840 3392
rect 70676 3340 70728 3392
rect 71688 3340 71740 3392
rect 61384 3272 61436 3324
rect 52828 3204 52880 3256
rect 53748 3204 53800 3256
rect 54024 3204 54076 3256
rect 43352 3136 43404 3188
rect 64788 3204 64840 3256
rect 251824 3340 251876 3392
rect 289820 3340 289872 3392
rect 299112 3340 299164 3392
rect 302884 3340 302936 3392
rect 310980 3340 311032 3392
rect 71872 3272 71924 3324
rect 253204 3272 253256 3324
rect 61200 3136 61252 3188
rect 66904 3068 66956 3120
rect 68284 3136 68336 3188
rect 71044 3068 71096 3120
rect 77852 3204 77904 3256
rect 78588 3204 78640 3256
rect 81440 3204 81492 3256
rect 82728 3204 82780 3256
rect 75460 3136 75512 3188
rect 79324 3136 79376 3188
rect 82636 3136 82688 3188
rect 84844 3204 84896 3256
rect 84936 3204 84988 3256
rect 85488 3204 85540 3256
rect 88524 3204 88576 3256
rect 89628 3204 89680 3256
rect 254584 3204 254636 3256
rect 269304 3204 269356 3256
rect 89720 3068 89772 3120
rect 255964 3136 256016 3188
rect 272892 3136 272944 3188
rect 288440 3272 288492 3324
rect 303804 3272 303856 3324
rect 339500 3272 339552 3324
rect 340788 3272 340840 3324
rect 341156 3340 341208 3392
rect 350540 3340 350592 3392
rect 353668 3340 353720 3392
rect 353760 3340 353812 3392
rect 375656 3340 375708 3392
rect 276480 3204 276532 3256
rect 288532 3204 288584 3256
rect 291936 3204 291988 3256
rect 316684 3204 316736 3256
rect 318064 3204 318116 3256
rect 348424 3272 348476 3324
rect 348976 3272 349028 3324
rect 362132 3272 362184 3324
rect 362868 3272 362920 3324
rect 364524 3272 364576 3324
rect 404268 3340 404320 3392
rect 422760 3408 422812 3460
rect 424324 3408 424376 3460
rect 425152 3408 425204 3460
rect 467932 3408 467984 3460
rect 469036 3408 469088 3460
rect 578608 3408 578660 3460
rect 409788 3340 409840 3392
rect 433984 3340 434036 3392
rect 435824 3340 435876 3392
rect 438124 3340 438176 3392
rect 394516 3272 394568 3324
rect 400220 3272 400272 3324
rect 405004 3272 405056 3324
rect 416872 3272 416924 3324
rect 420184 3272 420236 3324
rect 446588 3272 446640 3324
rect 503628 3272 503680 3324
rect 514024 3340 514076 3392
rect 517888 3340 517940 3392
rect 514392 3272 514444 3324
rect 516876 3272 516928 3324
rect 525064 3340 525116 3392
rect 527824 3340 527876 3392
rect 567844 3340 567896 3392
rect 350264 3204 350316 3256
rect 357256 3204 357308 3256
rect 357348 3204 357400 3256
rect 376024 3204 376076 3256
rect 409144 3204 409196 3256
rect 432328 3204 432380 3256
rect 437020 3204 437072 3256
rect 446220 3204 446272 3256
rect 496544 3204 496596 3256
rect 512644 3204 512696 3256
rect 577412 3272 577464 3324
rect 570236 3204 570288 3256
rect 94504 3068 94556 3120
rect 95148 3068 95200 3120
rect 95700 3068 95752 3120
rect 96528 3068 96580 3120
rect 98092 3068 98144 3120
rect 99196 3068 99248 3120
rect 101588 3068 101640 3120
rect 102048 3068 102100 3120
rect 102784 3068 102836 3120
rect 103428 3068 103480 3120
rect 105176 3068 105228 3120
rect 106188 3068 106240 3120
rect 106372 3068 106424 3120
rect 107476 3068 107528 3120
rect 77944 3000 77996 3052
rect 93308 3000 93360 3052
rect 102600 3000 102652 3052
rect 79048 2932 79100 2984
rect 86132 2932 86184 2984
rect 96896 2932 96948 2984
rect 257344 3068 257396 3120
rect 277676 3068 277728 3120
rect 290464 3136 290516 3188
rect 295524 3136 295576 3188
rect 319444 3136 319496 3188
rect 325240 3136 325292 3188
rect 350540 3136 350592 3188
rect 350632 3136 350684 3188
rect 358912 3136 358964 3188
rect 367284 3136 367336 3188
rect 407028 3136 407080 3188
rect 429936 3136 429988 3188
rect 431224 3136 431276 3188
rect 278872 3068 278924 3120
rect 309784 3068 309836 3120
rect 103980 2864 104032 2916
rect 258816 3000 258868 3052
rect 293132 3000 293184 3052
rect 312544 3000 312596 3052
rect 315764 3000 315816 3052
rect 324228 3000 324280 3052
rect 335912 3000 335964 3052
rect 112352 2932 112404 2984
rect 113088 2932 113140 2984
rect 113548 2932 113600 2984
rect 114468 2932 114520 2984
rect 115940 2932 115992 2984
rect 116952 2932 117004 2984
rect 119436 2932 119488 2984
rect 119988 2932 120040 2984
rect 120632 2932 120684 2984
rect 121368 2932 121420 2984
rect 111156 2864 111208 2916
rect 258724 2932 258776 2984
rect 316960 2932 317012 2984
rect 345664 3068 345716 3120
rect 346676 3068 346728 3120
rect 370504 3068 370556 3120
rect 405648 3068 405700 3120
rect 426348 3068 426400 3120
rect 428464 3068 428516 3120
rect 475108 3068 475160 3120
rect 475384 3068 475436 3120
rect 477500 3068 477552 3120
rect 505744 3136 505796 3188
rect 563152 3136 563204 3188
rect 482284 3068 482336 3120
rect 524972 3068 525024 3120
rect 560760 3068 560812 3120
rect 336096 3000 336148 3052
rect 395896 3000 395948 3052
rect 401324 3000 401376 3052
rect 406384 3000 406436 3052
rect 410892 3000 410944 3052
rect 416596 3000 416648 3052
rect 431316 3000 431368 3052
rect 459652 3000 459704 3052
rect 489368 3000 489420 3052
rect 509884 3000 509936 3052
rect 523684 3000 523736 3052
rect 553584 3000 553636 3052
rect 344376 2932 344428 2984
rect 345480 2932 345532 2984
rect 351184 2932 351236 2984
rect 95884 2796 95936 2848
rect 114744 2796 114796 2848
rect 260104 2864 260156 2916
rect 275284 2864 275336 2916
rect 275928 2864 275980 2916
rect 319260 2864 319312 2916
rect 322848 2864 322900 2916
rect 327080 2864 327132 2916
rect 121828 2796 121880 2848
rect 261484 2796 261536 2848
rect 330024 2796 330076 2848
rect 343640 2796 343692 2848
rect 344560 2864 344612 2916
rect 354956 2932 355008 2984
rect 355968 2932 356020 2984
rect 356060 2932 356112 2984
rect 356704 2932 356756 2984
rect 356796 2932 356848 2984
rect 359464 2932 359516 2984
rect 374368 2932 374420 2984
rect 395988 2932 396040 2984
rect 402520 2932 402572 2984
rect 417424 2932 417476 2984
rect 428740 2932 428792 2984
rect 429844 2932 429896 2984
rect 448980 2932 449032 2984
rect 385868 2864 385920 2916
rect 387064 2864 387116 2916
rect 398196 2864 398248 2916
rect 403716 2864 403768 2916
rect 356060 2796 356112 2848
rect 356152 2796 356204 2848
rect 375840 2796 375892 2848
rect 388444 2796 388496 2848
rect 439596 2796 439648 2848
rect 481088 2932 481140 2984
rect 520924 2932 520976 2984
rect 546500 2932 546552 2984
rect 473912 2864 473964 2916
rect 521016 2864 521068 2916
rect 539324 2864 539376 2916
rect 466828 2796 466880 2848
rect 518164 2796 518216 2848
rect 532240 2796 532292 2848
rect 387064 2728 387116 2780
rect 462044 2728 462096 2780
rect 261024 1232 261076 1284
rect 23112 552 23164 604
rect 23388 552 23440 604
rect 164700 552 164752 604
rect 165528 552 165580 604
rect 165896 552 165948 604
rect 166908 552 166960 604
rect 169392 552 169444 604
rect 169668 552 169720 604
rect 182548 552 182600 604
rect 183468 552 183520 604
rect 183744 552 183796 604
rect 184756 552 184808 604
rect 187240 552 187292 604
rect 187608 552 187660 604
rect 189632 552 189684 604
rect 190368 552 190420 604
rect 281264 552 281316 604
rect 281448 552 281500 604
rect 384672 552 384724 604
rect 384948 552 385000 604
rect 405924 552 405976 604
rect 406108 552 406160 604
rect 463700 552 463752 604
rect 464436 552 464488 604
rect 469220 552 469272 604
rect 470324 552 470376 604
rect 471520 595 471572 604
rect 471520 561 471529 595
rect 471529 561 471563 595
rect 471563 561 471572 595
rect 471520 552 471572 561
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700369 8156 703520
rect 8114 700360 8170 700369
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 105464 700602 105492 703520
rect 137848 700670 137876 703520
rect 154132 700738 154160 703520
rect 170324 700942 170352 703520
rect 202800 701010 202828 703520
rect 202788 701004 202840 701010
rect 202788 700946 202840 700952
rect 170312 700936 170364 700942
rect 170312 700878 170364 700884
rect 154120 700732 154172 700738
rect 154120 700674 154172 700680
rect 137836 700664 137888 700670
rect 137836 700606 137888 700612
rect 105452 700596 105504 700602
rect 105452 700538 105504 700544
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 8114 700295 8170 700304
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 218992 700262 219020 703520
rect 218980 700256 219032 700262
rect 218980 700198 219032 700204
rect 235184 700058 235212 703520
rect 235172 700052 235224 700058
rect 235172 699994 235224 700000
rect 267660 699990 267688 703520
rect 267648 699984 267700 699990
rect 267648 699926 267700 699932
rect 283852 699922 283880 703520
rect 283840 699916 283892 699922
rect 283840 699858 283892 699864
rect 300136 699718 300164 703520
rect 328368 700868 328420 700874
rect 328368 700810 328420 700816
rect 300124 699712 300176 699718
rect 300124 699654 300176 699660
rect 300768 699712 300820 699718
rect 300768 699654 300820 699660
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 300780 584662 300808 699654
rect 321468 696992 321520 696998
rect 321468 696934 321520 696940
rect 320088 673532 320140 673538
rect 320088 673474 320140 673480
rect 315948 650072 316000 650078
rect 315948 650014 316000 650020
rect 313188 626612 313240 626618
rect 313188 626554 313240 626560
rect 309048 603152 309100 603158
rect 309048 603094 309100 603100
rect 300768 584656 300820 584662
rect 300768 584598 300820 584604
rect 298192 583704 298244 583710
rect 298192 583646 298244 583652
rect 256056 583636 256108 583642
rect 256056 583578 256108 583584
rect 245568 583568 245620 583574
rect 245568 583510 245620 583516
rect 6644 583500 6696 583506
rect 6644 583442 6696 583448
rect 4712 583432 4764 583438
rect 4712 583374 4764 583380
rect 3148 583228 3200 583234
rect 3148 583170 3200 583176
rect 3056 568336 3108 568342
rect 3056 568278 3108 568284
rect 3068 567361 3096 568278
rect 3054 567352 3110 567361
rect 3054 567287 3110 567296
rect 3056 553376 3108 553382
rect 3056 553318 3108 553324
rect 3068 553081 3096 553318
rect 3054 553072 3110 553081
rect 3054 553007 3110 553016
rect 3056 538688 3108 538694
rect 3054 538656 3056 538665
rect 3108 538656 3110 538665
rect 3054 538591 3110 538600
rect 3056 510264 3108 510270
rect 3056 510206 3108 510212
rect 3068 509969 3096 510206
rect 3054 509960 3110 509969
rect 3054 509895 3110 509904
rect 2780 495576 2832 495582
rect 2778 495544 2780 495553
rect 2832 495544 2834 495553
rect 2778 495479 2834 495488
rect 2964 481160 3016 481166
rect 2962 481128 2964 481137
rect 3016 481128 3018 481137
rect 2962 481063 3018 481072
rect 3160 452441 3188 583170
rect 3240 583024 3292 583030
rect 3240 582966 3292 582972
rect 3146 452432 3202 452441
rect 3146 452367 3202 452376
rect 3148 438864 3200 438870
rect 3148 438806 3200 438812
rect 3160 438025 3188 438806
rect 3146 438016 3202 438025
rect 3146 437951 3202 437960
rect 3148 424108 3200 424114
rect 3148 424050 3200 424056
rect 3160 423745 3188 424050
rect 3146 423736 3202 423745
rect 3146 423671 3202 423680
rect 3252 395049 3280 582966
rect 4068 582820 4120 582826
rect 4068 582762 4120 582768
rect 3884 582684 3936 582690
rect 3884 582626 3936 582632
rect 3700 582480 3752 582486
rect 3700 582422 3752 582428
rect 3332 578536 3384 578542
rect 3332 578478 3384 578484
rect 3238 395040 3294 395049
rect 3238 394975 3294 394984
rect 3240 380860 3292 380866
rect 3240 380802 3292 380808
rect 3252 380633 3280 380802
rect 3238 380624 3294 380633
rect 3238 380559 3294 380568
rect 3344 366217 3372 578478
rect 3608 578400 3660 578406
rect 3608 578342 3660 578348
rect 3424 578332 3476 578338
rect 3424 578274 3476 578280
rect 3330 366208 3386 366217
rect 3330 366143 3386 366152
rect 3332 324284 3384 324290
rect 3332 324226 3384 324232
rect 3344 323105 3372 324226
rect 3330 323096 3386 323105
rect 3330 323031 3386 323040
rect 2780 308848 2832 308854
rect 2778 308816 2780 308825
rect 2832 308816 2834 308825
rect 2778 308751 2834 308760
rect 2962 295216 3018 295225
rect 2962 295151 3018 295160
rect 2976 294409 3004 295151
rect 2962 294400 3018 294409
rect 2962 294335 3018 294344
rect 2780 252068 2832 252074
rect 2780 252010 2832 252016
rect 2792 251297 2820 252010
rect 2778 251288 2834 251297
rect 2778 251223 2834 251232
rect 3056 237380 3108 237386
rect 3056 237322 3108 237328
rect 3068 237017 3096 237322
rect 3054 237008 3110 237017
rect 3054 236943 3110 236952
rect 2780 165504 2832 165510
rect 2780 165446 2832 165452
rect 2792 165073 2820 165446
rect 2778 165064 2834 165073
rect 2778 164999 2834 165008
rect 3332 151768 3384 151774
rect 3332 151710 3384 151716
rect 3344 150793 3372 151710
rect 3330 150784 3386 150793
rect 3330 150719 3386 150728
rect 2780 136400 2832 136406
rect 2778 136368 2780 136377
rect 2832 136368 2834 136377
rect 2778 136303 2834 136312
rect 2780 122392 2832 122398
rect 2780 122334 2832 122340
rect 2792 122097 2820 122334
rect 2778 122088 2834 122097
rect 2778 122023 2834 122032
rect 3436 93265 3464 578274
rect 3516 578264 3568 578270
rect 3516 578206 3568 578212
rect 3528 107681 3556 578206
rect 3620 179489 3648 578342
rect 3712 193905 3740 582422
rect 3792 579896 3844 579902
rect 3792 579838 3844 579844
rect 3804 208185 3832 579838
rect 3896 222601 3924 582626
rect 3976 578468 4028 578474
rect 3976 578410 4028 578416
rect 3988 265713 4016 578410
rect 4080 280129 4108 582762
rect 4724 495582 4752 583374
rect 6276 583296 6328 583302
rect 4894 583264 4950 583273
rect 6276 583238 6328 583244
rect 4894 583199 4950 583208
rect 4804 581052 4856 581058
rect 4804 580994 4856 581000
rect 4712 495576 4764 495582
rect 4712 495518 4764 495524
rect 4066 280120 4122 280129
rect 4066 280055 4122 280064
rect 3974 265704 4030 265713
rect 3974 265639 4030 265648
rect 3882 222592 3938 222601
rect 3882 222527 3938 222536
rect 3790 208176 3846 208185
rect 3790 208111 3846 208120
rect 3698 193896 3754 193905
rect 3698 193831 3754 193840
rect 3606 179480 3662 179489
rect 3606 179415 3662 179424
rect 3514 107672 3570 107681
rect 3514 107607 3570 107616
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 2780 79892 2832 79898
rect 2780 79834 2832 79840
rect 2792 78985 2820 79834
rect 2778 78976 2834 78985
rect 2778 78911 2834 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 2780 50176 2832 50182
rect 2778 50144 2780 50153
rect 2832 50144 2834 50153
rect 2778 50079 2834 50088
rect 3148 35896 3200 35902
rect 3146 35864 3148 35873
rect 3200 35864 3202 35873
rect 3146 35799 3202 35808
rect 4816 8158 4844 580994
rect 4908 50182 4936 583199
rect 5448 582956 5500 582962
rect 5448 582898 5500 582904
rect 5356 582752 5408 582758
rect 5356 582694 5408 582700
rect 5264 582548 5316 582554
rect 5264 582490 5316 582496
rect 5172 582412 5224 582418
rect 5172 582354 5224 582360
rect 5080 579828 5132 579834
rect 5080 579770 5132 579776
rect 4988 579760 5040 579766
rect 4988 579702 5040 579708
rect 5000 79898 5028 579702
rect 5092 122398 5120 579770
rect 5184 136406 5212 582354
rect 5276 165510 5304 582490
rect 5368 252074 5396 582694
rect 5460 308854 5488 582898
rect 6184 579692 6236 579698
rect 6184 579634 6236 579640
rect 5448 308848 5500 308854
rect 5448 308790 5500 308796
rect 5356 252068 5408 252074
rect 5356 252010 5408 252016
rect 5264 165504 5316 165510
rect 5264 165446 5316 165452
rect 5172 136400 5224 136406
rect 5172 136342 5224 136348
rect 5080 122392 5132 122398
rect 5080 122334 5132 122340
rect 4988 79892 5040 79898
rect 4988 79834 5040 79840
rect 4896 50176 4948 50182
rect 4896 50118 4948 50124
rect 6196 35902 6224 579634
rect 6288 424114 6316 583238
rect 6552 580100 6604 580106
rect 6552 580042 6604 580048
rect 6460 580032 6512 580038
rect 6460 579974 6512 579980
rect 6368 579964 6420 579970
rect 6368 579906 6420 579912
rect 6380 481166 6408 579906
rect 6472 510270 6500 579974
rect 6564 538694 6592 580042
rect 6656 553382 6684 583442
rect 10324 583364 10376 583370
rect 10324 583306 10376 583312
rect 6736 580168 6788 580174
rect 6736 580110 6788 580116
rect 6748 568342 6776 580110
rect 6736 568336 6788 568342
rect 6736 568278 6788 568284
rect 6644 553376 6696 553382
rect 6644 553318 6696 553324
rect 6552 538688 6604 538694
rect 6552 538630 6604 538636
rect 6460 510264 6512 510270
rect 6460 510206 6512 510212
rect 6368 481160 6420 481166
rect 6368 481102 6420 481108
rect 10336 438870 10364 583306
rect 13084 583160 13136 583166
rect 13084 583102 13136 583108
rect 10324 438864 10376 438870
rect 10324 438806 10376 438812
rect 6276 424108 6328 424114
rect 6276 424050 6328 424056
rect 13096 380866 13124 583102
rect 14464 583092 14516 583098
rect 14464 583034 14516 583040
rect 13084 380860 13136 380866
rect 13084 380802 13136 380808
rect 13084 337408 13136 337414
rect 10322 337376 10378 337385
rect 13084 337350 13136 337356
rect 10322 337311 10378 337320
rect 6184 35896 6236 35902
rect 6184 35838 6236 35844
rect 2780 8152 2832 8158
rect 2780 8094 2832 8100
rect 4804 8152 4856 8158
rect 4804 8094 4856 8100
rect 2792 7177 2820 8094
rect 8852 7676 8904 7682
rect 8852 7618 8904 7624
rect 4068 7608 4120 7614
rect 4068 7550 4120 7556
rect 2778 7168 2834 7177
rect 2778 7103 2834 7112
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4830
rect 2884 480 2912 4898
rect 4080 480 4108 7550
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5276 480 5304 3402
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 8864 480 8892 7618
rect 10336 3466 10364 337311
rect 12440 5092 12492 5098
rect 12440 5034 12492 5040
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 10048 3324 10100 3330
rect 10048 3266 10100 3272
rect 10060 480 10088 3266
rect 11256 480 11284 3538
rect 12452 480 12480 5034
rect 13096 3330 13124 337350
rect 14476 324290 14504 583034
rect 15844 582888 15896 582894
rect 15844 582830 15896 582836
rect 14464 324284 14516 324290
rect 14464 324226 14516 324232
rect 15856 237386 15884 582830
rect 17224 582616 17276 582622
rect 17224 582558 17276 582564
rect 24122 582584 24178 582593
rect 15844 237380 15896 237386
rect 15844 237322 15896 237328
rect 17236 151774 17264 582558
rect 24122 582519 24178 582528
rect 19984 337476 20036 337482
rect 19984 337418 20036 337424
rect 17224 151768 17276 151774
rect 17224 151710 17276 151716
rect 18328 9036 18380 9042
rect 18328 8978 18380 8984
rect 13636 8968 13688 8974
rect 13636 8910 13688 8916
rect 13084 3324 13136 3330
rect 13084 3266 13136 3272
rect 13648 480 13676 8910
rect 17224 5160 17276 5166
rect 17224 5102 17276 5108
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14844 480 14872 3470
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 16040 480 16068 3402
rect 17236 480 17264 5102
rect 18340 480 18368 8978
rect 19524 3800 19576 3806
rect 19524 3742 19576 3748
rect 19536 480 19564 3742
rect 19996 3602 20024 337418
rect 24136 64870 24164 582519
rect 245580 579972 245608 583510
rect 247682 582720 247738 582729
rect 247682 582655 247738 582664
rect 247696 579972 247724 582655
rect 256068 579972 256096 583578
rect 293958 583128 294014 583137
rect 293958 583063 294014 583072
rect 289728 581596 289780 581602
rect 289728 581538 289780 581544
rect 287612 581528 287664 581534
rect 287612 581470 287664 581476
rect 283472 581460 283524 581466
rect 283472 581402 283524 581408
rect 281356 581392 281408 581398
rect 281356 581334 281408 581340
rect 275008 581324 275060 581330
rect 275008 581266 275060 581272
rect 268660 581256 268712 581262
rect 268660 581198 268712 581204
rect 264520 581120 264572 581126
rect 264520 581062 264572 581068
rect 262404 580304 262456 580310
rect 262404 580246 262456 580252
rect 262416 579972 262444 580246
rect 264532 579972 264560 581062
rect 268672 579972 268700 581198
rect 275020 579972 275048 581266
rect 281368 579972 281396 581334
rect 283484 579972 283512 581402
rect 287624 579972 287652 581470
rect 289740 579972 289768 581538
rect 293972 579972 294000 583063
rect 296076 581664 296128 581670
rect 296076 581606 296128 581612
rect 296088 579972 296116 581606
rect 298204 579972 298232 583646
rect 302424 581732 302476 581738
rect 302424 581674 302476 581680
rect 300308 580372 300360 580378
rect 300308 580314 300360 580320
rect 300320 579972 300348 580314
rect 302436 579972 302464 581674
rect 304540 581188 304592 581194
rect 304540 581130 304592 581136
rect 304552 579972 304580 581130
rect 306564 580236 306616 580242
rect 306564 580178 306616 580184
rect 306576 579972 306604 580178
rect 309060 579986 309088 603094
rect 311808 592068 311860 592074
rect 311808 592010 311860 592016
rect 311820 580802 311848 592010
rect 311360 580774 311848 580802
rect 311360 579986 311388 580774
rect 313200 579986 313228 626554
rect 315960 580802 315988 650014
rect 317328 638988 317380 638994
rect 317328 638930 317380 638936
rect 315592 580774 315988 580802
rect 315592 580122 315620 580774
rect 315408 580094 315620 580122
rect 315408 579986 315436 580094
rect 317340 579986 317368 638930
rect 308706 579958 309088 579986
rect 310822 579958 311388 579986
rect 312938 579958 313228 579986
rect 315054 579958 315436 579986
rect 317170 579958 317368 579986
rect 320100 579850 320128 673474
rect 321480 579986 321508 696934
rect 324228 685908 324280 685914
rect 324228 685850 324280 685856
rect 324240 579986 324268 685850
rect 325516 584452 325568 584458
rect 325516 584394 325568 584400
rect 321402 579958 321508 579986
rect 323426 579958 324268 579986
rect 325528 579972 325556 584394
rect 328380 580122 328408 700810
rect 329748 700800 329800 700806
rect 329748 700742 329800 700748
rect 328104 580094 328408 580122
rect 328104 579986 328132 580094
rect 327658 579958 328132 579986
rect 329760 579972 329788 700742
rect 332520 699718 332548 703520
rect 336648 700188 336700 700194
rect 336648 700130 336700 700136
rect 335268 700120 335320 700126
rect 335268 700062 335320 700068
rect 332508 699712 332560 699718
rect 332508 699654 332560 699660
rect 331864 584520 331916 584526
rect 331864 584462 331916 584468
rect 331876 579972 331904 584462
rect 335280 580802 335308 700062
rect 334360 580774 335308 580802
rect 334360 579986 334388 580774
rect 336660 579986 336688 700130
rect 343548 699848 343600 699854
rect 343548 699790 343600 699796
rect 340788 699780 340840 699786
rect 340788 699722 340840 699728
rect 338212 584588 338264 584594
rect 338212 584530 338264 584536
rect 334006 579958 334388 579986
rect 336122 579958 336688 579986
rect 338224 579972 338252 584530
rect 340800 579986 340828 699722
rect 343560 580802 343588 699790
rect 348804 699718 348832 703520
rect 364996 703474 365024 703520
rect 364996 703446 365208 703474
rect 358820 701004 358872 701010
rect 358820 700946 358872 700952
rect 356060 700052 356112 700058
rect 356060 699994 356112 700000
rect 351920 699984 351972 699990
rect 351920 699926 351972 699932
rect 346400 699712 346452 699718
rect 346400 699654 346452 699660
rect 347780 699712 347832 699718
rect 347780 699654 347832 699660
rect 348792 699712 348844 699718
rect 348792 699654 348844 699660
rect 344468 584724 344520 584730
rect 344468 584666 344520 584672
rect 343008 580774 343588 580802
rect 343008 579986 343036 580774
rect 340354 579958 340828 579986
rect 342378 579958 343036 579986
rect 344480 579972 344508 584666
rect 346412 579986 346440 699654
rect 346412 579958 346610 579986
rect 319286 579822 320128 579850
rect 347792 579850 347820 699654
rect 350816 584656 350868 584662
rect 350816 584598 350868 584604
rect 350828 579972 350856 584598
rect 351932 580122 351960 699926
rect 354680 699916 354732 699922
rect 354680 699858 354732 699864
rect 351932 580094 352512 580122
rect 352484 579986 352512 580094
rect 354692 579986 354720 699858
rect 356072 580802 356100 699994
rect 356072 580774 356560 580802
rect 356532 579986 356560 580774
rect 358832 579986 358860 700946
rect 362960 700936 363012 700942
rect 362960 700878 363012 700884
rect 360200 700256 360252 700262
rect 360200 700198 360252 700204
rect 360212 580802 360240 700198
rect 360212 580774 360792 580802
rect 360764 579986 360792 580774
rect 362972 579986 363000 700878
rect 364340 700664 364392 700670
rect 364340 700606 364392 700612
rect 364352 580802 364380 700606
rect 365180 687818 365208 703446
rect 367100 700732 367152 700738
rect 367100 700674 367152 700680
rect 364616 687812 364668 687818
rect 364616 687754 364668 687760
rect 365168 687812 365220 687818
rect 365168 687754 365220 687760
rect 364628 685846 364656 687754
rect 364616 685840 364668 685846
rect 364616 685782 364668 685788
rect 364524 676252 364576 676258
rect 364524 676194 364576 676200
rect 364536 669338 364564 676194
rect 364536 669310 364748 669338
rect 364720 650026 364748 669310
rect 364536 649998 364748 650026
rect 364536 630714 364564 649998
rect 364536 630686 364656 630714
rect 364628 618254 364656 630686
rect 364616 618248 364668 618254
rect 364616 618190 364668 618196
rect 364524 608660 364576 608666
rect 364524 608602 364576 608608
rect 364536 601746 364564 608602
rect 364536 601718 364656 601746
rect 364628 598942 364656 601718
rect 364616 598936 364668 598942
rect 364616 598878 364668 598884
rect 364708 589348 364760 589354
rect 364708 589290 364760 589296
rect 364720 584730 364748 589290
rect 364708 584724 364760 584730
rect 364708 584666 364760 584672
rect 364352 580774 365024 580802
rect 364996 579986 365024 580774
rect 367112 579986 367140 700674
rect 368480 700596 368532 700602
rect 368480 700538 368532 700544
rect 368492 580802 368520 700538
rect 374000 700528 374052 700534
rect 374000 700470 374052 700476
rect 371240 700460 371292 700466
rect 371240 700402 371292 700408
rect 368492 580774 369256 580802
rect 369228 579986 369256 580774
rect 352484 579958 352958 579986
rect 354692 579958 355074 579986
rect 356532 579958 357190 579986
rect 358832 579958 359306 579986
rect 360764 579958 361330 579986
rect 362972 579958 363446 579986
rect 364996 579958 365562 579986
rect 367112 579958 367678 579986
rect 369228 579958 369794 579986
rect 371252 579850 371280 700402
rect 374012 579972 374040 700470
rect 375380 700392 375432 700398
rect 375380 700334 375432 700340
rect 378138 700360 378194 700369
rect 375392 580122 375420 700334
rect 378138 700295 378194 700304
rect 379520 700324 379572 700330
rect 375392 580094 375696 580122
rect 375668 579986 375696 580094
rect 378152 579986 378180 700295
rect 379520 700266 379572 700272
rect 379532 580122 379560 700266
rect 397472 699786 397500 703520
rect 413664 699854 413692 703520
rect 413652 699848 413704 699854
rect 413652 699790 413704 699796
rect 397460 699780 397512 699786
rect 397460 699722 397512 699728
rect 429856 688634 429884 703520
rect 462332 700126 462360 703520
rect 478524 700194 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700188 478564 700194
rect 478512 700130 478564 700136
rect 462320 700120 462372 700126
rect 462320 700062 462372 700068
rect 429384 688628 429436 688634
rect 429384 688570 429436 688576
rect 429844 688628 429896 688634
rect 429844 688570 429896 688576
rect 429396 685930 429424 688570
rect 494900 686089 494928 703446
rect 527192 700874 527220 703520
rect 527180 700868 527232 700874
rect 527180 700810 527232 700816
rect 543476 700806 543504 703520
rect 543464 700800 543516 700806
rect 543464 700742 543516 700748
rect 559668 688634 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 559104 688628 559156 688634
rect 559104 688570 559156 688576
rect 559656 688628 559708 688634
rect 559656 688570 559708 688576
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 429304 685902 429424 685930
rect 494242 685944 494298 685953
rect 429304 684486 429332 685902
rect 559116 685930 559144 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 494242 685879 494298 685888
rect 559024 685902 559144 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 429292 684480 429344 684486
rect 429292 684422 429344 684428
rect 382280 681760 382332 681766
rect 382280 681702 382332 681708
rect 379532 580094 379744 580122
rect 379716 579986 379744 580094
rect 382292 579986 382320 681702
rect 494256 678994 494284 685879
rect 559024 684486 559052 685902
rect 580172 685850 580224 685856
rect 559012 684480 559064 684486
rect 559012 684422 559064 684428
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 386420 667956 386472 667962
rect 386420 667898 386472 667904
rect 383660 652792 383712 652798
rect 383660 652734 383712 652740
rect 375668 579958 376142 579986
rect 378152 579958 378258 579986
rect 379716 579958 380282 579986
rect 382292 579958 382398 579986
rect 383672 579850 383700 652734
rect 386432 579986 386460 667898
rect 429660 666596 429712 666602
rect 429660 666538 429712 666544
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 429672 659682 429700 666538
rect 429488 659654 429700 659682
rect 494164 659682 494192 666538
rect 559392 659682 559420 666538
rect 494164 659654 494284 659682
rect 429488 647290 429516 659654
rect 494256 654158 494284 659654
rect 559208 659654 559420 659682
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 429384 647284 429436 647290
rect 429384 647226 429436 647232
rect 429476 647284 429528 647290
rect 429476 647226 429528 647232
rect 429396 640422 429424 647226
rect 494072 644450 494100 654094
rect 559208 647290 559236 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 494072 644422 494284 644450
rect 429384 640416 429436 640422
rect 429384 640358 429436 640364
rect 429476 640416 429528 640422
rect 429476 640358 429528 640364
rect 429488 630698 429516 640358
rect 494256 634846 494284 644422
rect 559116 640422 559144 647226
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 429292 630692 429344 630698
rect 429292 630634 429344 630640
rect 429476 630692 429528 630698
rect 429476 630634 429528 630640
rect 429304 630578 429332 630634
rect 429304 630550 429424 630578
rect 387800 623824 387852 623830
rect 387800 623766 387852 623772
rect 387812 580122 387840 623766
rect 429396 621058 429424 630550
rect 494072 625138 494100 634782
rect 559208 630698 559236 640358
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 559024 630578 559052 630634
rect 559024 630550 559144 630578
rect 494072 625110 494284 625138
rect 429396 621030 429516 621058
rect 429488 611386 429516 621030
rect 494256 615534 494284 625110
rect 559116 621058 559144 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 559116 621030 559236 621058
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 429292 611380 429344 611386
rect 429292 611322 429344 611328
rect 429476 611380 429528 611386
rect 429476 611322 429528 611328
rect 429304 611266 429332 611322
rect 429304 611238 429424 611266
rect 391940 610020 391992 610026
rect 391940 609962 391992 609968
rect 390560 594856 390612 594862
rect 390560 594798 390612 594804
rect 387812 580094 388392 580122
rect 388364 579986 388392 580094
rect 390572 579986 390600 594798
rect 391952 580802 391980 609962
rect 429396 608598 429424 611238
rect 429384 608592 429436 608598
rect 429384 608534 429436 608540
rect 494072 605826 494100 615470
rect 559208 611386 559236 621030
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 559024 611266 559052 611322
rect 559024 611238 559144 611266
rect 559116 608598 559144 611238
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 494072 605798 494284 605826
rect 429568 601724 429620 601730
rect 429568 601666 429620 601672
rect 429580 598942 429608 601666
rect 429568 598936 429620 598942
rect 429568 598878 429620 598884
rect 494256 596222 494284 605798
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 559300 598942 559328 601666
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 494072 596142 494192 596158
rect 494164 596034 494192 596142
rect 494164 596006 494284 596034
rect 429660 589348 429712 589354
rect 429660 589290 429712 589296
rect 429672 584594 429700 589290
rect 429660 584588 429712 584594
rect 429660 584530 429712 584536
rect 494256 584526 494284 596006
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 494244 584520 494296 584526
rect 494244 584462 494296 584468
rect 559392 584458 559420 589290
rect 559380 584452 559432 584458
rect 559380 584394 559432 584400
rect 471244 583704 471296 583710
rect 471244 583646 471296 583652
rect 399208 583500 399260 583506
rect 399208 583442 399260 583448
rect 391952 580774 392440 580802
rect 392412 579986 392440 580774
rect 395068 580168 395120 580174
rect 395068 580110 395120 580116
rect 386432 579958 386630 579986
rect 388364 579958 388746 579986
rect 390572 579958 390862 579986
rect 392412 579958 392978 579986
rect 395080 579972 395108 580110
rect 397092 580100 397144 580106
rect 397092 580042 397144 580048
rect 397104 579972 397132 580042
rect 399220 579972 399248 583442
rect 405556 583432 405608 583438
rect 405556 583374 405608 583380
rect 400956 580032 401008 580038
rect 401008 579980 401350 579986
rect 400956 579974 401350 579980
rect 400968 579958 401350 579974
rect 403176 579970 403466 579986
rect 405568 579972 405596 583374
rect 411904 583364 411956 583370
rect 411904 583306 411956 583312
rect 409788 583296 409840 583302
rect 409788 583238 409840 583244
rect 407672 583228 407724 583234
rect 407672 583170 407724 583176
rect 407684 579972 407712 583170
rect 409800 579972 409828 583238
rect 411916 579972 411944 583306
rect 460294 583264 460350 583273
rect 460294 583199 460350 583208
rect 418160 583160 418212 583166
rect 418160 583102 418212 583108
rect 414020 583024 414072 583030
rect 414020 582966 414072 582972
rect 414032 579972 414060 582966
rect 418172 579972 418200 583102
rect 424508 583092 424560 583098
rect 424508 583034 424560 583040
rect 420274 582992 420330 583001
rect 420274 582927 420330 582936
rect 422392 582956 422444 582962
rect 420288 579972 420316 582927
rect 422392 582898 422444 582904
rect 422404 579972 422432 582898
rect 424520 579972 424548 583034
rect 437112 582888 437164 582894
rect 426622 582856 426678 582865
rect 437112 582830 437164 582836
rect 426622 582791 426678 582800
rect 430856 582820 430908 582826
rect 426636 579972 426664 582791
rect 430856 582762 430908 582768
rect 430868 579972 430896 582762
rect 432972 582752 433024 582758
rect 432972 582694 433024 582700
rect 432984 579972 433012 582694
rect 434996 582684 435048 582690
rect 434996 582626 435048 582632
rect 435008 579972 435036 582626
rect 437124 579972 437152 582830
rect 449808 582616 449860 582622
rect 449808 582558 449860 582564
rect 445576 582548 445628 582554
rect 445576 582490 445628 582496
rect 443460 582480 443512 582486
rect 443460 582422 443512 582428
rect 443472 579972 443500 582422
rect 445588 579972 445616 582490
rect 447692 582412 447744 582418
rect 447692 582354 447744 582360
rect 447704 579972 447732 582354
rect 449820 579972 449848 582558
rect 460308 579972 460336 583199
rect 462410 582584 462466 582593
rect 462410 582519 462466 582528
rect 462424 579972 462452 582519
rect 469588 581732 469640 581738
rect 469588 581674 469640 581680
rect 466644 581052 466696 581058
rect 466644 580994 466696 581000
rect 466656 579972 466684 580994
rect 403164 579964 403466 579970
rect 403216 579958 403466 579964
rect 403164 579906 403216 579912
rect 438860 579896 438912 579902
rect 347792 579822 348726 579850
rect 371252 579822 371910 579850
rect 383672 579822 384514 579850
rect 438912 579844 439254 579850
rect 438860 579838 439254 579844
rect 438872 579822 439254 579838
rect 451568 579834 451950 579850
rect 451556 579828 451950 579834
rect 451608 579822 451950 579828
rect 451556 579770 451608 579776
rect 458272 579760 458324 579766
rect 458206 579708 458272 579714
rect 458206 579702 458324 579708
rect 458206 579686 458312 579702
rect 464264 579698 464554 579714
rect 464252 579692 464554 579698
rect 464304 579686 464554 579692
rect 464252 579634 464304 579640
rect 270802 579426 271184 579442
rect 415688 579426 416070 579442
rect 428384 579426 428766 579442
rect 453592 579426 453974 579442
rect 455800 579426 456090 579442
rect 270802 579420 271196 579426
rect 270802 579414 271144 579420
rect 271144 579362 271196 579368
rect 415676 579420 416070 579426
rect 415728 579414 416070 579420
rect 428372 579420 428766 579426
rect 415676 579362 415728 579368
rect 428424 579414 428766 579420
rect 453580 579420 453974 579426
rect 428372 579362 428424 579368
rect 453632 579414 453974 579420
rect 455788 579420 456090 579426
rect 453580 579362 453632 579368
rect 455840 579414 456090 579420
rect 455788 579362 455840 579368
rect 252100 579352 252152 579358
rect 231122 579320 231178 579329
rect 230874 579278 231122 579306
rect 232962 579320 233018 579329
rect 232898 579278 232962 579306
rect 231122 579255 231178 579264
rect 235262 579320 235318 579329
rect 235014 579278 235262 579306
rect 232962 579255 233018 579264
rect 237194 579320 237250 579329
rect 237130 579278 237194 579306
rect 235262 579255 235318 579264
rect 239402 579320 239458 579329
rect 239246 579278 239402 579306
rect 237194 579255 237250 579264
rect 241426 579320 241482 579329
rect 241362 579278 241426 579306
rect 239402 579255 239458 579264
rect 241426 579255 241482 579264
rect 243266 579320 243322 579329
rect 249522 579320 249578 579329
rect 243322 579278 243478 579306
rect 243266 579255 243322 579264
rect 249578 579278 249734 579306
rect 251850 579300 252100 579306
rect 254216 579352 254268 579358
rect 251850 579294 252152 579300
rect 253966 579300 254216 579306
rect 258448 579352 258500 579358
rect 253966 579294 254268 579300
rect 258198 579300 258448 579306
rect 260656 579352 260708 579358
rect 258198 579294 258500 579300
rect 260314 579300 260656 579306
rect 266912 579352 266964 579358
rect 260314 579294 260708 579300
rect 266662 579300 266912 579306
rect 273076 579352 273128 579358
rect 266662 579294 266964 579300
rect 272918 579300 273076 579306
rect 277308 579352 277360 579358
rect 272918 579294 273128 579300
rect 277150 579300 277308 579306
rect 279608 579352 279660 579358
rect 277150 579294 277360 579300
rect 279266 579300 279608 579306
rect 285680 579352 285732 579358
rect 279266 579294 279660 579300
rect 285614 579300 285680 579306
rect 292120 579352 292172 579358
rect 285614 579294 285732 579300
rect 291870 579300 292120 579306
rect 291870 579294 292172 579300
rect 441068 579352 441120 579358
rect 468574 579320 468630 579329
rect 441120 579300 441370 579306
rect 441068 579294 441370 579300
rect 251850 579278 252140 579294
rect 253966 579278 254256 579294
rect 258198 579278 258488 579294
rect 260314 579278 260696 579294
rect 266662 579278 266952 579294
rect 272918 579278 273116 579294
rect 277150 579278 277348 579294
rect 279266 579278 279648 579294
rect 285614 579278 285720 579294
rect 291870 579278 292160 579294
rect 441080 579278 441370 579294
rect 249522 579255 249578 579264
rect 468630 579278 468786 579306
rect 468574 579255 468630 579264
rect 469600 557530 469628 581674
rect 469772 581664 469824 581670
rect 469772 581606 469824 581612
rect 469680 580372 469732 580378
rect 469680 580314 469732 580320
rect 469588 557524 469640 557530
rect 469588 557466 469640 557472
rect 469692 534070 469720 580314
rect 469680 534064 469732 534070
rect 469680 534006 469732 534012
rect 469784 510610 469812 581606
rect 470508 581596 470560 581602
rect 470508 581538 470560 581544
rect 470416 581528 470468 581534
rect 470416 581470 470468 581476
rect 470324 581460 470376 581466
rect 470324 581402 470376 581408
rect 470232 581392 470284 581398
rect 470232 581334 470284 581340
rect 470140 581324 470192 581330
rect 470140 581266 470192 581272
rect 469956 581256 470008 581262
rect 469956 581198 470008 581204
rect 469864 580304 469916 580310
rect 469864 580246 469916 580252
rect 469772 510604 469824 510610
rect 469772 510546 469824 510552
rect 231044 340190 231426 340218
rect 232516 340190 232898 340218
rect 244752 340190 245226 340218
rect 290292 340190 290766 340218
rect 291764 340190 292238 340218
rect 294708 340190 295182 340218
rect 300136 340190 300518 340218
rect 325068 340190 325542 340218
rect 327552 340190 327934 340218
rect 337396 340190 337778 340218
rect 340340 340190 340722 340218
rect 374564 340190 375038 340218
rect 386800 340190 387274 340218
rect 392610 340190 393084 340218
rect 399510 340190 399892 340218
rect 422970 340190 423444 340218
rect 229112 340054 230046 340082
rect 71044 338088 71096 338094
rect 71044 338030 71096 338036
rect 66904 338020 66956 338026
rect 66904 337962 66956 337968
rect 61384 337952 61436 337958
rect 61384 337894 61436 337900
rect 57244 337884 57296 337890
rect 57244 337826 57296 337832
rect 50344 337816 50396 337822
rect 50344 337758 50396 337764
rect 32404 337748 32456 337754
rect 32404 337690 32456 337696
rect 28264 337544 28316 337550
rect 28264 337486 28316 337492
rect 24124 64864 24176 64870
rect 24124 64806 24176 64812
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 21916 7744 21968 7750
rect 21916 7686 21968 7692
rect 20720 4072 20772 4078
rect 20720 4014 20772 4020
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 20732 480 20760 4014
rect 21928 480 21956 7686
rect 23400 610 23428 11698
rect 27896 9104 27948 9110
rect 27896 9046 27948 9052
rect 26700 7812 26752 7818
rect 26700 7754 26752 7760
rect 24308 3664 24360 3670
rect 24308 3606 24360 3612
rect 23112 604 23164 610
rect 23112 546 23164 552
rect 23388 604 23440 610
rect 23388 546 23440 552
rect 23124 480 23152 546
rect 24320 480 24348 3606
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25516 480 25544 3538
rect 26712 480 26740 7754
rect 27908 480 27936 9046
rect 28276 4078 28304 337486
rect 31668 13116 31720 13122
rect 31668 13058 31720 13064
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 28264 4072 28316 4078
rect 28264 4014 28316 4020
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 29104 480 29132 3334
rect 30300 480 30328 7822
rect 31680 626 31708 13058
rect 32416 3806 32444 337690
rect 39304 337680 39356 337686
rect 39304 337622 39356 337628
rect 35164 337612 35216 337618
rect 35164 337554 35216 337560
rect 33876 7948 33928 7954
rect 33876 7890 33928 7896
rect 32404 3800 32456 3806
rect 32404 3742 32456 3748
rect 32680 3732 32732 3738
rect 32680 3674 32732 3680
rect 31496 598 31708 626
rect 31496 480 31524 598
rect 32692 480 32720 3674
rect 33888 480 33916 7890
rect 34980 4140 35032 4146
rect 34980 4082 35032 4088
rect 34992 480 35020 4082
rect 35176 3398 35204 337554
rect 37372 8016 37424 8022
rect 37372 7958 37424 7964
rect 35164 3392 35216 3398
rect 35164 3334 35216 3340
rect 36176 3392 36228 3398
rect 36176 3334 36228 3340
rect 36188 480 36216 3334
rect 37384 480 37412 7958
rect 38568 3800 38620 3806
rect 38568 3742 38620 3748
rect 38580 480 38608 3742
rect 39316 3398 39344 337622
rect 49332 9240 49384 9246
rect 49332 9182 49384 9188
rect 44548 9172 44600 9178
rect 44548 9114 44600 9120
rect 40960 8084 41012 8090
rect 40960 8026 41012 8032
rect 39764 3868 39816 3874
rect 39764 3810 39816 3816
rect 39304 3392 39356 3398
rect 39304 3334 39356 3340
rect 39776 480 39804 3810
rect 40972 480 41000 8026
rect 42156 3324 42208 3330
rect 42156 3266 42208 3272
rect 42168 480 42196 3266
rect 43352 3188 43404 3194
rect 43352 3130 43404 3136
rect 43364 480 43392 3130
rect 44560 480 44588 9114
rect 48136 5228 48188 5234
rect 48136 5170 48188 5176
rect 46940 4004 46992 4010
rect 46940 3946 46992 3952
rect 45744 3936 45796 3942
rect 45744 3878 45796 3884
rect 45756 480 45784 3878
rect 46952 480 46980 3946
rect 48148 480 48176 5170
rect 49344 480 49372 9182
rect 50356 4146 50384 337758
rect 56508 10396 56560 10402
rect 56508 10338 56560 10344
rect 53748 10328 53800 10334
rect 53748 10270 53800 10276
rect 51630 6216 51686 6225
rect 51630 6151 51686 6160
rect 50344 4140 50396 4146
rect 50344 4082 50396 4088
rect 50528 4072 50580 4078
rect 50528 4014 50580 4020
rect 50540 480 50568 4014
rect 51644 480 51672 6151
rect 53760 3262 53788 10270
rect 55220 6180 55272 6186
rect 55220 6122 55272 6128
rect 52828 3256 52880 3262
rect 52828 3198 52880 3204
rect 53748 3256 53800 3262
rect 53748 3198 53800 3204
rect 54024 3256 54076 3262
rect 54024 3198 54076 3204
rect 52840 480 52868 3198
rect 54036 480 54064 3198
rect 55232 480 55260 6122
rect 56520 3482 56548 10338
rect 56428 3454 56548 3482
rect 56428 480 56456 3454
rect 57256 3330 57284 337826
rect 60648 10464 60700 10470
rect 60648 10406 60700 10412
rect 58808 6248 58860 6254
rect 58808 6190 58860 6196
rect 57612 4140 57664 4146
rect 57612 4082 57664 4088
rect 57244 3324 57296 3330
rect 57244 3266 57296 3272
rect 57624 480 57652 4082
rect 58820 480 58848 6190
rect 60660 3398 60688 10406
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60016 480 60044 3334
rect 61396 3330 61424 337894
rect 64788 10532 64840 10538
rect 64788 10474 64840 10480
rect 62396 6316 62448 6322
rect 62396 6258 62448 6264
rect 61384 3324 61436 3330
rect 61384 3266 61436 3272
rect 61200 3188 61252 3194
rect 61200 3130 61252 3136
rect 61212 480 61240 3130
rect 62408 480 62436 6258
rect 64800 3398 64828 10474
rect 65984 6384 66036 6390
rect 65984 6326 66036 6332
rect 63592 3392 63644 3398
rect 63592 3334 63644 3340
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 63604 480 63632 3334
rect 64788 3256 64840 3262
rect 64788 3198 64840 3204
rect 64800 480 64828 3198
rect 65996 480 66024 6326
rect 66916 3126 66944 337962
rect 69480 6452 69532 6458
rect 69480 6394 69532 6400
rect 67180 5296 67232 5302
rect 67180 5238 67232 5244
rect 66904 3120 66956 3126
rect 66904 3062 66956 3068
rect 67192 480 67220 5238
rect 68284 3188 68336 3194
rect 68284 3130 68336 3136
rect 68296 480 68324 3130
rect 69492 480 69520 6394
rect 70676 3392 70728 3398
rect 70676 3334 70728 3340
rect 70688 480 70716 3334
rect 71056 3126 71084 338030
rect 79324 337340 79376 337346
rect 79324 337282 79376 337288
rect 77944 337000 77996 337006
rect 77944 336942 77996 336948
rect 74448 13252 74500 13258
rect 74448 13194 74500 13200
rect 71688 13184 71740 13190
rect 71688 13126 71740 13132
rect 71700 3398 71728 13126
rect 73068 6520 73120 6526
rect 73068 6462 73120 6468
rect 71688 3392 71740 3398
rect 71688 3334 71740 3340
rect 71872 3324 71924 3330
rect 71872 3266 71924 3272
rect 71044 3120 71096 3126
rect 71044 3062 71096 3068
rect 71884 480 71912 3266
rect 73080 480 73108 6462
rect 74460 3380 74488 13194
rect 76656 6588 76708 6594
rect 76656 6530 76708 6536
rect 74276 3352 74488 3380
rect 74276 480 74304 3352
rect 75460 3188 75512 3194
rect 75460 3130 75512 3136
rect 75472 480 75500 3130
rect 76668 480 76696 6530
rect 77852 3256 77904 3262
rect 77852 3198 77904 3204
rect 77864 480 77892 3198
rect 77956 3058 77984 336942
rect 78588 14476 78640 14482
rect 78588 14418 78640 14424
rect 78600 3262 78628 14418
rect 78588 3256 78640 3262
rect 78588 3198 78640 3204
rect 79336 3194 79364 337282
rect 132500 337272 132552 337278
rect 132498 337240 132500 337249
rect 142068 337272 142120 337278
rect 132552 337240 132554 337249
rect 84844 337204 84896 337210
rect 132498 337175 132554 337184
rect 142066 337240 142068 337249
rect 151820 337272 151872 337278
rect 142120 337240 142122 337249
rect 142066 337175 142122 337184
rect 151818 337240 151820 337249
rect 161388 337272 161440 337278
rect 151872 337240 151874 337249
rect 151818 337175 151874 337184
rect 161386 337240 161388 337249
rect 171140 337272 171192 337278
rect 161440 337240 161442 337249
rect 161386 337175 161442 337184
rect 171138 337240 171140 337249
rect 180708 337272 180760 337278
rect 171192 337240 171194 337249
rect 171138 337175 171194 337184
rect 180706 337240 180708 337249
rect 190460 337272 190512 337278
rect 180760 337240 180762 337249
rect 180706 337175 180762 337184
rect 190458 337240 190460 337249
rect 200028 337272 200080 337278
rect 190512 337240 190514 337249
rect 190458 337175 190514 337184
rect 200026 337240 200028 337249
rect 209780 337272 209832 337278
rect 200080 337240 200082 337249
rect 200026 337175 200082 337184
rect 209778 337240 209780 337249
rect 219348 337272 219400 337278
rect 209832 337240 209834 337249
rect 209778 337175 209834 337184
rect 219346 337240 219348 337249
rect 219400 337240 219402 337249
rect 219346 337175 219402 337184
rect 84844 337146 84896 337152
rect 82728 14544 82780 14550
rect 82728 14486 82780 14492
rect 80244 8152 80296 8158
rect 80244 8094 80296 8100
rect 79324 3188 79376 3194
rect 79324 3130 79376 3136
rect 77944 3052 77996 3058
rect 77944 2994 77996 3000
rect 79048 2984 79100 2990
rect 79048 2926 79100 2932
rect 79060 480 79088 2926
rect 80256 480 80284 8094
rect 82740 3262 82768 14486
rect 83832 8220 83884 8226
rect 83832 8162 83884 8168
rect 81440 3256 81492 3262
rect 81440 3198 81492 3204
rect 82728 3256 82780 3262
rect 82728 3198 82780 3204
rect 81452 480 81480 3198
rect 82636 3188 82688 3194
rect 82636 3130 82688 3136
rect 82648 480 82676 3130
rect 83844 480 83872 8162
rect 84856 3262 84884 337146
rect 100668 337136 100720 337142
rect 100668 337078 100720 337084
rect 95884 337068 95936 337074
rect 95884 337010 95936 337016
rect 92388 14748 92440 14754
rect 92388 14690 92440 14696
rect 89628 14680 89680 14686
rect 89628 14622 89680 14628
rect 85488 14612 85540 14618
rect 85488 14554 85540 14560
rect 85500 3262 85528 14554
rect 87328 8288 87380 8294
rect 87328 8230 87380 8236
rect 84844 3256 84896 3262
rect 84844 3198 84896 3204
rect 84936 3256 84988 3262
rect 84936 3198 84988 3204
rect 85488 3256 85540 3262
rect 85488 3198 85540 3204
rect 84948 480 84976 3198
rect 86132 2984 86184 2990
rect 86132 2926 86184 2932
rect 86144 480 86172 2926
rect 87340 480 87368 8230
rect 89640 3262 89668 14622
rect 91008 10600 91060 10606
rect 91008 10542 91060 10548
rect 91020 3482 91048 10542
rect 92400 3482 92428 14690
rect 95148 10668 95200 10674
rect 95148 10610 95200 10616
rect 90928 3454 91048 3482
rect 92124 3454 92428 3482
rect 88524 3256 88576 3262
rect 88524 3198 88576 3204
rect 89628 3256 89680 3262
rect 89628 3198 89680 3204
rect 88536 480 88564 3198
rect 89720 3120 89772 3126
rect 89720 3062 89772 3068
rect 89732 480 89760 3062
rect 90928 480 90956 3454
rect 92124 480 92152 3454
rect 95160 3126 95188 10610
rect 94504 3120 94556 3126
rect 94504 3062 94556 3068
rect 95148 3120 95200 3126
rect 95148 3062 95200 3068
rect 95700 3120 95752 3126
rect 95700 3062 95752 3068
rect 93308 3052 93360 3058
rect 93308 2994 93360 3000
rect 93320 480 93348 2994
rect 94516 480 94544 3062
rect 95712 480 95740 3062
rect 95896 2854 95924 337010
rect 99288 14884 99340 14890
rect 99288 14826 99340 14832
rect 96528 14816 96580 14822
rect 96528 14758 96580 14764
rect 96540 3126 96568 14758
rect 99196 10736 99248 10742
rect 99196 10678 99248 10684
rect 99208 3126 99236 10678
rect 96528 3120 96580 3126
rect 96528 3062 96580 3068
rect 98092 3120 98144 3126
rect 98092 3062 98144 3068
rect 99196 3120 99248 3126
rect 99196 3062 99248 3068
rect 96896 2984 96948 2990
rect 96896 2926 96948 2932
rect 95884 2848 95936 2854
rect 95884 2790 95936 2796
rect 96908 480 96936 2926
rect 98104 480 98132 3062
rect 99300 480 99328 14826
rect 100680 3482 100708 337078
rect 107568 337000 107620 337006
rect 107568 336942 107620 336948
rect 102784 336932 102836 336938
rect 102784 336874 102836 336880
rect 102048 10804 102100 10810
rect 102048 10746 102100 10752
rect 100496 3454 100708 3482
rect 100496 480 100524 3454
rect 102060 3126 102088 10746
rect 102796 3210 102824 336874
rect 107476 15020 107528 15026
rect 107476 14962 107528 14968
rect 103428 14952 103480 14958
rect 103428 14894 103480 14900
rect 102612 3182 102824 3210
rect 101588 3120 101640 3126
rect 101588 3062 101640 3068
rect 102048 3120 102100 3126
rect 102048 3062 102100 3068
rect 101600 480 101628 3062
rect 102612 3058 102640 3182
rect 103440 3126 103468 14894
rect 106188 10872 106240 10878
rect 106188 10814 106240 10820
rect 106200 3126 106228 10814
rect 107488 3126 107516 14962
rect 102784 3120 102836 3126
rect 102784 3062 102836 3068
rect 103428 3120 103480 3126
rect 103428 3062 103480 3068
rect 105176 3120 105228 3126
rect 105176 3062 105228 3068
rect 106188 3120 106240 3126
rect 106188 3062 106240 3068
rect 106372 3120 106424 3126
rect 106372 3062 106424 3068
rect 107476 3120 107528 3126
rect 107476 3062 107528 3068
rect 102600 3052 102652 3058
rect 102600 2994 102652 3000
rect 102796 480 102824 3062
rect 103980 2916 104032 2922
rect 103980 2858 104032 2864
rect 103992 480 104020 2858
rect 105188 480 105216 3062
rect 106384 480 106412 3062
rect 107580 480 107608 336942
rect 118608 336864 118660 336870
rect 118608 336806 118660 336812
rect 114468 15156 114520 15162
rect 114468 15098 114520 15104
rect 110328 15088 110380 15094
rect 110328 15030 110380 15036
rect 108948 10940 109000 10946
rect 108948 10882 109000 10888
rect 108960 3482 108988 10882
rect 110340 3482 110368 15030
rect 113088 11008 113140 11014
rect 113088 10950 113140 10956
rect 108776 3454 108988 3482
rect 109972 3454 110368 3482
rect 108776 480 108804 3454
rect 109972 480 110000 3454
rect 113100 2990 113128 10950
rect 114480 2990 114508 15098
rect 117228 14408 117280 14414
rect 117228 14350 117280 14356
rect 117136 10260 117188 10266
rect 117136 10202 117188 10208
rect 117148 3618 117176 10202
rect 116964 3590 117176 3618
rect 116964 2990 116992 3590
rect 117240 3482 117268 14350
rect 117148 3454 117268 3482
rect 112352 2984 112404 2990
rect 112352 2926 112404 2932
rect 113088 2984 113140 2990
rect 113088 2926 113140 2932
rect 113548 2984 113600 2990
rect 113548 2926 113600 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 115940 2984 115992 2990
rect 115940 2926 115992 2932
rect 116952 2984 117004 2990
rect 116952 2926 117004 2932
rect 111156 2916 111208 2922
rect 111156 2858 111208 2864
rect 111168 480 111196 2858
rect 112364 480 112392 2926
rect 113560 480 113588 2926
rect 114744 2848 114796 2854
rect 114744 2790 114796 2796
rect 114756 480 114784 2790
rect 115952 480 115980 2926
rect 117148 480 117176 3454
rect 118620 3346 118648 336806
rect 125508 336796 125560 336802
rect 125508 336738 125560 336744
rect 121368 14340 121420 14346
rect 121368 14282 121420 14288
rect 119988 10192 120040 10198
rect 119988 10134 120040 10140
rect 118252 3318 118648 3346
rect 118252 480 118280 3318
rect 120000 2990 120028 10134
rect 121380 2990 121408 14282
rect 125416 14272 125468 14278
rect 125416 14214 125468 14220
rect 124128 10124 124180 10130
rect 124128 10066 124180 10072
rect 124140 3482 124168 10066
rect 125428 4214 125456 14214
rect 124220 4208 124272 4214
rect 124220 4150 124272 4156
rect 125416 4208 125468 4214
rect 125416 4150 125468 4156
rect 123036 3454 124168 3482
rect 119436 2984 119488 2990
rect 119436 2926 119488 2932
rect 119988 2984 120040 2990
rect 119988 2926 120040 2932
rect 120632 2984 120684 2990
rect 120632 2926 120684 2932
rect 121368 2984 121420 2990
rect 121368 2926 121420 2932
rect 119448 480 119476 2926
rect 120644 480 120672 2926
rect 121828 2848 121880 2854
rect 121828 2790 121880 2796
rect 121840 480 121868 2790
rect 123036 480 123064 3454
rect 124232 480 124260 4150
rect 125520 3482 125548 336738
rect 186228 13796 186280 13802
rect 186228 13738 186280 13744
rect 183468 13728 183520 13734
rect 183468 13670 183520 13676
rect 179328 13660 179380 13666
rect 179328 13602 179380 13608
rect 176568 13592 176620 13598
rect 176568 13534 176620 13540
rect 172428 13524 172480 13530
rect 172428 13466 172480 13472
rect 168288 13456 168340 13462
rect 168288 13398 168340 13404
rect 165528 13388 165580 13394
rect 165528 13330 165580 13336
rect 160008 13320 160060 13326
rect 160008 13262 160060 13268
rect 155868 12232 155920 12238
rect 155868 12174 155920 12180
rect 151728 12164 151780 12170
rect 151728 12106 151780 12112
rect 148968 12096 149020 12102
rect 148968 12038 149020 12044
rect 144828 12028 144880 12034
rect 144828 11970 144880 11976
rect 142068 11960 142120 11966
rect 142068 11902 142120 11908
rect 128268 11892 128320 11898
rect 128268 11834 128320 11840
rect 126888 11824 126940 11830
rect 126888 11766 126940 11772
rect 126900 3482 126928 11766
rect 128280 3482 128308 11834
rect 139676 9376 139728 9382
rect 139676 9318 139728 9324
rect 136088 9308 136140 9314
rect 136088 9250 136140 9256
rect 132590 8936 132646 8945
rect 132590 8871 132646 8880
rect 129002 7576 129058 7585
rect 129002 7511 129058 7520
rect 125428 3454 125548 3482
rect 126624 3454 126928 3482
rect 127820 3454 128308 3482
rect 125428 480 125456 3454
rect 126624 480 126652 3454
rect 127820 480 127848 3454
rect 129016 480 129044 7511
rect 131396 6656 131448 6662
rect 131396 6598 131448 6604
rect 130200 5364 130252 5370
rect 130200 5306 130252 5312
rect 130212 480 130240 5306
rect 131408 480 131436 6598
rect 132604 480 132632 8871
rect 134892 7540 134944 7546
rect 134892 7482 134944 7488
rect 133788 5432 133840 5438
rect 133788 5374 133840 5380
rect 133800 480 133828 5374
rect 134904 480 134932 7482
rect 136100 480 136128 9250
rect 138480 7472 138532 7478
rect 138480 7414 138532 7420
rect 137284 5500 137336 5506
rect 137284 5442 137336 5448
rect 137296 480 137324 5442
rect 138492 480 138520 7414
rect 139688 480 139716 9318
rect 141976 7404 142028 7410
rect 141976 7346 142028 7352
rect 140872 4208 140924 4214
rect 140872 4150 140924 4156
rect 140884 480 140912 4150
rect 141988 3482 142016 7346
rect 142080 4214 142108 11902
rect 143448 10056 143500 10062
rect 143448 9998 143500 10004
rect 142068 4208 142120 4214
rect 142068 4150 142120 4156
rect 143460 3482 143488 9998
rect 144840 3482 144868 11970
rect 147588 9988 147640 9994
rect 147588 9930 147640 9936
rect 145656 7336 145708 7342
rect 145656 7278 145708 7284
rect 141988 3454 142108 3482
rect 142080 480 142108 3454
rect 143276 3454 143488 3482
rect 144472 3454 144868 3482
rect 143276 480 143304 3454
rect 144472 480 144500 3454
rect 145668 480 145696 7278
rect 147600 3482 147628 9930
rect 148980 3482 149008 12038
rect 151636 9920 151688 9926
rect 151636 9862 151688 9868
rect 149244 7268 149296 7274
rect 149244 7210 149296 7216
rect 146864 3454 147628 3482
rect 148060 3454 149008 3482
rect 146864 480 146892 3454
rect 148060 480 148088 3454
rect 149256 480 149284 7210
rect 151648 4214 151676 9862
rect 150440 4208 150492 4214
rect 150440 4150 150492 4156
rect 151636 4208 151688 4214
rect 151636 4150 151688 4156
rect 150452 480 150480 4150
rect 151740 3482 151768 12106
rect 154488 9852 154540 9858
rect 154488 9794 154540 9800
rect 152740 7200 152792 7206
rect 152740 7142 152792 7148
rect 151556 3454 151768 3482
rect 151556 480 151584 3454
rect 152752 480 152780 7142
rect 154500 3482 154528 9794
rect 155880 3482 155908 12174
rect 158628 9784 158680 9790
rect 158628 9726 158680 9732
rect 156328 7132 156380 7138
rect 156328 7074 156380 7080
rect 153948 3454 154528 3482
rect 155144 3454 155908 3482
rect 153948 480 153976 3454
rect 155144 480 155172 3454
rect 156340 480 156368 7074
rect 158640 3482 158668 9726
rect 159916 7064 159968 7070
rect 159916 7006 159968 7012
rect 158720 4208 158772 4214
rect 158720 4150 158772 4156
rect 157536 3454 158668 3482
rect 157536 480 157564 3454
rect 158732 480 158760 4150
rect 159928 480 159956 7006
rect 160020 4214 160048 13262
rect 162768 12300 162820 12306
rect 162768 12242 162820 12248
rect 161388 9716 161440 9722
rect 161388 9658 161440 9664
rect 160008 4208 160060 4214
rect 160008 4150 160060 4156
rect 161400 3482 161428 9658
rect 161124 3454 161428 3482
rect 161124 480 161152 3454
rect 162780 626 162808 12242
rect 163504 6724 163556 6730
rect 163504 6666 163556 6672
rect 162320 598 162808 626
rect 162320 480 162348 598
rect 163516 480 163544 6666
rect 165540 610 165568 13330
rect 166908 12368 166960 12374
rect 166908 12310 166960 12316
rect 166920 610 166948 12310
rect 167092 6792 167144 6798
rect 167092 6734 167144 6740
rect 164700 604 164752 610
rect 164700 546 164752 552
rect 165528 604 165580 610
rect 165528 546 165580 552
rect 165896 604 165948 610
rect 165896 546 165948 552
rect 166908 604 166960 610
rect 166908 546 166960 552
rect 164712 480 164740 546
rect 165908 480 165936 546
rect 167104 480 167132 6734
rect 168300 626 168328 13398
rect 169668 12436 169720 12442
rect 169668 12378 169720 12384
rect 168208 598 168328 626
rect 169680 610 169708 12378
rect 170588 6860 170640 6866
rect 170588 6802 170640 6808
rect 169392 604 169444 610
rect 168208 480 168236 598
rect 169392 546 169444 552
rect 169668 604 169720 610
rect 169668 546 169720 552
rect 169404 480 169432 546
rect 170600 480 170628 6802
rect 172440 3346 172468 13466
rect 173808 11688 173860 11694
rect 173808 11630 173860 11636
rect 173820 3346 173848 11630
rect 176476 11620 176528 11626
rect 176476 11562 176528 11568
rect 174176 6112 174228 6118
rect 174176 6054 174228 6060
rect 171796 3318 172468 3346
rect 172992 3318 173848 3346
rect 171796 480 171824 3318
rect 172992 480 173020 3318
rect 174188 480 174216 6054
rect 175372 4208 175424 4214
rect 175372 4150 175424 4156
rect 175384 480 175412 4150
rect 176488 3482 176516 11562
rect 176580 4214 176608 13534
rect 177764 6044 177816 6050
rect 177764 5986 177816 5992
rect 176568 4208 176620 4214
rect 176568 4150 176620 4156
rect 176488 3454 176608 3482
rect 176580 480 176608 3454
rect 177776 480 177804 5986
rect 179340 3346 179368 13602
rect 180708 11552 180760 11558
rect 180708 11494 180760 11500
rect 180720 3346 180748 11494
rect 181352 5976 181404 5982
rect 181352 5918 181404 5924
rect 178972 3318 179368 3346
rect 180168 3318 180748 3346
rect 178972 480 179000 3318
rect 180168 480 180196 3318
rect 181364 480 181392 5918
rect 183480 610 183508 13670
rect 184848 11484 184900 11490
rect 184848 11426 184900 11432
rect 184860 6066 184888 11426
rect 184768 6038 184888 6066
rect 184768 610 184796 6038
rect 184848 5908 184900 5914
rect 184848 5850 184900 5856
rect 182548 604 182600 610
rect 182548 546 182600 552
rect 183468 604 183520 610
rect 183468 546 183520 552
rect 183744 604 183796 610
rect 183744 546 183796 552
rect 184756 604 184808 610
rect 184756 546 184808 552
rect 182560 480 182588 546
rect 183756 480 183784 546
rect 184860 480 184888 5850
rect 186240 626 186268 13738
rect 190368 13048 190420 13054
rect 190368 12990 190420 12996
rect 187608 11416 187660 11422
rect 187608 11358 187660 11364
rect 186056 598 186268 626
rect 187620 610 187648 11358
rect 188436 5840 188488 5846
rect 188436 5782 188488 5788
rect 187240 604 187292 610
rect 186056 480 186084 598
rect 187240 546 187292 552
rect 187608 604 187660 610
rect 187608 546 187660 552
rect 187252 480 187280 546
rect 188448 480 188476 5782
rect 190380 610 190408 12990
rect 206928 12980 206980 12986
rect 206928 12922 206980 12928
rect 191748 11348 191800 11354
rect 191748 11290 191800 11296
rect 191760 3346 191788 11290
rect 194508 11280 194560 11286
rect 194508 11222 194560 11228
rect 193220 9444 193272 9450
rect 193220 9386 193272 9392
rect 192024 5772 192076 5778
rect 192024 5714 192076 5720
rect 190840 3318 191788 3346
rect 189632 604 189684 610
rect 189632 546 189684 552
rect 190368 604 190420 610
rect 190368 546 190420 552
rect 189644 480 189672 546
rect 190840 480 190868 3318
rect 192036 480 192064 5714
rect 193232 480 193260 9386
rect 194520 3482 194548 11222
rect 198648 11212 198700 11218
rect 198648 11154 198700 11160
rect 196808 9512 196860 9518
rect 196808 9454 196860 9460
rect 195612 5704 195664 5710
rect 195612 5646 195664 5652
rect 194428 3454 194548 3482
rect 194428 480 194456 3454
rect 195624 480 195652 5646
rect 196820 480 196848 9454
rect 198660 3346 198688 11154
rect 203892 9648 203944 9654
rect 203892 9590 203944 9596
rect 200396 9580 200448 9586
rect 200396 9522 200448 9528
rect 199200 5636 199252 5642
rect 199200 5578 199252 5584
rect 198016 3318 198688 3346
rect 198016 480 198044 3318
rect 199212 480 199240 5578
rect 200408 480 200436 9522
rect 202696 5568 202748 5574
rect 202696 5510 202748 5516
rect 201500 4412 201552 4418
rect 201500 4354 201552 4360
rect 201512 480 201540 4354
rect 202708 480 202736 5510
rect 203904 480 203932 9590
rect 205088 4344 205140 4350
rect 205088 4286 205140 4292
rect 205100 480 205128 4286
rect 206940 3346 206968 12922
rect 211068 12912 211120 12918
rect 211068 12854 211120 12860
rect 207480 8900 207532 8906
rect 207480 8842 207532 8848
rect 206296 3318 206968 3346
rect 206296 480 206324 3318
rect 207492 480 207520 8842
rect 210976 8832 211028 8838
rect 210976 8774 211028 8780
rect 208674 4856 208730 4865
rect 208674 4791 208730 4800
rect 208688 480 208716 4791
rect 209872 4208 209924 4214
rect 209872 4150 209924 4156
rect 209884 480 209912 4150
rect 210988 3482 211016 8774
rect 211080 4214 211108 12854
rect 213828 12844 213880 12850
rect 213828 12786 213880 12792
rect 212264 4752 212316 4758
rect 212264 4694 212316 4700
rect 211068 4208 211120 4214
rect 211068 4150 211120 4156
rect 210988 3454 211108 3482
rect 211080 480 211108 3454
rect 212276 480 212304 4694
rect 213840 3346 213868 12786
rect 217968 12776 218020 12782
rect 217968 12718 218020 12724
rect 214656 8764 214708 8770
rect 214656 8706 214708 8712
rect 213472 3318 213868 3346
rect 213472 480 213500 3318
rect 214668 480 214696 8706
rect 215852 4684 215904 4690
rect 215852 4626 215904 4632
rect 215864 480 215892 4626
rect 217980 3346 218008 12718
rect 220728 12708 220780 12714
rect 220728 12650 220780 12656
rect 218152 8696 218204 8702
rect 218152 8638 218204 8644
rect 217060 3318 218008 3346
rect 217060 480 217088 3318
rect 218164 480 218192 8638
rect 219348 4616 219400 4622
rect 219348 4558 219400 4564
rect 219360 480 219388 4558
rect 220740 3346 220768 12650
rect 224868 12640 224920 12646
rect 224868 12582 224920 12588
rect 221740 8628 221792 8634
rect 221740 8570 221792 8576
rect 220556 3318 220768 3346
rect 220556 480 220584 3318
rect 221752 480 221780 8570
rect 222936 4548 222988 4554
rect 222936 4490 222988 4496
rect 222948 480 222976 4490
rect 224880 3346 224908 12582
rect 229008 12572 229060 12578
rect 229008 12514 229060 12520
rect 225328 8560 225380 8566
rect 225328 8502 225380 8508
rect 224144 3318 224908 3346
rect 224144 480 224172 3318
rect 225340 480 225368 8502
rect 228916 8492 228968 8498
rect 228916 8434 228968 8440
rect 227720 7608 227772 7614
rect 227720 7550 227772 7556
rect 226524 4480 226576 4486
rect 226524 4422 226576 4428
rect 226536 480 226564 4422
rect 227732 480 227760 7550
rect 228928 480 228956 8434
rect 229020 7614 229048 12514
rect 229008 7608 229060 7614
rect 229008 7550 229060 7556
rect 229112 4282 229140 340054
rect 229192 337272 229244 337278
rect 229190 337240 229192 337249
rect 229244 337240 229246 337249
rect 229190 337175 229246 337184
rect 230492 4894 230520 340068
rect 230584 340054 230966 340082
rect 230584 4962 230612 340054
rect 231044 337770 231072 340190
rect 230768 337742 231072 337770
rect 230768 321570 230796 337742
rect 231964 337385 231992 340068
rect 232056 340054 232438 340082
rect 231950 337376 232006 337385
rect 231950 337311 232006 337320
rect 230756 321564 230808 321570
rect 230756 321506 230808 321512
rect 230940 321564 230992 321570
rect 230940 321506 230992 321512
rect 230952 318782 230980 321506
rect 230940 318776 230992 318782
rect 230940 318718 230992 318724
rect 230848 309188 230900 309194
rect 230848 309130 230900 309136
rect 230860 205578 230888 309130
rect 230768 205550 230888 205578
rect 230768 202881 230796 205550
rect 230754 202872 230810 202881
rect 230754 202807 230810 202816
rect 231030 202872 231086 202881
rect 231030 202807 231086 202816
rect 231044 193254 231072 202807
rect 230848 193248 230900 193254
rect 230848 193190 230900 193196
rect 231032 193248 231084 193254
rect 231032 193190 231084 193196
rect 230860 186266 230888 193190
rect 230768 186238 230888 186266
rect 230768 183569 230796 186238
rect 230754 183560 230810 183569
rect 230754 183495 230810 183504
rect 231030 183560 231086 183569
rect 231030 183495 231086 183504
rect 231044 173942 231072 183495
rect 230848 173936 230900 173942
rect 230848 173878 230900 173884
rect 231032 173936 231084 173942
rect 231032 173878 231084 173884
rect 230860 166954 230888 173878
rect 230768 166926 230888 166954
rect 230768 157418 230796 166926
rect 230756 157412 230808 157418
rect 230756 157354 230808 157360
rect 230848 157344 230900 157350
rect 230848 157286 230900 157292
rect 230860 104854 230888 157286
rect 230848 104848 230900 104854
rect 230848 104790 230900 104796
rect 230848 95260 230900 95266
rect 230848 95202 230900 95208
rect 230860 61470 230888 95202
rect 230848 61464 230900 61470
rect 230848 61406 230900 61412
rect 230756 48340 230808 48346
rect 230756 48282 230808 48288
rect 230768 38758 230796 48282
rect 230756 38752 230808 38758
rect 230756 38694 230808 38700
rect 230756 37324 230808 37330
rect 230756 37266 230808 37272
rect 230768 12510 230796 37266
rect 230756 12504 230808 12510
rect 230756 12446 230808 12452
rect 230664 11144 230716 11150
rect 230664 11086 230716 11092
rect 230676 7682 230704 11086
rect 230664 7676 230716 7682
rect 230664 7618 230716 7624
rect 231308 7608 231360 7614
rect 231308 7550 231360 7556
rect 230572 4956 230624 4962
rect 230572 4898 230624 4904
rect 230480 4888 230532 4894
rect 230480 4830 230532 4836
rect 230112 4820 230164 4826
rect 230112 4762 230164 4768
rect 229100 4276 229152 4282
rect 229100 4218 229152 4224
rect 230124 480 230152 4762
rect 231320 480 231348 7550
rect 232056 3369 232084 340054
rect 232516 337770 232544 340190
rect 232240 337742 232544 337770
rect 232240 321570 232268 337742
rect 232228 321564 232280 321570
rect 232228 321506 232280 321512
rect 232412 321564 232464 321570
rect 232412 321506 232464 321512
rect 232424 313970 232452 321506
rect 232332 313942 232452 313970
rect 232332 205578 232360 313942
rect 232240 205550 232360 205578
rect 232240 202881 232268 205550
rect 232226 202872 232282 202881
rect 232226 202807 232282 202816
rect 232318 202736 232374 202745
rect 232318 202671 232374 202680
rect 232332 186266 232360 202671
rect 232240 186238 232360 186266
rect 232240 183569 232268 186238
rect 232226 183560 232282 183569
rect 232226 183495 232282 183504
rect 232318 183424 232374 183433
rect 232318 183359 232374 183368
rect 232332 182170 232360 183359
rect 232320 182164 232372 182170
rect 232320 182106 232372 182112
rect 232320 172576 232372 172582
rect 232240 172524 232320 172530
rect 232240 172518 232372 172524
rect 232240 172514 232360 172518
rect 232228 172508 232360 172514
rect 232280 172502 232360 172508
rect 232228 172450 232280 172456
rect 232240 172419 232268 172450
rect 232228 164212 232280 164218
rect 232228 164154 232280 164160
rect 232240 162874 232268 164154
rect 232240 162846 232360 162874
rect 232332 104802 232360 162846
rect 232240 104774 232360 104802
rect 232240 100094 232268 104774
rect 232228 100088 232280 100094
rect 232228 100030 232280 100036
rect 232320 87032 232372 87038
rect 232320 86974 232372 86980
rect 232332 85542 232360 86974
rect 232320 85536 232372 85542
rect 232320 85478 232372 85484
rect 232320 75948 232372 75954
rect 232320 75890 232372 75896
rect 232332 66230 232360 75890
rect 232320 66224 232372 66230
rect 232320 66166 232372 66172
rect 232320 56636 232372 56642
rect 232320 56578 232372 56584
rect 232332 53106 232360 56578
rect 232320 53100 232372 53106
rect 232320 53042 232372 53048
rect 232228 38752 232280 38758
rect 232228 38694 232280 38700
rect 232240 34218 232268 38694
rect 232240 34190 232360 34218
rect 232332 28966 232360 34190
rect 232228 28960 232280 28966
rect 232228 28902 232280 28908
rect 232320 28960 232372 28966
rect 232320 28902 232372 28908
rect 232240 12322 232268 28902
rect 232148 12294 232268 12322
rect 232148 5030 232176 12294
rect 232504 8424 232556 8430
rect 232504 8366 232556 8372
rect 232136 5024 232188 5030
rect 232136 4966 232188 4972
rect 232042 3360 232098 3369
rect 232042 3295 232098 3304
rect 232516 480 232544 8366
rect 233436 7002 233464 340068
rect 233528 340054 233910 340082
rect 233528 337414 233556 340054
rect 234356 337482 234384 340068
rect 234724 340054 234922 340082
rect 235092 340054 235382 340082
rect 235644 340054 235842 340082
rect 236394 340054 236500 340082
rect 234344 337476 234396 337482
rect 234344 337418 234396 337424
rect 233516 337408 233568 337414
rect 233516 337350 233568 337356
rect 233884 337408 233936 337414
rect 233884 337350 233936 337356
rect 233896 9110 233924 337350
rect 234620 337272 234672 337278
rect 234618 337240 234620 337249
rect 234672 337240 234674 337249
rect 234618 337175 234674 337184
rect 233884 9104 233936 9110
rect 233884 9046 233936 9052
rect 233424 6996 233476 7002
rect 233424 6938 233476 6944
rect 234724 5098 234752 340054
rect 235092 335594 235120 340054
rect 234816 335566 235120 335594
rect 234816 8974 234844 335566
rect 235644 335510 235672 340054
rect 236184 335708 236236 335714
rect 236184 335650 236236 335656
rect 236092 335640 236144 335646
rect 236092 335582 236144 335588
rect 235080 335504 235132 335510
rect 235080 335446 235132 335452
rect 235632 335504 235684 335510
rect 235632 335446 235684 335452
rect 235092 321638 235120 335446
rect 235080 321632 235132 321638
rect 235080 321574 235132 321580
rect 235080 321496 235132 321502
rect 235080 321438 235132 321444
rect 235092 313970 235120 321438
rect 234908 313942 235120 313970
rect 234908 302274 234936 313942
rect 234908 302246 235120 302274
rect 235092 299470 235120 302246
rect 235080 299464 235132 299470
rect 235080 299406 235132 299412
rect 235172 299464 235224 299470
rect 235172 299406 235224 299412
rect 235184 282826 235212 299406
rect 235092 282798 235212 282826
rect 235092 280158 235120 282798
rect 235080 280152 235132 280158
rect 235080 280094 235132 280100
rect 235172 280152 235224 280158
rect 235172 280094 235224 280100
rect 235184 263514 235212 280094
rect 235092 263486 235212 263514
rect 235092 260846 235120 263486
rect 235080 260840 235132 260846
rect 235080 260782 235132 260788
rect 235172 260840 235224 260846
rect 235172 260782 235224 260788
rect 235184 244202 235212 260782
rect 235092 244174 235212 244202
rect 235092 231878 235120 244174
rect 235080 231872 235132 231878
rect 235080 231814 235132 231820
rect 235172 231872 235224 231878
rect 235172 231814 235224 231820
rect 235184 224890 235212 231814
rect 235092 224862 235212 224890
rect 235092 212566 235120 224862
rect 235080 212560 235132 212566
rect 235080 212502 235132 212508
rect 235172 212560 235224 212566
rect 235172 212502 235224 212508
rect 235184 205578 235212 212502
rect 235092 205550 235212 205578
rect 235092 193254 235120 205550
rect 235080 193248 235132 193254
rect 235080 193190 235132 193196
rect 235172 193248 235224 193254
rect 235172 193190 235224 193196
rect 235184 186266 235212 193190
rect 235092 186238 235212 186266
rect 235092 173942 235120 186238
rect 235080 173936 235132 173942
rect 235080 173878 235132 173884
rect 235172 173936 235224 173942
rect 235172 173878 235224 173884
rect 235184 166954 235212 173878
rect 235092 166926 235212 166954
rect 235092 154578 235120 166926
rect 235092 154550 235212 154578
rect 235184 147642 235212 154550
rect 235092 147614 235212 147642
rect 235092 140026 235120 147614
rect 236000 144900 236052 144906
rect 236000 144842 236052 144848
rect 234908 139998 235120 140026
rect 234908 135289 234936 139998
rect 236012 135289 236040 144842
rect 234894 135280 234950 135289
rect 234894 135215 234950 135224
rect 235170 135280 235226 135289
rect 235170 135215 235226 135224
rect 235998 135280 236054 135289
rect 235998 135215 236054 135224
rect 235184 122806 235212 135215
rect 235172 122800 235224 122806
rect 235172 122742 235224 122748
rect 235080 113212 235132 113218
rect 235080 113154 235132 113160
rect 235092 101454 235120 113154
rect 235080 101448 235132 101454
rect 235080 101390 235132 101396
rect 235264 101448 235316 101454
rect 235264 101390 235316 101396
rect 235276 96665 235304 101390
rect 235078 96656 235134 96665
rect 235078 96591 235134 96600
rect 235262 96656 235318 96665
rect 235262 96591 235318 96600
rect 235092 86986 235120 96591
rect 235092 86958 235212 86986
rect 235000 80102 235028 80133
rect 235184 80102 235212 86958
rect 234988 80096 235040 80102
rect 235172 80096 235224 80102
rect 235040 80044 235120 80050
rect 234988 80038 235120 80044
rect 235172 80038 235224 80044
rect 235000 80022 235120 80038
rect 235092 60738 235120 80022
rect 235000 60710 235120 60738
rect 235000 60602 235028 60710
rect 235000 60574 235120 60602
rect 235092 41426 235120 60574
rect 235000 41398 235120 41426
rect 235000 41290 235028 41398
rect 235000 41262 235120 41290
rect 235092 19394 235120 41262
rect 235000 19366 235120 19394
rect 235000 12458 235028 19366
rect 235000 12430 235120 12458
rect 235092 12322 235120 12430
rect 234908 12294 235120 12322
rect 234804 8968 234856 8974
rect 234804 8910 234856 8916
rect 234804 7676 234856 7682
rect 234804 7618 234856 7624
rect 234712 5092 234764 5098
rect 234712 5034 234764 5040
rect 233700 4888 233752 4894
rect 233700 4830 233752 4836
rect 233712 480 233740 4830
rect 234816 480 234844 7618
rect 234908 3534 234936 12294
rect 236000 8968 236052 8974
rect 236000 8910 236052 8916
rect 234896 3528 234948 3534
rect 234896 3470 234948 3476
rect 236012 480 236040 8910
rect 236104 5166 236132 335582
rect 236196 9042 236224 335650
rect 236472 321586 236500 340054
rect 236564 340054 236854 340082
rect 237024 340054 237314 340082
rect 236564 335646 236592 340054
rect 237024 335714 237052 340054
rect 237852 337754 237880 340068
rect 237840 337748 237892 337754
rect 237840 337690 237892 337696
rect 238312 337482 238340 340068
rect 238786 340054 238892 340082
rect 238300 337476 238352 337482
rect 238300 337418 238352 337424
rect 237012 335708 237064 335714
rect 237012 335650 237064 335656
rect 236552 335640 236604 335646
rect 236552 335582 236604 335588
rect 236288 321558 236500 321586
rect 236288 318782 236316 321558
rect 236276 318776 236328 318782
rect 236276 318718 236328 318724
rect 236276 309256 236328 309262
rect 236276 309198 236328 309204
rect 236288 309126 236316 309198
rect 236276 309120 236328 309126
rect 236276 309062 236328 309068
rect 236276 299600 236328 299606
rect 236276 299542 236328 299548
rect 236288 299470 236316 299542
rect 236276 299464 236328 299470
rect 236276 299406 236328 299412
rect 236276 289876 236328 289882
rect 236276 289818 236328 289824
rect 236288 289746 236316 289818
rect 236276 289740 236328 289746
rect 236276 289682 236328 289688
rect 236276 280288 236328 280294
rect 236276 280230 236328 280236
rect 236288 280158 236316 280230
rect 236276 280152 236328 280158
rect 236276 280094 236328 280100
rect 236276 270564 236328 270570
rect 236276 270506 236328 270512
rect 236288 270434 236316 270506
rect 236276 270428 236328 270434
rect 236276 270370 236328 270376
rect 236276 260976 236328 260982
rect 236276 260918 236328 260924
rect 236288 260846 236316 260918
rect 236276 260840 236328 260846
rect 236276 260782 236328 260788
rect 236276 251252 236328 251258
rect 236276 251194 236328 251200
rect 236288 251161 236316 251194
rect 236274 251152 236330 251161
rect 236274 251087 236330 251096
rect 236458 251152 236514 251161
rect 236458 251087 236514 251096
rect 236472 241534 236500 251087
rect 236276 241528 236328 241534
rect 236276 241470 236328 241476
rect 236460 241528 236512 241534
rect 236460 241470 236512 241476
rect 236288 231849 236316 241470
rect 236274 231840 236330 231849
rect 236274 231775 236330 231784
rect 236458 231840 236514 231849
rect 236458 231775 236514 231784
rect 236472 222222 236500 231775
rect 236276 222216 236328 222222
rect 236276 222158 236328 222164
rect 236460 222216 236512 222222
rect 236460 222158 236512 222164
rect 236288 212537 236316 222158
rect 236274 212528 236330 212537
rect 236274 212463 236330 212472
rect 236458 212528 236514 212537
rect 236458 212463 236514 212472
rect 236472 202910 236500 212463
rect 236276 202904 236328 202910
rect 236276 202846 236328 202852
rect 236460 202904 236512 202910
rect 236460 202846 236512 202852
rect 236288 193225 236316 202846
rect 236274 193216 236330 193225
rect 236274 193151 236330 193160
rect 236458 193216 236514 193225
rect 236458 193151 236514 193160
rect 236472 183598 236500 193151
rect 236276 183592 236328 183598
rect 236274 183560 236276 183569
rect 236460 183592 236512 183598
rect 236328 183560 236330 183569
rect 236274 183495 236330 183504
rect 236458 183560 236460 183569
rect 236512 183560 236514 183569
rect 236458 183495 236514 183504
rect 236472 173942 236500 183495
rect 236368 173936 236420 173942
rect 236366 173904 236368 173913
rect 236460 173936 236512 173942
rect 236420 173904 236422 173913
rect 236460 173878 236512 173884
rect 236550 173904 236606 173913
rect 236366 173839 236422 173848
rect 236550 173839 236606 173848
rect 236564 164257 236592 173839
rect 236274 164248 236330 164257
rect 236274 164183 236330 164192
rect 236550 164248 236606 164257
rect 236550 164183 236606 164192
rect 236288 144906 236316 164183
rect 236276 144900 236328 144906
rect 236276 144842 236328 144848
rect 236274 135280 236330 135289
rect 236274 135215 236330 135224
rect 236288 96626 236316 135215
rect 236276 96620 236328 96626
rect 236276 96562 236328 96568
rect 236276 87032 236328 87038
rect 236276 86974 236328 86980
rect 236288 85542 236316 86974
rect 236276 85536 236328 85542
rect 236276 85478 236328 85484
rect 236276 75948 236328 75954
rect 236276 75890 236328 75896
rect 236288 67658 236316 75890
rect 236276 67652 236328 67658
rect 236276 67594 236328 67600
rect 236368 67584 236420 67590
rect 236368 67526 236420 67532
rect 236380 61470 236408 67526
rect 236368 61464 236420 61470
rect 236368 61406 236420 61412
rect 236276 48408 236328 48414
rect 236276 48350 236328 48356
rect 236288 46918 236316 48350
rect 236276 46912 236328 46918
rect 236276 46854 236328 46860
rect 236460 37324 236512 37330
rect 236460 37266 236512 37272
rect 236472 31634 236500 37266
rect 236380 31606 236500 31634
rect 236380 28966 236408 31606
rect 236368 28960 236420 28966
rect 236368 28902 236420 28908
rect 236368 19372 236420 19378
rect 236368 19314 236420 19320
rect 236380 12458 236408 19314
rect 236380 12430 236500 12458
rect 236472 12322 236500 12430
rect 236288 12294 236500 12322
rect 236184 9036 236236 9042
rect 236184 8978 236236 8984
rect 236092 5160 236144 5166
rect 236092 5102 236144 5108
rect 236288 3466 236316 12294
rect 238864 7750 238892 340054
rect 238956 340054 239338 340082
rect 239508 340054 239798 340082
rect 240258 340054 240364 340082
rect 238956 11762 238984 340054
rect 239508 331242 239536 340054
rect 239140 331214 239536 331242
rect 239140 321706 239168 331214
rect 239128 321700 239180 321706
rect 239128 321642 239180 321648
rect 239128 321564 239180 321570
rect 239128 321506 239180 321512
rect 239140 318866 239168 321506
rect 239140 318838 239260 318866
rect 239232 318782 239260 318838
rect 239220 318776 239272 318782
rect 239220 318718 239272 318724
rect 239220 309188 239272 309194
rect 239220 309130 239272 309136
rect 239232 292602 239260 309130
rect 239220 292596 239272 292602
rect 239220 292538 239272 292544
rect 239220 289876 239272 289882
rect 239220 289818 239272 289824
rect 239232 282826 239260 289818
rect 239140 282798 239260 282826
rect 239140 280158 239168 282798
rect 239128 280152 239180 280158
rect 239128 280094 239180 280100
rect 239220 270564 239272 270570
rect 239220 270506 239272 270512
rect 239232 263514 239260 270506
rect 239140 263486 239260 263514
rect 239140 260846 239168 263486
rect 239128 260840 239180 260846
rect 239128 260782 239180 260788
rect 239220 251252 239272 251258
rect 239220 251194 239272 251200
rect 239232 244202 239260 251194
rect 239140 244174 239260 244202
rect 239140 241482 239168 244174
rect 239140 241454 239260 241482
rect 239232 224890 239260 241454
rect 239140 224862 239260 224890
rect 239140 222170 239168 224862
rect 239140 222142 239260 222170
rect 239232 205578 239260 222142
rect 239140 205550 239260 205578
rect 239140 193254 239168 205550
rect 239128 193248 239180 193254
rect 239128 193190 239180 193196
rect 239220 193248 239272 193254
rect 239220 193190 239272 193196
rect 239232 186266 239260 193190
rect 239140 186238 239260 186266
rect 239140 173942 239168 186238
rect 239128 173936 239180 173942
rect 239128 173878 239180 173884
rect 239220 173936 239272 173942
rect 239220 173878 239272 173884
rect 239232 166954 239260 173878
rect 239140 166926 239260 166954
rect 239140 154578 239168 166926
rect 239140 154550 239260 154578
rect 239232 147642 239260 154550
rect 239140 147614 239260 147642
rect 239140 138038 239168 147614
rect 239128 138032 239180 138038
rect 239128 137974 239180 137980
rect 239220 137964 239272 137970
rect 239220 137906 239272 137912
rect 239232 122806 239260 137906
rect 239220 122800 239272 122806
rect 239220 122742 239272 122748
rect 239128 118040 239180 118046
rect 239128 117982 239180 117988
rect 239140 99414 239168 117982
rect 239128 99408 239180 99414
rect 239128 99350 239180 99356
rect 239128 99272 239180 99278
rect 239128 99214 239180 99220
rect 239140 70514 239168 99214
rect 239128 70508 239180 70514
rect 239128 70450 239180 70456
rect 239128 70372 239180 70378
rect 239128 70314 239180 70320
rect 239140 31822 239168 70314
rect 239128 31816 239180 31822
rect 239128 31758 239180 31764
rect 239036 31748 239088 31754
rect 239036 31690 239088 31696
rect 239048 19446 239076 31690
rect 239036 19440 239088 19446
rect 239036 19382 239088 19388
rect 239036 19304 239088 19310
rect 239036 19246 239088 19252
rect 238944 11756 238996 11762
rect 238944 11698 238996 11704
rect 238852 7744 238904 7750
rect 238852 7686 238904 7692
rect 238392 6996 238444 7002
rect 238392 6938 238444 6944
rect 237196 4956 237248 4962
rect 237196 4898 237248 4904
rect 236276 3460 236328 3466
rect 236276 3402 236328 3408
rect 237208 480 237236 4898
rect 238404 480 238432 6938
rect 239048 3670 239076 19246
rect 239588 9036 239640 9042
rect 239588 8978 239640 8984
rect 239036 3664 239088 3670
rect 239036 3606 239088 3612
rect 239600 480 239628 8978
rect 240336 3602 240364 340054
rect 240428 340054 240810 340082
rect 240428 7818 240456 340054
rect 241256 337414 241284 340068
rect 241716 337618 241744 340068
rect 241808 340054 242282 340082
rect 242360 340054 242742 340082
rect 243096 340054 243202 340082
rect 243464 340054 243754 340082
rect 241704 337612 241756 337618
rect 241704 337554 241756 337560
rect 241244 337408 241296 337414
rect 241244 337350 241296 337356
rect 241612 335640 241664 335646
rect 241612 335582 241664 335588
rect 241426 40352 241482 40361
rect 241426 40287 241428 40296
rect 241480 40287 241482 40296
rect 241428 40258 241480 40264
rect 241426 16824 241482 16833
rect 241426 16759 241482 16768
rect 241440 16697 241468 16759
rect 241426 16688 241482 16697
rect 241426 16623 241482 16632
rect 241624 13122 241652 335582
rect 241612 13116 241664 13122
rect 241612 13058 241664 13064
rect 241808 7886 241836 340054
rect 242360 335646 242388 340054
rect 242348 335640 242400 335646
rect 242348 335582 242400 335588
rect 242992 332104 243044 332110
rect 242992 332046 243044 332052
rect 243004 7954 243032 332046
rect 242992 7948 243044 7954
rect 242992 7890 243044 7896
rect 241796 7880 241848 7886
rect 241796 7822 241848 7828
rect 240416 7812 240468 7818
rect 240416 7754 240468 7760
rect 241980 7744 242032 7750
rect 241980 7686 242032 7692
rect 240784 5024 240836 5030
rect 240784 4966 240836 4972
rect 240324 3596 240376 3602
rect 240324 3538 240376 3544
rect 240796 480 240824 4966
rect 241992 480 242020 7686
rect 243096 3738 243124 340054
rect 243464 332110 243492 340054
rect 244200 337822 244228 340068
rect 244188 337816 244240 337822
rect 244188 337758 244240 337764
rect 244660 337686 244688 340068
rect 244648 337680 244700 337686
rect 244648 337622 244700 337628
rect 244752 335594 244780 340190
rect 245686 340054 245792 340082
rect 244476 335566 244780 335594
rect 243452 332104 243504 332110
rect 243452 332046 243504 332052
rect 244476 311846 244504 335566
rect 244464 311840 244516 311846
rect 244464 311782 244516 311788
rect 244464 309188 244516 309194
rect 244464 309130 244516 309136
rect 244476 292618 244504 309130
rect 244384 292590 244504 292618
rect 244384 292482 244412 292590
rect 244384 292454 244504 292482
rect 244476 289814 244504 292454
rect 244464 289808 244516 289814
rect 244464 289750 244516 289756
rect 244464 280220 244516 280226
rect 244464 280162 244516 280168
rect 244476 273306 244504 280162
rect 244384 273278 244504 273306
rect 244384 273170 244412 273278
rect 244384 273142 244504 273170
rect 244476 259457 244504 273142
rect 244462 259448 244518 259457
rect 244462 259383 244518 259392
rect 244646 259448 244702 259457
rect 244646 259383 244702 259392
rect 244660 254538 244688 259383
rect 244476 254510 244688 254538
rect 244476 241505 244504 254510
rect 244278 241496 244334 241505
rect 244278 241431 244334 241440
rect 244462 241496 244518 241505
rect 244462 241431 244518 241440
rect 244292 231878 244320 241431
rect 244280 231872 244332 231878
rect 244280 231814 244332 231820
rect 244464 231872 244516 231878
rect 244464 231814 244516 231820
rect 244476 222193 244504 231814
rect 244278 222184 244334 222193
rect 244278 222119 244334 222128
rect 244462 222184 244518 222193
rect 244462 222119 244518 222128
rect 244292 212566 244320 222119
rect 244280 212560 244332 212566
rect 244280 212502 244332 212508
rect 244464 212560 244516 212566
rect 244464 212502 244516 212508
rect 244476 202881 244504 212502
rect 244278 202872 244334 202881
rect 244278 202807 244334 202816
rect 244462 202872 244518 202881
rect 244462 202807 244518 202816
rect 244292 193254 244320 202807
rect 244280 193248 244332 193254
rect 244280 193190 244332 193196
rect 244464 193248 244516 193254
rect 244464 193190 244516 193196
rect 244476 176746 244504 193190
rect 244384 176718 244504 176746
rect 244384 176610 244412 176718
rect 244384 176582 244504 176610
rect 244476 164218 244504 176582
rect 244280 164212 244332 164218
rect 244280 164154 244332 164160
rect 244464 164212 244516 164218
rect 244464 164154 244516 164160
rect 244292 154601 244320 164154
rect 244278 154592 244334 154601
rect 244278 154527 244334 154536
rect 244462 154592 244518 154601
rect 244462 154527 244518 154536
rect 244476 144906 244504 154527
rect 244280 144900 244332 144906
rect 244280 144842 244332 144848
rect 244464 144900 244516 144906
rect 244464 144842 244516 144848
rect 244292 135289 244320 144842
rect 244278 135280 244334 135289
rect 244278 135215 244334 135224
rect 244462 135280 244518 135289
rect 244462 135215 244518 135224
rect 244476 120766 244504 135215
rect 244464 120760 244516 120766
rect 244464 120702 244516 120708
rect 244648 120760 244700 120766
rect 244648 120702 244700 120708
rect 244660 115977 244688 120702
rect 244462 115968 244518 115977
rect 244462 115903 244518 115912
rect 244646 115968 244702 115977
rect 244646 115903 244702 115912
rect 244476 106264 244504 115903
rect 244384 106236 244504 106264
rect 244384 99414 244412 106236
rect 244372 99408 244424 99414
rect 244372 99350 244424 99356
rect 244464 99340 244516 99346
rect 244464 99282 244516 99288
rect 244476 70514 244504 99282
rect 244464 70508 244516 70514
rect 244464 70450 244516 70456
rect 244464 66292 244516 66298
rect 244464 66234 244516 66240
rect 244476 53854 244504 66234
rect 244372 53848 244424 53854
rect 244372 53790 244424 53796
rect 244464 53848 244516 53854
rect 244464 53790 244516 53796
rect 244384 44169 244412 53790
rect 244370 44160 244426 44169
rect 244370 44095 244426 44104
rect 244554 44160 244610 44169
rect 244554 44095 244610 44104
rect 244568 34542 244596 44095
rect 245016 40316 245068 40322
rect 245016 40258 245068 40264
rect 245028 40089 245056 40258
rect 245014 40080 245070 40089
rect 245014 40015 245070 40024
rect 244372 34536 244424 34542
rect 244372 34478 244424 34484
rect 244556 34536 244608 34542
rect 244556 34478 244608 34484
rect 244384 31906 244412 34478
rect 244384 31878 244504 31906
rect 244476 24818 244504 31878
rect 244464 24812 244516 24818
rect 244464 24754 244516 24760
rect 243176 9104 243228 9110
rect 243176 9046 243228 9052
rect 243084 3732 243136 3738
rect 243084 3674 243136 3680
rect 243188 480 243216 9046
rect 244372 8356 244424 8362
rect 244372 8298 244424 8304
rect 244384 8022 244412 8298
rect 244372 8016 244424 8022
rect 244372 7958 244424 7964
rect 245568 7812 245620 7818
rect 245568 7754 245620 7760
rect 244372 5092 244424 5098
rect 244372 5034 244424 5040
rect 244384 480 244412 5034
rect 245580 480 245608 7754
rect 245764 3806 245792 340054
rect 245948 340054 246146 340082
rect 245844 335504 245896 335510
rect 245844 335446 245896 335452
rect 245856 8090 245884 335446
rect 245844 8084 245896 8090
rect 245844 8026 245896 8032
rect 245948 3874 245976 340054
rect 246684 335510 246712 340068
rect 247144 337890 247172 340068
rect 247604 337958 247632 340068
rect 247592 337952 247644 337958
rect 247592 337894 247644 337900
rect 247132 337884 247184 337890
rect 247132 337826 247184 337832
rect 247684 336524 247736 336530
rect 247684 336466 247736 336472
rect 246672 335504 246724 335510
rect 246672 335446 246724 335452
rect 247132 334212 247184 334218
rect 247132 334154 247184 334160
rect 247144 331106 247172 334154
rect 247144 331078 247264 331106
rect 247236 302274 247264 331078
rect 247144 302246 247264 302274
rect 247144 302138 247172 302246
rect 247144 302110 247264 302138
rect 247236 282962 247264 302110
rect 247144 282934 247264 282962
rect 247144 282826 247172 282934
rect 247144 282798 247264 282826
rect 247236 263650 247264 282798
rect 247144 263622 247264 263650
rect 247144 263514 247172 263622
rect 247144 263486 247264 263514
rect 247236 244338 247264 263486
rect 247144 244310 247264 244338
rect 247144 244202 247172 244310
rect 247144 244174 247264 244202
rect 247236 225026 247264 244174
rect 247144 224998 247264 225026
rect 247144 224890 247172 224998
rect 247144 224862 247264 224890
rect 247236 205714 247264 224862
rect 247144 205686 247264 205714
rect 247144 205578 247172 205686
rect 247144 205550 247264 205578
rect 247236 186402 247264 205550
rect 247144 186374 247264 186402
rect 247144 186266 247172 186374
rect 247144 186238 247264 186266
rect 247236 167090 247264 186238
rect 247144 167062 247264 167090
rect 247144 166954 247172 167062
rect 247144 166926 247264 166954
rect 247236 164200 247264 166926
rect 247236 164172 247356 164200
rect 247328 154630 247356 164172
rect 247224 154624 247276 154630
rect 247224 154566 247276 154572
rect 247316 154624 247368 154630
rect 247316 154566 247368 154572
rect 247236 147778 247264 154566
rect 247236 147750 247356 147778
rect 247328 144945 247356 147750
rect 247130 144936 247186 144945
rect 247314 144936 247370 144945
rect 247130 144871 247132 144880
rect 247184 144871 247186 144880
rect 247224 144900 247276 144906
rect 247132 144842 247184 144848
rect 247314 144871 247370 144880
rect 247224 144842 247276 144848
rect 247236 128466 247264 144842
rect 247144 128438 247264 128466
rect 247144 128330 247172 128438
rect 247144 128302 247264 128330
rect 247236 106264 247264 128302
rect 247144 106236 247264 106264
rect 247144 96801 247172 106236
rect 247130 96792 247186 96801
rect 247130 96727 247186 96736
rect 247130 96656 247186 96665
rect 247130 96591 247132 96600
rect 247184 96591 247186 96600
rect 247132 96562 247184 96568
rect 247132 89684 247184 89690
rect 247132 89626 247184 89632
rect 247144 86986 247172 89626
rect 247144 86958 247264 86986
rect 247236 80238 247264 86958
rect 247224 80232 247276 80238
rect 247224 80174 247276 80180
rect 247224 77308 247276 77314
rect 247224 77250 247276 77256
rect 247236 67590 247264 77250
rect 247132 67584 247184 67590
rect 247132 67526 247184 67532
rect 247224 67584 247276 67590
rect 247224 67526 247276 67532
rect 247144 58018 247172 67526
rect 247144 57990 247264 58018
rect 247236 47002 247264 57990
rect 247144 46974 247264 47002
rect 247144 46918 247172 46974
rect 247132 46912 247184 46918
rect 247132 46854 247184 46860
rect 247132 34536 247184 34542
rect 247132 34478 247184 34484
rect 247144 31226 247172 34478
rect 247052 31198 247172 31226
rect 247052 26382 247080 31198
rect 247040 26376 247092 26382
rect 247040 26318 247092 26324
rect 247132 26376 247184 26382
rect 247132 26318 247184 26324
rect 247144 24834 247172 26318
rect 247144 24806 247264 24834
rect 247236 22166 247264 24806
rect 247224 22160 247276 22166
rect 247224 22102 247276 22108
rect 247132 22092 247184 22098
rect 247132 22034 247184 22040
rect 247144 9178 247172 22034
rect 247132 9172 247184 9178
rect 247132 9114 247184 9120
rect 246764 8356 246816 8362
rect 246764 8298 246816 8304
rect 245936 3868 245988 3874
rect 245936 3810 245988 3816
rect 245752 3800 245804 3806
rect 245752 3742 245804 3748
rect 246776 480 246804 8298
rect 247696 3942 247724 336466
rect 248156 334218 248184 340068
rect 248512 337748 248564 337754
rect 248512 337690 248564 337696
rect 248144 334212 248196 334218
rect 248144 334154 248196 334160
rect 248420 29232 248472 29238
rect 248418 29200 248420 29209
rect 248472 29200 248474 29209
rect 248418 29135 248474 29144
rect 248524 5234 248552 337690
rect 248616 336530 248644 340068
rect 248708 340054 249090 340082
rect 248604 336524 248656 336530
rect 248604 336466 248656 336472
rect 248512 5228 248564 5234
rect 248512 5170 248564 5176
rect 247960 5160 248012 5166
rect 247960 5102 248012 5108
rect 247684 3936 247736 3942
rect 247684 3878 247736 3884
rect 247972 480 248000 5102
rect 248708 4010 248736 340054
rect 249536 337754 249564 340068
rect 249904 340054 250102 340082
rect 249524 337748 249576 337754
rect 249524 337690 249576 337696
rect 249246 336696 249302 336705
rect 249246 336631 249302 336640
rect 249064 336252 249116 336258
rect 249064 336194 249116 336200
rect 249076 4078 249104 336194
rect 249260 327185 249288 336631
rect 249246 327176 249302 327185
rect 249246 327111 249302 327120
rect 249246 321464 249302 321473
rect 249246 321399 249302 321408
rect 249260 317665 249288 321399
rect 249246 317656 249302 317665
rect 249246 317591 249302 317600
rect 249246 298072 249302 298081
rect 249246 298007 249302 298016
rect 249260 288561 249288 298007
rect 249246 288552 249302 288561
rect 249246 288487 249302 288496
rect 249246 288416 249302 288425
rect 249246 288351 249302 288360
rect 249260 279041 249288 288351
rect 249246 279032 249302 279041
rect 249246 278967 249302 278976
rect 249430 277400 249486 277409
rect 249430 277335 249486 277344
rect 249444 267889 249472 277335
rect 249430 267880 249486 267889
rect 249430 267815 249486 267824
rect 249246 212528 249302 212537
rect 249246 212463 249302 212472
rect 249260 205465 249288 212463
rect 249246 205456 249302 205465
rect 249246 205391 249302 205400
rect 249614 202872 249670 202881
rect 249614 202807 249670 202816
rect 249628 196625 249656 202807
rect 249614 196616 249670 196625
rect 249614 196551 249670 196560
rect 249246 191584 249302 191593
rect 249246 191519 249302 191528
rect 249260 182209 249288 191519
rect 249246 182200 249302 182209
rect 249246 182135 249302 182144
rect 249430 180568 249486 180577
rect 249430 180503 249486 180512
rect 249444 173913 249472 180503
rect 249430 173904 249486 173913
rect 249430 173839 249486 173848
rect 249800 80776 249852 80782
rect 249800 80718 249852 80724
rect 249812 75993 249840 80718
rect 249798 75984 249854 75993
rect 249798 75919 249854 75928
rect 249904 9246 249932 340054
rect 250444 337408 250496 337414
rect 250444 337350 250496 337356
rect 250168 328500 250220 328506
rect 250168 328442 250220 328448
rect 250180 314022 250208 328442
rect 250168 314016 250220 314022
rect 250168 313958 250220 313964
rect 250168 313880 250220 313886
rect 250168 313822 250220 313828
rect 250180 292618 250208 313822
rect 250088 292590 250208 292618
rect 250088 289814 250116 292590
rect 250076 289808 250128 289814
rect 250076 289750 250128 289756
rect 250352 289808 250404 289814
rect 250352 289750 250404 289756
rect 250364 288425 250392 289750
rect 250074 288416 250130 288425
rect 250074 288351 250130 288360
rect 250350 288416 250406 288425
rect 250350 288351 250406 288360
rect 250088 278798 250116 288351
rect 250076 278792 250128 278798
rect 250076 278734 250128 278740
rect 250168 278792 250220 278798
rect 250168 278734 250220 278740
rect 250180 273358 250208 278734
rect 250168 273352 250220 273358
rect 250168 273294 250220 273300
rect 250076 273216 250128 273222
rect 250076 273158 250128 273164
rect 250088 269074 250116 273158
rect 250076 269068 250128 269074
rect 250076 269010 250128 269016
rect 250168 259480 250220 259486
rect 250168 259422 250220 259428
rect 250180 259350 250208 259422
rect 250168 259344 250220 259350
rect 250168 259286 250220 259292
rect 250352 251116 250404 251122
rect 250352 251058 250404 251064
rect 250364 231878 250392 251058
rect 250076 231872 250128 231878
rect 250076 231814 250128 231820
rect 250352 231872 250404 231878
rect 250352 231814 250404 231820
rect 250088 227202 250116 231814
rect 250088 227174 250392 227202
rect 250364 212566 250392 227174
rect 250076 212560 250128 212566
rect 250076 212502 250128 212508
rect 250352 212560 250404 212566
rect 250352 212502 250404 212508
rect 250088 211138 250116 212502
rect 250076 211132 250128 211138
rect 250076 211074 250128 211080
rect 250260 211132 250312 211138
rect 250260 211074 250312 211080
rect 250272 201498 250300 211074
rect 250272 201482 250392 201498
rect 250076 201476 250128 201482
rect 250272 201476 250404 201482
rect 250272 201470 250352 201476
rect 250076 201418 250128 201424
rect 250352 201418 250404 201424
rect 250088 200122 250116 201418
rect 250076 200116 250128 200122
rect 250076 200058 250128 200064
rect 250076 186312 250128 186318
rect 250076 186254 250128 186260
rect 250088 177342 250116 186254
rect 250076 177336 250128 177342
rect 250076 177278 250128 177284
rect 250352 177336 250404 177342
rect 250352 177278 250404 177284
rect 250364 154737 250392 177278
rect 250350 154728 250406 154737
rect 250350 154663 250406 154672
rect 250074 154592 250130 154601
rect 250074 154527 250130 154536
rect 250088 149682 250116 154527
rect 249996 149654 250116 149682
rect 249996 144922 250024 149654
rect 249996 144894 250300 144922
rect 250272 143546 250300 144894
rect 250260 143540 250312 143546
rect 250260 143482 250312 143488
rect 250352 133952 250404 133958
rect 250352 133894 250404 133900
rect 250364 124137 250392 133894
rect 250166 124128 250222 124137
rect 250166 124063 250222 124072
rect 250350 124128 250406 124137
rect 250350 124063 250406 124072
rect 250180 96694 250208 124063
rect 250076 96688 250128 96694
rect 250076 96630 250128 96636
rect 250168 96688 250220 96694
rect 250168 96630 250220 96636
rect 250088 91882 250116 96630
rect 250088 91854 250208 91882
rect 250180 91610 250208 91854
rect 250088 91582 250208 91610
rect 250088 80782 250116 91582
rect 250076 80776 250128 80782
rect 250076 80718 250128 80724
rect 250074 75984 250130 75993
rect 250074 75919 250130 75928
rect 250088 75886 250116 75919
rect 250076 75880 250128 75886
rect 250076 75822 250128 75828
rect 250076 66292 250128 66298
rect 250076 66234 250128 66240
rect 250088 56794 250116 66234
rect 250088 56766 250208 56794
rect 250180 56658 250208 56766
rect 250088 56630 250208 56658
rect 250088 56574 250116 56630
rect 250076 56568 250128 56574
rect 250076 56510 250128 56516
rect 250076 51060 250128 51066
rect 250076 51002 250128 51008
rect 250088 47002 250116 51002
rect 250088 46974 250208 47002
rect 250180 46918 250208 46974
rect 250168 46912 250220 46918
rect 250168 46854 250220 46860
rect 250076 37324 250128 37330
rect 250076 37266 250128 37272
rect 250088 31770 250116 37266
rect 250088 31742 250300 31770
rect 250272 31634 250300 31742
rect 250180 31606 250300 31634
rect 250180 26246 250208 31606
rect 249984 26240 250036 26246
rect 249984 26182 250036 26188
rect 250168 26240 250220 26246
rect 250168 26182 250220 26188
rect 249892 9240 249944 9246
rect 249892 9182 249944 9188
rect 249156 7880 249208 7886
rect 249156 7822 249208 7828
rect 249064 4072 249116 4078
rect 249064 4014 249116 4020
rect 248696 4004 248748 4010
rect 248696 3946 248748 3952
rect 249168 480 249196 7822
rect 249996 6225 250024 26182
rect 250352 9172 250404 9178
rect 250352 9114 250404 9120
rect 249982 6216 250038 6225
rect 249982 6151 250038 6160
rect 250364 480 250392 9114
rect 250456 4146 250484 337350
rect 250548 336258 250576 340068
rect 250640 340054 251022 340082
rect 251284 340054 251574 340082
rect 250536 336252 250588 336258
rect 250536 336194 250588 336200
rect 250640 334490 250668 340054
rect 250628 334484 250680 334490
rect 250628 334426 250680 334432
rect 251178 87136 251234 87145
rect 251178 87071 251180 87080
rect 251232 87071 251234 87080
rect 251180 87042 251232 87048
rect 251086 16688 251142 16697
rect 251086 16623 251088 16632
rect 251140 16623 251142 16632
rect 251088 16594 251140 16600
rect 251284 10334 251312 340054
rect 252020 338026 252048 340068
rect 252008 338020 252060 338026
rect 252008 337962 252060 337968
rect 252480 337754 252508 340068
rect 252664 340054 253046 340082
rect 251456 337748 251508 337754
rect 251456 337690 251508 337696
rect 252468 337748 252520 337754
rect 252468 337690 252520 337696
rect 251468 321638 251496 337690
rect 251824 336728 251876 336734
rect 251824 336670 251876 336676
rect 251456 321632 251508 321638
rect 251456 321574 251508 321580
rect 251548 321428 251600 321434
rect 251548 321370 251600 321376
rect 251560 294710 251588 321370
rect 251548 294704 251600 294710
rect 251548 294646 251600 294652
rect 251456 289876 251508 289882
rect 251456 289818 251508 289824
rect 251468 280158 251496 289818
rect 251456 280152 251508 280158
rect 251456 280094 251508 280100
rect 251456 270564 251508 270570
rect 251456 270506 251508 270512
rect 251468 260846 251496 270506
rect 251456 260840 251508 260846
rect 251456 260782 251508 260788
rect 251456 251252 251508 251258
rect 251456 251194 251508 251200
rect 251468 241505 251496 251194
rect 251454 241496 251510 241505
rect 251454 241431 251510 241440
rect 251638 241496 251694 241505
rect 251638 241431 251694 241440
rect 251652 231878 251680 241431
rect 251456 231872 251508 231878
rect 251456 231814 251508 231820
rect 251640 231872 251692 231878
rect 251640 231814 251692 231820
rect 251468 222193 251496 231814
rect 251454 222184 251510 222193
rect 251454 222119 251510 222128
rect 251638 222184 251694 222193
rect 251638 222119 251694 222128
rect 251652 212566 251680 222119
rect 251456 212560 251508 212566
rect 251456 212502 251508 212508
rect 251640 212560 251692 212566
rect 251640 212502 251692 212508
rect 251468 202881 251496 212502
rect 251454 202872 251510 202881
rect 251454 202807 251510 202816
rect 251638 202872 251694 202881
rect 251638 202807 251694 202816
rect 251652 193254 251680 202807
rect 251456 193248 251508 193254
rect 251456 193190 251508 193196
rect 251640 193248 251692 193254
rect 251640 193190 251692 193196
rect 251468 183569 251496 193190
rect 251454 183560 251510 183569
rect 251454 183495 251510 183504
rect 251638 183560 251694 183569
rect 251638 183495 251694 183504
rect 251652 173942 251680 183495
rect 251456 173936 251508 173942
rect 251456 173878 251508 173884
rect 251640 173936 251692 173942
rect 251640 173878 251692 173884
rect 251468 164218 251496 173878
rect 251456 164212 251508 164218
rect 251456 164154 251508 164160
rect 251640 164212 251692 164218
rect 251640 164154 251692 164160
rect 251652 154601 251680 164154
rect 251454 154592 251510 154601
rect 251454 154527 251510 154536
rect 251638 154592 251694 154601
rect 251638 154527 251694 154536
rect 251468 138122 251496 154527
rect 251376 138094 251496 138122
rect 251376 137986 251404 138094
rect 251376 137958 251496 137986
rect 251468 125594 251496 137958
rect 251456 125588 251508 125594
rect 251456 125530 251508 125536
rect 251456 116000 251508 116006
rect 251456 115942 251508 115948
rect 251468 106282 251496 115942
rect 251456 106276 251508 106282
rect 251456 106218 251508 106224
rect 251456 96688 251508 96694
rect 251456 96630 251508 96636
rect 251468 86970 251496 96630
rect 251456 86964 251508 86970
rect 251456 86906 251508 86912
rect 251456 77308 251508 77314
rect 251456 77250 251508 77256
rect 251468 50946 251496 77250
rect 251376 50918 251496 50946
rect 251376 46918 251404 50918
rect 251364 46912 251416 46918
rect 251364 46854 251416 46860
rect 251456 37324 251508 37330
rect 251456 37266 251508 37272
rect 251468 35902 251496 37266
rect 251456 35896 251508 35902
rect 251456 35838 251508 35844
rect 251456 26308 251508 26314
rect 251456 26250 251508 26256
rect 251468 21457 251496 26250
rect 251454 21448 251510 21457
rect 251454 21383 251510 21392
rect 251272 10328 251324 10334
rect 251272 10270 251324 10276
rect 251362 8392 251418 8401
rect 251362 8327 251418 8336
rect 251376 6186 251404 8327
rect 251364 6180 251416 6186
rect 251364 6122 251416 6128
rect 251456 5228 251508 5234
rect 251456 5170 251508 5176
rect 250444 4140 250496 4146
rect 250444 4082 250496 4088
rect 251468 480 251496 5170
rect 251836 3398 251864 336670
rect 252664 10402 252692 340054
rect 253204 337544 253256 337550
rect 253204 337486 253256 337492
rect 252652 10396 252704 10402
rect 252652 10338 252704 10344
rect 252652 7948 252704 7954
rect 252652 7890 252704 7896
rect 251824 3392 251876 3398
rect 251824 3334 251876 3340
rect 252664 480 252692 7890
rect 253216 3330 253244 337486
rect 253492 337414 253520 340068
rect 253480 337408 253532 337414
rect 253480 337350 253532 337356
rect 253846 76120 253902 76129
rect 253846 76055 253848 76064
rect 253900 76055 253902 76064
rect 253848 76026 253900 76032
rect 253848 40112 253900 40118
rect 253846 40080 253848 40089
rect 253900 40080 253902 40089
rect 253846 40015 253902 40024
rect 253848 9240 253900 9246
rect 253848 9182 253900 9188
rect 253204 3324 253256 3330
rect 253204 3266 253256 3272
rect 253860 480 253888 9182
rect 253952 6254 253980 340068
rect 254044 340054 254518 340082
rect 254044 10470 254072 340054
rect 254964 338094 254992 340068
rect 255438 340054 255544 340082
rect 254952 338088 255004 338094
rect 254952 338030 255004 338036
rect 254584 337748 254636 337754
rect 254584 337690 254636 337696
rect 254032 10464 254084 10470
rect 254032 10406 254084 10412
rect 253940 6248 253992 6254
rect 253940 6190 253992 6196
rect 254596 3262 254624 337690
rect 255516 6322 255544 340054
rect 255608 340054 255990 340082
rect 255608 10538 255636 340054
rect 255964 337612 256016 337618
rect 255964 337554 256016 337560
rect 255596 10532 255648 10538
rect 255596 10474 255648 10480
rect 255504 6316 255556 6322
rect 255504 6258 255556 6264
rect 255044 3460 255096 3466
rect 255044 3402 255096 3408
rect 254584 3256 254636 3262
rect 254584 3198 254636 3204
rect 255056 480 255084 3402
rect 255976 3194 256004 337554
rect 256436 336734 256464 340068
rect 256804 340054 256910 340082
rect 256988 340054 257462 340082
rect 256424 336728 256476 336734
rect 256424 336670 256476 336676
rect 256240 8016 256292 8022
rect 256240 7958 256292 7964
rect 255964 3188 256016 3194
rect 255964 3130 256016 3136
rect 256252 480 256280 7958
rect 256804 6390 256832 340054
rect 256792 6384 256844 6390
rect 256792 6326 256844 6332
rect 256988 5302 257016 340054
rect 257344 337408 257396 337414
rect 257344 337350 257396 337356
rect 256976 5296 257028 5302
rect 256976 5238 257028 5244
rect 257356 3126 257384 337350
rect 257908 337278 257936 340068
rect 258276 340054 258382 340082
rect 258552 340054 258934 340082
rect 257896 337272 257948 337278
rect 257896 337214 257948 337220
rect 258172 334620 258224 334626
rect 258172 334562 258224 334568
rect 257894 29336 257950 29345
rect 257894 29271 257950 29280
rect 257908 29238 257936 29271
rect 257896 29232 257948 29238
rect 257896 29174 257948 29180
rect 258184 13190 258212 334562
rect 258172 13184 258224 13190
rect 258172 13126 258224 13132
rect 258276 6458 258304 340054
rect 258552 334626 258580 340054
rect 259380 337550 259408 340068
rect 259472 340054 259854 340082
rect 260116 340054 260406 340082
rect 259368 337544 259420 337550
rect 259368 337486 259420 337492
rect 258724 337476 258776 337482
rect 258724 337418 258776 337424
rect 258540 334620 258592 334626
rect 258540 334562 258592 334568
rect 258264 6452 258316 6458
rect 258264 6394 258316 6400
rect 257436 4004 257488 4010
rect 257436 3946 257488 3952
rect 257344 3120 257396 3126
rect 257344 3062 257396 3068
rect 257448 480 257476 3946
rect 258632 3528 258684 3534
rect 258632 3470 258684 3476
rect 258644 480 258672 3470
rect 258736 2990 258764 337418
rect 258816 337272 258868 337278
rect 258816 337214 258868 337220
rect 258828 3058 258856 337214
rect 259276 76084 259328 76090
rect 259276 76026 259328 76032
rect 259288 75970 259316 76026
rect 259366 75984 259422 75993
rect 259288 75942 259366 75970
rect 259366 75919 259422 75928
rect 259366 16688 259422 16697
rect 259366 16623 259368 16632
rect 259420 16623 259422 16632
rect 259368 16594 259420 16600
rect 259472 6526 259500 340054
rect 260116 337822 260144 340054
rect 259644 337816 259696 337822
rect 259644 337758 259696 337764
rect 260104 337816 260156 337822
rect 260104 337758 260156 337764
rect 259656 331226 259684 337758
rect 260104 337680 260156 337686
rect 260104 337622 260156 337628
rect 259644 331220 259696 331226
rect 259644 331162 259696 331168
rect 259828 331220 259880 331226
rect 259828 331162 259880 331168
rect 259840 328438 259868 331162
rect 259828 328432 259880 328438
rect 259828 328374 259880 328380
rect 259920 318844 259972 318850
rect 259920 318786 259972 318792
rect 259932 311914 259960 318786
rect 259736 311908 259788 311914
rect 259736 311850 259788 311856
rect 259920 311908 259972 311914
rect 259920 311850 259972 311856
rect 259748 309126 259776 311850
rect 259736 309120 259788 309126
rect 259736 309062 259788 309068
rect 259644 299600 259696 299606
rect 259644 299542 259696 299548
rect 259656 299470 259684 299542
rect 259644 299464 259696 299470
rect 259644 299406 259696 299412
rect 259828 299464 259880 299470
rect 259828 299406 259880 299412
rect 259840 289898 259868 299406
rect 259748 289870 259868 289898
rect 259748 289814 259776 289870
rect 259736 289808 259788 289814
rect 259736 289750 259788 289756
rect 259920 289808 259972 289814
rect 259920 289750 259972 289756
rect 259932 280265 259960 289750
rect 259550 280256 259606 280265
rect 259550 280191 259606 280200
rect 259918 280256 259974 280265
rect 259918 280191 259974 280200
rect 259564 280158 259592 280191
rect 259552 280152 259604 280158
rect 259552 280094 259604 280100
rect 259552 273080 259604 273086
rect 259552 273022 259604 273028
rect 259564 260846 259592 273022
rect 259552 260840 259604 260846
rect 259552 260782 259604 260788
rect 259552 253768 259604 253774
rect 259552 253710 259604 253716
rect 259564 251190 259592 253710
rect 259552 251184 259604 251190
rect 259552 251126 259604 251132
rect 259644 244180 259696 244186
rect 259644 244122 259696 244128
rect 259656 241398 259684 244122
rect 259644 241392 259696 241398
rect 259644 241334 259696 241340
rect 259828 241392 259880 241398
rect 259828 241334 259880 241340
rect 259840 222222 259868 241334
rect 259644 222216 259696 222222
rect 259644 222158 259696 222164
rect 259828 222216 259880 222222
rect 259828 222158 259880 222164
rect 259656 222086 259684 222158
rect 259644 222080 259696 222086
rect 259644 222022 259696 222028
rect 259828 222080 259880 222086
rect 259828 222022 259880 222028
rect 259840 215234 259868 222022
rect 259748 215206 259868 215234
rect 259748 205578 259776 215206
rect 259656 205550 259776 205578
rect 259656 202881 259684 205550
rect 259642 202872 259698 202881
rect 259642 202807 259698 202816
rect 259918 202872 259974 202881
rect 259918 202807 259974 202816
rect 259932 193254 259960 202807
rect 259736 193248 259788 193254
rect 259736 193190 259788 193196
rect 259920 193248 259972 193254
rect 259920 193190 259972 193196
rect 259748 186266 259776 193190
rect 259656 186238 259776 186266
rect 259656 179586 259684 186238
rect 259644 179580 259696 179586
rect 259644 179522 259696 179528
rect 259736 174004 259788 174010
rect 259736 173946 259788 173952
rect 259748 169114 259776 173946
rect 259736 169108 259788 169114
rect 259736 169050 259788 169056
rect 259920 169108 259972 169114
rect 259920 169050 259972 169056
rect 259932 164257 259960 169050
rect 259642 164248 259698 164257
rect 259918 164248 259974 164257
rect 259642 164183 259644 164192
rect 259696 164183 259698 164192
rect 259828 164212 259880 164218
rect 259644 164154 259696 164160
rect 259918 164183 259974 164192
rect 259828 164154 259880 164160
rect 259840 154222 259868 164154
rect 259828 154216 259880 154222
rect 259828 154158 259880 154164
rect 259644 145036 259696 145042
rect 259644 144978 259696 144984
rect 259656 137850 259684 144978
rect 259656 137822 259776 137850
rect 259748 128382 259776 137822
rect 259736 128376 259788 128382
rect 259736 128318 259788 128324
rect 259828 128308 259880 128314
rect 259828 128250 259880 128256
rect 259840 125526 259868 128250
rect 259736 125520 259788 125526
rect 259736 125462 259788 125468
rect 259828 125520 259880 125526
rect 259828 125462 259880 125468
rect 259748 116113 259776 125462
rect 259734 116104 259790 116113
rect 259734 116039 259790 116048
rect 259642 115968 259698 115977
rect 259642 115903 259698 115912
rect 259656 109018 259684 115903
rect 259656 108990 259868 109018
rect 259840 106282 259868 108990
rect 259552 106276 259604 106282
rect 259552 106218 259604 106224
rect 259828 106276 259880 106282
rect 259828 106218 259880 106224
rect 259564 96665 259592 106218
rect 259550 96656 259606 96665
rect 259550 96591 259606 96600
rect 259734 96656 259790 96665
rect 259734 96591 259790 96600
rect 259748 91746 259776 96591
rect 259748 91718 259868 91746
rect 259840 86986 259868 91718
rect 259840 86958 259960 86986
rect 259932 77738 259960 86958
rect 259748 77710 259960 77738
rect 259748 66298 259776 77710
rect 259644 66292 259696 66298
rect 259644 66234 259696 66240
rect 259736 66292 259788 66298
rect 259736 66234 259788 66240
rect 259656 56642 259684 66234
rect 259644 56636 259696 56642
rect 259644 56578 259696 56584
rect 259552 56568 259604 56574
rect 259552 56510 259604 56516
rect 259564 47002 259592 56510
rect 259564 46974 259684 47002
rect 259656 37210 259684 46974
rect 259656 37182 259868 37210
rect 259840 27674 259868 37182
rect 259736 27668 259788 27674
rect 259736 27610 259788 27616
rect 259828 27668 259880 27674
rect 259828 27610 259880 27616
rect 259748 22114 259776 27610
rect 259656 22086 259776 22114
rect 259656 13258 259684 22086
rect 259644 13252 259696 13258
rect 259644 13194 259696 13200
rect 259828 8084 259880 8090
rect 259828 8026 259880 8032
rect 259460 6520 259512 6526
rect 259460 6462 259512 6468
rect 258816 3052 258868 3058
rect 258816 2994 258868 3000
rect 258724 2984 258776 2990
rect 258724 2926 258776 2932
rect 259840 480 259868 8026
rect 260116 2922 260144 337622
rect 260852 337346 260880 340068
rect 261036 340054 261326 340082
rect 261496 340054 261878 340082
rect 260840 337340 260892 337346
rect 260840 337282 260892 337288
rect 260932 335640 260984 335646
rect 260932 335582 260984 335588
rect 260654 87136 260710 87145
rect 260654 87071 260656 87080
rect 260708 87071 260710 87080
rect 260656 87042 260708 87048
rect 260944 14482 260972 335582
rect 260932 14476 260984 14482
rect 260932 14418 260984 14424
rect 261036 6594 261064 340054
rect 261392 337612 261444 337618
rect 261392 337554 261444 337560
rect 261404 334370 261432 337554
rect 261496 335646 261524 340054
rect 262324 337754 262352 340068
rect 262416 340054 262798 340082
rect 263060 340054 263350 340082
rect 262312 337748 262364 337754
rect 262312 337690 262364 337696
rect 261484 335640 261536 335646
rect 261484 335582 261536 335588
rect 261404 334342 261524 334370
rect 261024 6588 261076 6594
rect 261024 6530 261076 6536
rect 260104 2916 260156 2922
rect 260104 2858 260156 2864
rect 261496 2854 261524 334342
rect 262416 8158 262444 340054
rect 263060 333062 263088 340054
rect 263796 337210 263824 340068
rect 263888 340054 264270 340082
rect 264440 340054 264822 340082
rect 263784 337204 263836 337210
rect 263784 337146 263836 337152
rect 263692 335640 263744 335646
rect 263692 335582 263744 335588
rect 262588 333056 262640 333062
rect 262588 332998 262640 333004
rect 263048 333056 263100 333062
rect 263048 332998 263100 333004
rect 262600 331226 262628 332998
rect 262588 331220 262640 331226
rect 262588 331162 262640 331168
rect 262772 331220 262824 331226
rect 262772 331162 262824 331168
rect 262784 317506 262812 331162
rect 262692 317478 262812 317506
rect 262692 315994 262720 317478
rect 262680 315988 262732 315994
rect 262680 315930 262732 315936
rect 262588 298240 262640 298246
rect 262588 298182 262640 298188
rect 262600 298110 262628 298182
rect 262588 298104 262640 298110
rect 262588 298046 262640 298052
rect 262588 297968 262640 297974
rect 262588 297910 262640 297916
rect 262600 280106 262628 297910
rect 262508 280078 262628 280106
rect 262508 270570 262536 280078
rect 262496 270564 262548 270570
rect 262496 270506 262548 270512
rect 262680 270564 262732 270570
rect 262680 270506 262732 270512
rect 262692 269090 262720 270506
rect 262600 269062 262720 269090
rect 262600 260914 262628 269062
rect 262588 260908 262640 260914
rect 262588 260850 262640 260856
rect 262600 259486 262628 259517
rect 262588 259480 262640 259486
rect 262640 259428 262720 259434
rect 262588 259422 262720 259428
rect 262600 259406 262720 259422
rect 262692 241602 262720 259406
rect 262680 241596 262732 241602
rect 262680 241538 262732 241544
rect 262588 241528 262640 241534
rect 262588 241470 262640 241476
rect 262600 235362 262628 241470
rect 262600 235334 262812 235362
rect 262784 222222 262812 235334
rect 262680 222216 262732 222222
rect 262680 222158 262732 222164
rect 262772 222216 262824 222222
rect 262772 222158 262824 222164
rect 262692 212514 262720 222158
rect 262692 212486 262812 212514
rect 262784 207942 262812 212486
rect 262588 207936 262640 207942
rect 262588 207878 262640 207884
rect 262772 207936 262824 207942
rect 262772 207878 262824 207884
rect 262600 202881 262628 207878
rect 262586 202872 262642 202881
rect 262586 202807 262642 202816
rect 262678 202736 262734 202745
rect 262678 202671 262734 202680
rect 262692 186266 262720 202671
rect 262600 186238 262720 186266
rect 262600 183569 262628 186238
rect 262586 183560 262642 183569
rect 262586 183495 262642 183504
rect 262770 183560 262826 183569
rect 262770 183495 262826 183504
rect 262784 178922 262812 183495
rect 262692 178894 262812 178922
rect 262692 161498 262720 178894
rect 262588 161492 262640 161498
rect 262588 161434 262640 161440
rect 262680 161492 262732 161498
rect 262680 161434 262732 161440
rect 262600 143546 262628 161434
rect 262588 143540 262640 143546
rect 262588 143482 262640 143488
rect 262864 143540 262916 143546
rect 262864 143482 262916 143488
rect 262876 120714 262904 143482
rect 262600 120686 262904 120714
rect 262600 109018 262628 120686
rect 262600 108990 262812 109018
rect 262784 101402 262812 108990
rect 262600 101374 262812 101402
rect 262600 98410 262628 101374
rect 262600 98382 262720 98410
rect 262692 60382 262720 98382
rect 262680 60376 262732 60382
rect 262680 60318 262732 60324
rect 262772 55276 262824 55282
rect 262772 55218 262824 55224
rect 262784 47054 262812 55218
rect 262772 47048 262824 47054
rect 262772 46990 262824 46996
rect 262680 46912 262732 46918
rect 262680 46854 262732 46860
rect 262692 35850 262720 46854
rect 262864 40112 262916 40118
rect 262862 40080 262864 40089
rect 262916 40080 262918 40089
rect 262862 40015 262918 40024
rect 262600 35822 262720 35850
rect 262600 26330 262628 35822
rect 262862 29336 262918 29345
rect 262862 29271 262918 29280
rect 262876 29073 262904 29271
rect 262862 29064 262918 29073
rect 262862 28999 262918 29008
rect 262600 26302 262720 26330
rect 262692 22114 262720 26302
rect 262600 22086 262720 22114
rect 262600 14550 262628 22086
rect 263704 14618 263732 335582
rect 263692 14612 263744 14618
rect 263692 14554 263744 14560
rect 262588 14544 262640 14550
rect 262588 14486 262640 14492
rect 263888 8226 263916 340054
rect 264440 335646 264468 340054
rect 265268 337074 265296 340068
rect 265452 340054 265742 340082
rect 265912 340054 266294 340082
rect 265256 337068 265308 337074
rect 265256 337010 265308 337016
rect 264428 335640 264480 335646
rect 264428 335582 264480 335588
rect 265072 335640 265124 335646
rect 265452 335594 265480 340054
rect 265912 335646 265940 340054
rect 266740 337414 266768 340068
rect 266924 340054 267214 340082
rect 267384 340054 267674 340082
rect 266728 337408 266780 337414
rect 266728 337350 266780 337356
rect 265072 335582 265124 335588
rect 264980 258052 265032 258058
rect 264980 257994 265032 258000
rect 264992 248441 265020 257994
rect 264978 248432 265034 248441
rect 264978 248367 265034 248376
rect 264980 190460 265032 190466
rect 264980 190402 265032 190408
rect 264992 180849 265020 190402
rect 264978 180840 265034 180849
rect 264978 180775 265034 180784
rect 264980 153128 265032 153134
rect 264980 153070 265032 153076
rect 264992 151774 265020 153070
rect 264980 151768 265032 151774
rect 264980 151710 265032 151716
rect 265084 143614 265112 335582
rect 265268 335566 265480 335594
rect 265900 335640 265952 335646
rect 265900 335582 265952 335588
rect 266452 335640 266504 335646
rect 266924 335594 266952 340054
rect 267384 335646 267412 340054
rect 268212 336938 268240 340068
rect 268396 340054 268686 340082
rect 269146 340054 269252 340082
rect 268200 336932 268252 336938
rect 268200 336874 268252 336880
rect 266452 335582 266504 335588
rect 265268 280226 265296 335566
rect 265256 280220 265308 280226
rect 265256 280162 265308 280168
rect 265256 280084 265308 280090
rect 265256 280026 265308 280032
rect 265268 277409 265296 280026
rect 265254 277400 265310 277409
rect 265254 277335 265310 277344
rect 265438 277400 265494 277409
rect 265438 277335 265494 277344
rect 265452 267782 265480 277335
rect 265256 267776 265308 267782
rect 265256 267718 265308 267724
rect 265440 267776 265492 267782
rect 265440 267718 265492 267724
rect 265268 264330 265296 267718
rect 265176 264302 265296 264330
rect 265176 259457 265204 264302
rect 265162 259448 265218 259457
rect 265162 259383 265218 259392
rect 265346 259448 265402 259457
rect 265346 259383 265402 259392
rect 265360 258058 265388 259383
rect 265348 258052 265400 258058
rect 265348 257994 265400 258000
rect 265162 248432 265218 248441
rect 265162 248367 265218 248376
rect 265176 234666 265204 248367
rect 265164 234660 265216 234666
rect 265164 234602 265216 234608
rect 265256 234524 265308 234530
rect 265256 234466 265308 234472
rect 265268 227202 265296 234466
rect 265268 227174 265388 227202
rect 265360 222222 265388 227174
rect 265164 222216 265216 222222
rect 265164 222158 265216 222164
rect 265348 222216 265400 222222
rect 265348 222158 265400 222164
rect 265176 212566 265204 222158
rect 265164 212560 265216 212566
rect 265256 212560 265308 212566
rect 265216 212508 265256 212514
rect 265164 212502 265308 212508
rect 265176 212486 265296 212502
rect 265176 202881 265204 212486
rect 265162 202872 265218 202881
rect 265162 202807 265218 202816
rect 265346 202872 265402 202881
rect 265346 202807 265402 202816
rect 265360 193254 265388 202807
rect 265256 193248 265308 193254
rect 265256 193190 265308 193196
rect 265348 193248 265400 193254
rect 265348 193190 265400 193196
rect 265268 190466 265296 193190
rect 265256 190460 265308 190466
rect 265256 190402 265308 190408
rect 265162 180840 265218 180849
rect 265162 180775 265164 180784
rect 265216 180775 265218 180784
rect 265256 180804 265308 180810
rect 265164 180746 265216 180752
rect 265256 180746 265308 180752
rect 265268 179382 265296 180746
rect 265256 179376 265308 179382
rect 265256 179318 265308 179324
rect 265348 161492 265400 161498
rect 265348 161434 265400 161440
rect 265360 153134 265388 161434
rect 265348 153128 265400 153134
rect 265348 153070 265400 153076
rect 265072 143608 265124 143614
rect 265072 143550 265124 143556
rect 265072 143472 265124 143478
rect 265072 143414 265124 143420
rect 265084 14686 265112 143414
rect 265256 142180 265308 142186
rect 265256 142122 265308 142128
rect 265268 142066 265296 142122
rect 265268 142038 265388 142066
rect 265360 133770 265388 142038
rect 265268 133742 265388 133770
rect 265268 130506 265296 133742
rect 265268 130478 265388 130506
rect 265360 125633 265388 130478
rect 265162 125624 265218 125633
rect 265162 125559 265164 125568
rect 265216 125559 265218 125568
rect 265346 125624 265402 125633
rect 265346 125559 265348 125568
rect 265164 125530 265216 125536
rect 265400 125559 265402 125568
rect 265348 125530 265400 125536
rect 265360 118538 265388 125530
rect 265268 118510 265388 118538
rect 265268 106350 265296 118510
rect 265164 106344 265216 106350
rect 265164 106286 265216 106292
rect 265256 106344 265308 106350
rect 265256 106286 265308 106292
rect 265176 104854 265204 106286
rect 265164 104848 265216 104854
rect 265164 104790 265216 104796
rect 265164 96620 265216 96626
rect 265164 96562 265216 96568
rect 265176 96393 265204 96562
rect 265162 96384 265218 96393
rect 265162 96319 265218 96328
rect 265254 89040 265310 89049
rect 265254 88975 265310 88984
rect 265268 82822 265296 88975
rect 265256 82816 265308 82822
rect 265256 82758 265308 82764
rect 265256 73228 265308 73234
rect 265256 73170 265308 73176
rect 265268 69578 265296 73170
rect 265268 69550 265480 69578
rect 265452 65906 265480 69550
rect 265360 65878 265480 65906
rect 265360 63510 265388 65878
rect 265348 63504 265400 63510
rect 265348 63446 265400 63452
rect 265256 53848 265308 53854
rect 265256 53790 265308 53796
rect 265268 50674 265296 53790
rect 265176 50646 265296 50674
rect 265176 50402 265204 50646
rect 265176 50374 265296 50402
rect 265268 41478 265296 50374
rect 265256 41472 265308 41478
rect 265256 41414 265308 41420
rect 265256 35964 265308 35970
rect 265256 35906 265308 35912
rect 265268 27606 265296 35906
rect 265256 27600 265308 27606
rect 265256 27542 265308 27548
rect 265164 18012 265216 18018
rect 265164 17954 265216 17960
rect 265072 14680 265124 14686
rect 265072 14622 265124 14628
rect 265176 8294 265204 17954
rect 266464 14754 266492 335582
rect 266740 335566 266952 335594
rect 267372 335640 267424 335646
rect 268396 335594 268424 340054
rect 269028 337408 269080 337414
rect 269028 337350 269080 337356
rect 267372 335582 267424 335588
rect 267844 335566 268424 335594
rect 266740 321722 266768 335566
rect 266740 321694 266860 321722
rect 266832 321450 266860 321694
rect 266740 321422 266860 321450
rect 266740 298110 266768 321422
rect 267844 321314 267872 335566
rect 267752 321286 267872 321314
rect 267752 309194 267780 321286
rect 267740 309188 267792 309194
rect 267740 309130 267792 309136
rect 267832 309188 267884 309194
rect 267832 309130 267884 309136
rect 267844 299606 267872 309130
rect 267832 299600 267884 299606
rect 267832 299542 267884 299548
rect 267740 299464 267792 299470
rect 267740 299406 267792 299412
rect 267752 298110 267780 299406
rect 266728 298104 266780 298110
rect 266728 298046 266780 298052
rect 267740 298104 267792 298110
rect 267740 298046 267792 298052
rect 266728 288448 266780 288454
rect 266728 288390 266780 288396
rect 267740 288448 267792 288454
rect 267740 288390 267792 288396
rect 266740 280140 266768 288390
rect 266740 280112 266860 280140
rect 266832 270609 266860 280112
rect 266818 270600 266874 270609
rect 267752 270570 267780 288390
rect 266818 270535 266874 270544
rect 267740 270564 267792 270570
rect 267740 270506 267792 270512
rect 267832 270564 267884 270570
rect 267832 270506 267884 270512
rect 266634 270464 266690 270473
rect 266634 270399 266690 270408
rect 266648 260914 266676 270399
rect 266636 260908 266688 260914
rect 266636 260850 266688 260856
rect 266728 260908 266780 260914
rect 266728 260850 266780 260856
rect 266740 254674 266768 260850
rect 267844 259486 267872 270506
rect 267740 259480 267792 259486
rect 267738 259448 267740 259457
rect 267832 259480 267884 259486
rect 267792 259448 267794 259457
rect 267832 259422 267884 259428
rect 267922 259448 267978 259457
rect 267738 259383 267794 259392
rect 267922 259383 267978 259392
rect 267936 258058 267964 259383
rect 267924 258052 267976 258058
rect 267924 257994 267976 258000
rect 268108 258052 268160 258058
rect 268108 257994 268160 258000
rect 266556 254646 266768 254674
rect 266556 253858 266584 254646
rect 266556 253830 266676 253858
rect 266648 241534 266676 253830
rect 268120 248441 268148 257994
rect 267738 248432 267794 248441
rect 267738 248367 267794 248376
rect 268106 248432 268162 248441
rect 268106 248367 268162 248376
rect 266636 241528 266688 241534
rect 266636 241470 266688 241476
rect 266728 241528 266780 241534
rect 266728 241470 266780 241476
rect 266740 234870 266768 241470
rect 267752 240106 267780 248367
rect 267740 240100 267792 240106
rect 267740 240042 267792 240048
rect 266728 234864 266780 234870
rect 266728 234806 266780 234812
rect 267924 231804 267976 231810
rect 267924 231746 267976 231752
rect 266728 230512 266780 230518
rect 266728 230454 266780 230460
rect 266740 217410 266768 230454
rect 266740 217382 266860 217410
rect 266832 212566 266860 217382
rect 267936 212566 267964 231746
rect 266636 212560 266688 212566
rect 266636 212502 266688 212508
rect 266820 212560 266872 212566
rect 266820 212502 266872 212508
rect 267832 212560 267884 212566
rect 267832 212502 267884 212508
rect 267924 212560 267976 212566
rect 267924 212502 267976 212508
rect 266648 205698 266676 212502
rect 267844 211138 267872 212502
rect 267832 211132 267884 211138
rect 267832 211074 267884 211080
rect 267924 211132 267976 211138
rect 267924 211074 267976 211080
rect 266636 205692 266688 205698
rect 266636 205634 266688 205640
rect 266728 205624 266780 205630
rect 266728 205566 266780 205572
rect 266740 198150 266768 205566
rect 266728 198144 266780 198150
rect 266728 198086 266780 198092
rect 266636 198076 266688 198082
rect 266636 198018 266688 198024
rect 266648 186386 266676 198018
rect 267936 193254 267964 211074
rect 267832 193248 267884 193254
rect 267752 193196 267832 193202
rect 267752 193190 267884 193196
rect 267924 193248 267976 193254
rect 267924 193190 267976 193196
rect 267752 193174 267872 193190
rect 267752 186386 267780 193174
rect 266636 186380 266688 186386
rect 266636 186322 266688 186328
rect 267740 186380 267792 186386
rect 267740 186322 267792 186328
rect 266728 186244 266780 186250
rect 266728 186186 266780 186192
rect 266740 178786 266768 186186
rect 267740 183592 267792 183598
rect 267740 183534 267792 183540
rect 266740 178758 266860 178786
rect 266832 173942 266860 178758
rect 266636 173936 266688 173942
rect 266636 173878 266688 173884
rect 266820 173936 266872 173942
rect 266820 173878 266872 173884
rect 266648 167634 266676 173878
rect 267752 171170 267780 183534
rect 267752 171142 267872 171170
rect 267844 171086 267872 171142
rect 267832 171080 267884 171086
rect 267832 171022 267884 171028
rect 266648 167606 266768 167634
rect 266740 125594 266768 167606
rect 267832 162784 267884 162790
rect 267832 162726 267884 162732
rect 267844 161430 267872 162726
rect 267832 161424 267884 161430
rect 267832 161366 267884 161372
rect 267832 151836 267884 151842
rect 267832 151778 267884 151784
rect 267844 147914 267872 151778
rect 267844 147886 267964 147914
rect 267936 147642 267964 147886
rect 267844 147614 267964 147642
rect 267844 133906 267872 147614
rect 267752 133878 267872 133906
rect 267752 125594 267780 133878
rect 266544 125588 266596 125594
rect 266544 125530 266596 125536
rect 266728 125588 266780 125594
rect 266728 125530 266780 125536
rect 267740 125588 267792 125594
rect 267740 125530 267792 125536
rect 267924 125588 267976 125594
rect 267924 125530 267976 125536
rect 266556 118674 266584 125530
rect 267936 120698 267964 125530
rect 267832 120692 267884 120698
rect 267832 120634 267884 120640
rect 267924 120692 267976 120698
rect 267924 120634 267976 120640
rect 266556 118646 266676 118674
rect 266648 108746 266676 118646
rect 267844 114510 267872 120634
rect 267832 114504 267884 114510
rect 267832 114446 267884 114452
rect 266648 108718 266768 108746
rect 266740 106282 266768 108718
rect 266728 106276 266780 106282
rect 266728 106218 266780 106224
rect 267832 106208 267884 106214
rect 267832 106150 267884 106156
rect 267844 104854 267872 106150
rect 267832 104848 267884 104854
rect 267832 104790 267884 104796
rect 266636 96688 266688 96694
rect 266636 96630 266688 96636
rect 266648 91746 266676 96630
rect 267924 95260 267976 95266
rect 267924 95202 267976 95208
rect 267936 92478 267964 95202
rect 267924 92472 267976 92478
rect 267924 92414 267976 92420
rect 268108 92472 268160 92478
rect 268108 92414 268160 92420
rect 266556 91718 266676 91746
rect 266556 89706 266584 91718
rect 266556 89678 266676 89706
rect 266648 77314 266676 89678
rect 268120 82929 268148 92414
rect 267830 82920 267886 82929
rect 267830 82855 267886 82864
rect 268106 82920 268162 82929
rect 268106 82855 268162 82864
rect 267844 82822 267872 82855
rect 267832 82816 267884 82822
rect 267832 82758 267884 82764
rect 268016 82816 268068 82822
rect 268016 82758 268068 82764
rect 268028 81433 268056 82758
rect 267830 81424 267886 81433
rect 267830 81359 267886 81368
rect 268014 81424 268070 81433
rect 268014 81359 268070 81368
rect 266636 77308 266688 77314
rect 266636 77250 266688 77256
rect 266728 77308 266780 77314
rect 266728 77250 266780 77256
rect 266740 74526 266768 77250
rect 266728 74520 266780 74526
rect 266728 74462 266780 74468
rect 267844 71806 267872 81359
rect 267832 71800 267884 71806
rect 267832 71742 267884 71748
rect 268016 71800 268068 71806
rect 268016 71742 268068 71748
rect 266912 64932 266964 64938
rect 266912 64874 266964 64880
rect 266924 44198 266952 64874
rect 268028 62121 268056 71742
rect 267830 62112 267886 62121
rect 267830 62047 267886 62056
rect 268014 62112 268070 62121
rect 268014 62047 268070 62056
rect 267844 52494 267872 62047
rect 267832 52488 267884 52494
rect 267832 52430 267884 52436
rect 268016 52488 268068 52494
rect 268016 52430 268068 52436
rect 268028 46986 268056 52430
rect 268016 46980 268068 46986
rect 268016 46922 268068 46928
rect 267740 46912 267792 46918
rect 267740 46854 267792 46860
rect 266636 44192 266688 44198
rect 266636 44134 266688 44140
rect 266912 44192 266964 44198
rect 266912 44134 266964 44140
rect 266648 41410 266676 44134
rect 266636 41404 266688 41410
rect 266636 41346 266688 41352
rect 267752 40202 267780 46854
rect 267752 40174 267964 40202
rect 266636 34468 266688 34474
rect 266636 34410 266688 34416
rect 266648 31770 266676 34410
rect 266648 31742 266768 31770
rect 266740 24954 266768 31742
rect 267936 31090 267964 40174
rect 267844 31062 267964 31090
rect 266728 24948 266780 24954
rect 266728 24890 266780 24896
rect 266636 24812 266688 24818
rect 266636 24754 266688 24760
rect 266452 14748 266504 14754
rect 266452 14690 266504 14696
rect 266648 10606 266676 24754
rect 267844 18086 267872 31062
rect 268016 22160 268068 22166
rect 268016 22102 268068 22108
rect 267832 18080 267884 18086
rect 267832 18022 267884 18028
rect 267740 18012 267792 18018
rect 267740 17954 267792 17960
rect 267752 10674 267780 17954
rect 268028 10878 268056 22102
rect 268016 10872 268068 10878
rect 268016 10814 268068 10820
rect 267740 10668 267792 10674
rect 267740 10610 267792 10616
rect 266636 10600 266688 10606
rect 266636 10542 266688 10548
rect 265164 8288 265216 8294
rect 265164 8230 265216 8236
rect 263876 8220 263928 8226
rect 263876 8162 263928 8168
rect 267004 8220 267056 8226
rect 267004 8162 267056 8168
rect 262404 8152 262456 8158
rect 262404 8094 262456 8100
rect 263416 8152 263468 8158
rect 263416 8094 263468 8100
rect 262220 3596 262272 3602
rect 262220 3538 262272 3544
rect 261484 2848 261536 2854
rect 261484 2790 261536 2796
rect 261024 1284 261076 1290
rect 261024 1226 261076 1232
rect 261036 480 261064 1226
rect 262232 480 262260 3538
rect 263428 480 263456 8094
rect 264612 3868 264664 3874
rect 264612 3810 264664 3816
rect 264624 480 264652 3810
rect 265808 3664 265860 3670
rect 265808 3606 265860 3612
rect 265820 480 265848 3606
rect 267016 480 267044 8162
rect 269040 4146 269068 337350
rect 269224 14822 269252 340054
rect 269684 337482 269712 340068
rect 269868 340054 270158 340082
rect 269672 337476 269724 337482
rect 269672 337418 269724 337424
rect 269868 335594 269896 340054
rect 269316 335566 269896 335594
rect 269212 14816 269264 14822
rect 269212 14758 269264 14764
rect 269316 10742 269344 335566
rect 270500 172508 270552 172514
rect 270500 172450 270552 172456
rect 270512 162897 270540 172450
rect 270498 162888 270554 162897
rect 270498 162823 270554 162832
rect 270500 130416 270552 130422
rect 270500 130358 270552 130364
rect 270512 125633 270540 130358
rect 270498 125624 270554 125633
rect 270498 125559 270554 125568
rect 270406 110528 270462 110537
rect 270406 110463 270408 110472
rect 270460 110463 270462 110472
rect 270408 110434 270460 110440
rect 270500 22228 270552 22234
rect 270500 22170 270552 22176
rect 270512 10810 270540 22170
rect 270604 16658 270632 340068
rect 271156 337142 271184 340068
rect 271248 340054 271630 340082
rect 271984 340054 272090 340082
rect 271144 337136 271196 337142
rect 271144 337078 271196 337084
rect 271248 334354 271276 340054
rect 271788 337476 271840 337482
rect 271788 337418 271840 337424
rect 271328 337340 271380 337346
rect 271328 337282 271380 337288
rect 270776 334348 270828 334354
rect 270776 334290 270828 334296
rect 271236 334348 271288 334354
rect 271236 334290 271288 334296
rect 270788 308394 270816 334290
rect 271340 334234 271368 337282
rect 271156 334206 271368 334234
rect 270788 308366 271000 308394
rect 270972 294001 271000 308366
rect 270774 293992 270830 294001
rect 270774 293927 270830 293936
rect 270958 293992 271014 294001
rect 270958 293927 271014 293936
rect 270788 292534 270816 293927
rect 270776 292528 270828 292534
rect 270776 292470 270828 292476
rect 270776 285660 270828 285666
rect 270776 285602 270828 285608
rect 270788 273306 270816 285602
rect 270696 273278 270816 273306
rect 270696 263634 270724 273278
rect 270684 263628 270736 263634
rect 270684 263570 270736 263576
rect 270684 263492 270736 263498
rect 270684 263434 270736 263440
rect 270696 260846 270724 263434
rect 270684 260840 270736 260846
rect 270684 260782 270736 260788
rect 270776 251116 270828 251122
rect 270776 251058 270828 251064
rect 270788 241602 270816 251058
rect 270776 241596 270828 241602
rect 270776 241538 270828 241544
rect 270684 241460 270736 241466
rect 270684 241402 270736 241408
rect 270696 240145 270724 241402
rect 270682 240136 270738 240145
rect 270682 240071 270738 240080
rect 270682 240000 270738 240009
rect 270682 239935 270738 239944
rect 270696 225010 270724 239935
rect 270684 225004 270736 225010
rect 270684 224946 270736 224952
rect 270684 220856 270736 220862
rect 270684 220798 270736 220804
rect 270696 205698 270724 220798
rect 270684 205692 270736 205698
rect 270684 205634 270736 205640
rect 270684 202904 270736 202910
rect 270682 202872 270684 202881
rect 270736 202872 270738 202881
rect 270682 202807 270738 202816
rect 270682 202736 270738 202745
rect 270682 202671 270738 202680
rect 270696 186386 270724 202671
rect 270684 186380 270736 186386
rect 270684 186322 270736 186328
rect 270684 183592 270736 183598
rect 270682 183560 270684 183569
rect 270736 183560 270738 183569
rect 270682 183495 270738 183504
rect 270866 183424 270922 183433
rect 270866 183359 270922 183368
rect 270880 176474 270908 183359
rect 270788 176446 270908 176474
rect 270788 172514 270816 176446
rect 270776 172508 270828 172514
rect 270776 172450 270828 172456
rect 270682 162888 270738 162897
rect 270682 162823 270738 162832
rect 270696 144906 270724 162823
rect 270684 144900 270736 144906
rect 270684 144842 270736 144848
rect 270684 140004 270736 140010
rect 270684 139946 270736 139952
rect 270696 130422 270724 139946
rect 270684 130416 270736 130422
rect 270684 130358 270736 130364
rect 270682 125624 270738 125633
rect 270682 125559 270684 125568
rect 270736 125559 270738 125568
rect 270684 125530 270736 125536
rect 270684 120692 270736 120698
rect 270684 120634 270736 120640
rect 270696 106282 270724 120634
rect 270684 106276 270736 106282
rect 270684 106218 270736 106224
rect 270684 106140 270736 106146
rect 270684 106082 270736 106088
rect 270696 100094 270724 106082
rect 270684 100088 270736 100094
rect 270684 100030 270736 100036
rect 270868 100088 270920 100094
rect 270868 100030 270920 100036
rect 270880 95282 270908 100030
rect 270788 95254 270908 95282
rect 270788 84182 270816 95254
rect 270776 84176 270828 84182
rect 270776 84118 270828 84124
rect 270776 74588 270828 74594
rect 270776 74530 270828 74536
rect 270788 66314 270816 74530
rect 270696 66286 270816 66314
rect 270696 66230 270724 66286
rect 270684 66224 270736 66230
rect 270684 66166 270736 66172
rect 270684 42900 270736 42906
rect 270684 42842 270736 42848
rect 270696 29730 270724 42842
rect 270696 29702 270816 29730
rect 270788 22234 270816 29702
rect 270776 22228 270828 22234
rect 270776 22170 270828 22176
rect 270592 16652 270644 16658
rect 270592 16594 270644 16600
rect 270592 16516 270644 16522
rect 270592 16458 270644 16464
rect 270604 14890 270632 16458
rect 270592 14884 270644 14890
rect 270592 14826 270644 14832
rect 270500 10804 270552 10810
rect 270500 10746 270552 10752
rect 269304 10736 269356 10742
rect 269304 10678 269356 10684
rect 270500 8288 270552 8294
rect 270500 8230 270552 8236
rect 268108 4140 268160 4146
rect 268108 4082 268160 4088
rect 269028 4140 269080 4146
rect 269028 4082 269080 4088
rect 268120 480 268148 4082
rect 269304 3256 269356 3262
rect 269304 3198 269356 3204
rect 269316 480 269344 3198
rect 270512 480 270540 8230
rect 271156 4418 271184 334206
rect 271144 4412 271196 4418
rect 271144 4354 271196 4360
rect 271800 626 271828 337418
rect 271984 14958 272012 340054
rect 272628 337278 272656 340068
rect 272720 340054 273102 340082
rect 273364 340054 273562 340082
rect 272616 337272 272668 337278
rect 272616 337214 272668 337220
rect 272720 334354 272748 340054
rect 272800 337272 272852 337278
rect 272800 337214 272852 337220
rect 272248 334348 272300 334354
rect 272248 334290 272300 334296
rect 272708 334348 272760 334354
rect 272708 334290 272760 334296
rect 272260 311982 272288 334290
rect 272812 334234 272840 337214
rect 272536 334206 272840 334234
rect 272248 311976 272300 311982
rect 272248 311918 272300 311924
rect 272248 311840 272300 311846
rect 272248 311782 272300 311788
rect 272260 303634 272288 311782
rect 272260 303606 272380 303634
rect 272352 295458 272380 303606
rect 272340 295452 272392 295458
rect 272340 295394 272392 295400
rect 272248 295316 272300 295322
rect 272248 295258 272300 295264
rect 272260 265690 272288 295258
rect 272168 265662 272288 265690
rect 272168 260846 272196 265662
rect 272156 260840 272208 260846
rect 272156 260782 272208 260788
rect 272156 260704 272208 260710
rect 272156 260646 272208 260652
rect 272168 244458 272196 260646
rect 272156 244452 272208 244458
rect 272156 244394 272208 244400
rect 272156 241596 272208 241602
rect 272156 241538 272208 241544
rect 272168 240106 272196 241538
rect 272156 240100 272208 240106
rect 272156 240042 272208 240048
rect 272248 234524 272300 234530
rect 272248 234466 272300 234472
rect 272260 230489 272288 234466
rect 272246 230480 272302 230489
rect 272246 230415 272302 230424
rect 272430 230480 272486 230489
rect 272430 230415 272486 230424
rect 272444 224754 272472 230415
rect 272260 224726 272472 224754
rect 272260 215370 272288 224726
rect 272168 215342 272288 215370
rect 272168 202881 272196 215342
rect 272154 202872 272210 202881
rect 272154 202807 272210 202816
rect 272246 190496 272302 190505
rect 272246 190431 272302 190440
rect 272260 180810 272288 190431
rect 272248 180804 272300 180810
rect 272248 180746 272300 180752
rect 272432 180804 272484 180810
rect 272432 180746 272484 180752
rect 272444 162897 272472 180746
rect 272246 162888 272302 162897
rect 272246 162823 272302 162832
rect 272430 162888 272486 162897
rect 272430 162823 272486 162832
rect 272260 153270 272288 162823
rect 272156 153264 272208 153270
rect 272156 153206 272208 153212
rect 272248 153264 272300 153270
rect 272248 153206 272300 153212
rect 272168 144906 272196 153206
rect 272156 144900 272208 144906
rect 272156 144842 272208 144848
rect 272248 144900 272300 144906
rect 272248 144842 272300 144848
rect 272260 139890 272288 144842
rect 272168 139862 272288 139890
rect 272168 130422 272196 139862
rect 272156 130416 272208 130422
rect 272156 130358 272208 130364
rect 272340 130416 272392 130422
rect 272340 130358 272392 130364
rect 272352 125633 272380 130358
rect 272154 125624 272210 125633
rect 272154 125559 272156 125568
rect 272208 125559 272210 125568
rect 272338 125624 272394 125633
rect 272338 125559 272394 125568
rect 272156 125530 272208 125536
rect 272156 120692 272208 120698
rect 272156 120634 272208 120640
rect 272168 109070 272196 120634
rect 272156 109064 272208 109070
rect 272156 109006 272208 109012
rect 272156 108928 272208 108934
rect 272156 108870 272208 108876
rect 272168 106282 272196 108870
rect 272156 106276 272208 106282
rect 272156 106218 272208 106224
rect 272248 106276 272300 106282
rect 272248 106218 272300 106224
rect 272260 104854 272288 106218
rect 272248 104848 272300 104854
rect 272248 104790 272300 104796
rect 272340 96552 272392 96558
rect 272340 96494 272392 96500
rect 272352 77246 272380 96494
rect 272248 77240 272300 77246
rect 272248 77182 272300 77188
rect 272340 77240 272392 77246
rect 272340 77182 272392 77188
rect 272260 75886 272288 77182
rect 272248 75880 272300 75886
rect 272248 75822 272300 75828
rect 272156 66292 272208 66298
rect 272156 66234 272208 66240
rect 272168 60790 272196 66234
rect 272156 60784 272208 60790
rect 272156 60726 272208 60732
rect 272156 60648 272208 60654
rect 272156 60590 272208 60596
rect 272168 44198 272196 60590
rect 272156 44192 272208 44198
rect 272156 44134 272208 44140
rect 272432 44192 272484 44198
rect 272432 44134 272484 44140
rect 272444 34542 272472 44134
rect 272248 34536 272300 34542
rect 272248 34478 272300 34484
rect 272432 34536 272484 34542
rect 272432 34478 272484 34484
rect 272260 22166 272288 34478
rect 272248 22160 272300 22166
rect 272248 22102 272300 22108
rect 271972 14952 272024 14958
rect 271972 14894 272024 14900
rect 272536 4350 272564 334206
rect 273168 63708 273220 63714
rect 273168 63650 273220 63656
rect 273180 63617 273208 63650
rect 273166 63608 273222 63617
rect 273166 63543 273222 63552
rect 273364 15026 273392 340054
rect 274100 337006 274128 340068
rect 274284 340054 274574 340082
rect 274744 340054 275034 340082
rect 274088 337000 274140 337006
rect 274088 336942 274140 336948
rect 274284 335628 274312 340054
rect 273640 335600 274312 335628
rect 273640 313478 273668 335600
rect 273628 313472 273680 313478
rect 273628 313414 273680 313420
rect 273444 311908 273496 311914
rect 273444 311850 273496 311856
rect 273456 311794 273484 311850
rect 273456 311766 273576 311794
rect 273548 293162 273576 311766
rect 273548 293134 273668 293162
rect 273640 282826 273668 293134
rect 273548 282798 273668 282826
rect 273548 280158 273576 282798
rect 273536 280152 273588 280158
rect 273536 280094 273588 280100
rect 273628 280152 273680 280158
rect 273628 280094 273680 280100
rect 273640 263514 273668 280094
rect 273548 263486 273668 263514
rect 273548 260846 273576 263486
rect 273536 260840 273588 260846
rect 273536 260782 273588 260788
rect 273628 260840 273680 260846
rect 273628 260782 273680 260788
rect 273640 244202 273668 260782
rect 273548 244174 273668 244202
rect 273548 240106 273576 244174
rect 273536 240100 273588 240106
rect 273536 240042 273588 240048
rect 273628 240100 273680 240106
rect 273628 240042 273680 240048
rect 273640 224890 273668 240042
rect 273548 224862 273668 224890
rect 273548 215370 273576 224862
rect 273456 215342 273576 215370
rect 273456 215286 273484 215342
rect 273444 215280 273496 215286
rect 273444 215222 273496 215228
rect 273628 215280 273680 215286
rect 273628 215222 273680 215228
rect 273640 207754 273668 215222
rect 273548 207726 273668 207754
rect 273548 202842 273576 207726
rect 273536 202836 273588 202842
rect 273536 202778 273588 202784
rect 273628 202836 273680 202842
rect 273628 202778 273680 202784
rect 273640 186266 273668 202778
rect 273548 186238 273668 186266
rect 273548 183530 273576 186238
rect 273536 183524 273588 183530
rect 273536 183466 273588 183472
rect 273628 183524 273680 183530
rect 273628 183466 273680 183472
rect 273640 157434 273668 183466
rect 273456 157406 273668 157434
rect 273456 157298 273484 157406
rect 273456 157270 273576 157298
rect 273548 137850 273576 157270
rect 273548 137822 273668 137850
rect 273640 128330 273668 137822
rect 273548 128302 273668 128330
rect 273548 118794 273576 128302
rect 273536 118788 273588 118794
rect 273536 118730 273588 118736
rect 273536 118652 273588 118658
rect 273536 118594 273588 118600
rect 273548 104854 273576 118594
rect 273536 104848 273588 104854
rect 273536 104790 273588 104796
rect 273628 95260 273680 95266
rect 273628 95202 273680 95208
rect 273640 70514 273668 95202
rect 273628 70508 273680 70514
rect 273628 70450 273680 70456
rect 273536 67652 273588 67658
rect 273536 67594 273588 67600
rect 273548 60738 273576 67594
rect 273456 60722 273576 60738
rect 273444 60716 273576 60722
rect 273496 60710 273576 60716
rect 273628 60716 273680 60722
rect 273444 60658 273496 60664
rect 273628 60658 273680 60664
rect 273640 51134 273668 60658
rect 273628 51128 273680 51134
rect 273628 51070 273680 51076
rect 273536 51060 273588 51066
rect 273536 51002 273588 51008
rect 273548 48278 273576 51002
rect 273536 48272 273588 48278
rect 273536 48214 273588 48220
rect 273536 38684 273588 38690
rect 273536 38626 273588 38632
rect 273548 22114 273576 38626
rect 273456 22086 273576 22114
rect 273456 16590 273484 22086
rect 273444 16584 273496 16590
rect 273444 16526 273496 16532
rect 274744 15094 274772 340054
rect 275572 337550 275600 340068
rect 275560 337544 275612 337550
rect 275560 337486 275612 337492
rect 275928 337544 275980 337550
rect 275928 337486 275980 337492
rect 274732 15088 274784 15094
rect 274732 15030 274784 15036
rect 273352 15020 273404 15026
rect 273352 14962 273404 14968
rect 274088 6180 274140 6186
rect 274088 6122 274140 6128
rect 272524 4344 272576 4350
rect 272524 4286 272576 4292
rect 272892 3188 272944 3194
rect 272892 3130 272944 3136
rect 271708 598 271828 626
rect 271708 480 271736 598
rect 272904 480 272932 3130
rect 274100 480 274128 6122
rect 275940 2922 275968 337486
rect 276032 11014 276060 340068
rect 276124 340054 276506 340082
rect 276124 15162 276152 340054
rect 277044 337686 277072 340068
rect 277518 340054 277624 340082
rect 277032 337680 277084 337686
rect 277032 337622 277084 337628
rect 276112 15156 276164 15162
rect 276112 15098 276164 15104
rect 276020 11008 276072 11014
rect 276020 10950 276072 10956
rect 277596 10266 277624 340054
rect 277688 340054 277978 340082
rect 277688 14414 277716 340054
rect 278516 336870 278544 340068
rect 278792 340054 278990 340082
rect 279068 340054 279450 340082
rect 278504 336864 278556 336870
rect 278504 336806 278556 336812
rect 278792 334830 278820 340054
rect 278780 334824 278832 334830
rect 278780 334766 278832 334772
rect 278964 334824 279016 334830
rect 278964 334766 279016 334772
rect 278872 328500 278924 328506
rect 278872 328442 278924 328448
rect 278686 157720 278742 157729
rect 278686 157655 278742 157664
rect 278700 157593 278728 157655
rect 278686 157584 278742 157593
rect 278686 157519 278742 157528
rect 278884 157434 278912 328442
rect 278792 157406 278912 157434
rect 278792 157298 278820 157406
rect 278792 157270 278912 157298
rect 278686 110528 278742 110537
rect 278686 110463 278688 110472
rect 278740 110463 278742 110472
rect 278688 110434 278740 110440
rect 278884 109154 278912 157270
rect 278792 109126 278912 109154
rect 278792 109002 278820 109126
rect 278780 108996 278832 109002
rect 278780 108938 278832 108944
rect 278872 99408 278924 99414
rect 278872 99350 278924 99356
rect 278884 80186 278912 99350
rect 278792 80158 278912 80186
rect 278686 63744 278742 63753
rect 278686 63679 278688 63688
rect 278740 63679 278742 63688
rect 278688 63650 278740 63656
rect 278792 41290 278820 80158
rect 278792 41262 278912 41290
rect 277676 14408 277728 14414
rect 277676 14350 277728 14356
rect 278884 14346 278912 41262
rect 278872 14340 278924 14346
rect 278872 14282 278924 14288
rect 277584 10260 277636 10266
rect 277584 10202 277636 10208
rect 278976 10198 279004 334766
rect 279068 328506 279096 340054
rect 279988 337618 280016 340068
rect 280356 340054 280462 340082
rect 280632 340054 280922 340082
rect 281184 340054 281474 340082
rect 281644 340054 281934 340082
rect 282104 340054 282394 340082
rect 282946 340054 283144 340082
rect 279976 337612 280028 337618
rect 279976 337554 280028 337560
rect 280252 335640 280304 335646
rect 280252 335582 280304 335588
rect 279056 328500 279108 328506
rect 279056 328442 279108 328448
rect 280066 110800 280122 110809
rect 280066 110735 280122 110744
rect 280080 110537 280108 110735
rect 280066 110528 280122 110537
rect 280066 110463 280122 110472
rect 279056 108996 279108 109002
rect 279056 108938 279108 108944
rect 279068 99414 279096 108938
rect 279056 99408 279108 99414
rect 279056 99350 279108 99356
rect 280264 14278 280292 335582
rect 280252 14272 280304 14278
rect 280252 14214 280304 14220
rect 278964 10192 279016 10198
rect 278964 10134 279016 10140
rect 280356 10130 280384 340054
rect 280632 335646 280660 340054
rect 281184 336802 281212 340054
rect 281448 337612 281500 337618
rect 281448 337554 281500 337560
rect 281172 336796 281224 336802
rect 281172 336738 281224 336744
rect 280620 335640 280672 335646
rect 280620 335582 280672 335588
rect 280344 10124 280396 10130
rect 280344 10066 280396 10072
rect 280068 6248 280120 6254
rect 280068 6190 280120 6196
rect 276480 3256 276532 3262
rect 276480 3198 276532 3204
rect 275284 2916 275336 2922
rect 275284 2858 275336 2864
rect 275928 2916 275980 2922
rect 275928 2858 275980 2864
rect 275296 480 275324 2858
rect 276492 480 276520 3198
rect 277676 3120 277728 3126
rect 277676 3062 277728 3068
rect 278872 3120 278924 3126
rect 278872 3062 278924 3068
rect 277688 480 277716 3062
rect 278884 480 278912 3062
rect 280080 480 280108 6190
rect 281460 610 281488 337554
rect 281540 335640 281592 335646
rect 281540 335582 281592 335588
rect 281552 11898 281580 335582
rect 281540 11892 281592 11898
rect 281540 11834 281592 11840
rect 281644 11830 281672 340054
rect 282104 335646 282132 340054
rect 282092 335640 282144 335646
rect 282092 335582 282144 335588
rect 283012 335640 283064 335646
rect 283012 335582 283064 335588
rect 282642 157448 282698 157457
rect 282642 157383 282644 157392
rect 282696 157383 282698 157392
rect 282644 157354 282696 157360
rect 282918 87272 282974 87281
rect 282918 87207 282974 87216
rect 282826 87136 282882 87145
rect 282932 87122 282960 87207
rect 282882 87094 282960 87122
rect 282826 87071 282882 87080
rect 282734 40216 282790 40225
rect 282918 40216 282974 40225
rect 282790 40174 282918 40202
rect 282734 40151 282790 40160
rect 282918 40151 282974 40160
rect 281632 11824 281684 11830
rect 281632 11766 281684 11772
rect 283024 6662 283052 335582
rect 283116 7585 283144 340054
rect 283208 340054 283406 340082
rect 283576 340054 283866 340082
rect 283102 7576 283158 7585
rect 283102 7511 283158 7520
rect 283012 6656 283064 6662
rect 283012 6598 283064 6604
rect 283208 5370 283236 340054
rect 283576 335646 283604 340054
rect 284404 338094 284432 340068
rect 284588 340054 284878 340082
rect 285140 340054 285338 340082
rect 285798 340054 285904 340082
rect 284392 338088 284444 338094
rect 284392 338030 284444 338036
rect 283564 335640 283616 335646
rect 283564 335582 283616 335588
rect 284484 335232 284536 335238
rect 284484 335174 284536 335180
rect 284300 331968 284352 331974
rect 284300 331910 284352 331916
rect 284312 5438 284340 331910
rect 284392 283620 284444 283626
rect 284392 283562 284444 283568
rect 284404 273970 284432 283562
rect 284392 273964 284444 273970
rect 284392 273906 284444 273912
rect 284496 8945 284524 335174
rect 284588 331974 284616 340054
rect 285140 332586 285168 340054
rect 285588 337680 285640 337686
rect 285588 337622 285640 337628
rect 284668 332580 284720 332586
rect 284668 332522 284720 332528
rect 285128 332580 285180 332586
rect 285128 332522 285180 332528
rect 284576 331968 284628 331974
rect 284576 331910 284628 331916
rect 284680 321314 284708 332522
rect 284680 321286 284800 321314
rect 284772 318782 284800 321286
rect 284760 318776 284812 318782
rect 284760 318718 284812 318724
rect 284944 314220 284996 314226
rect 284944 314162 284996 314168
rect 284956 306377 284984 314162
rect 284758 306368 284814 306377
rect 284758 306303 284814 306312
rect 284942 306368 284998 306377
rect 284942 306303 284998 306312
rect 284772 296750 284800 306303
rect 284760 296744 284812 296750
rect 284666 296712 284722 296721
rect 284852 296744 284904 296750
rect 284760 296686 284812 296692
rect 284850 296712 284852 296721
rect 284904 296712 284906 296721
rect 284666 296647 284722 296656
rect 284850 296647 284906 296656
rect 284680 288130 284708 296647
rect 284680 288102 284892 288130
rect 284864 283626 284892 288102
rect 284852 283620 284904 283626
rect 284852 283562 284904 283568
rect 284760 273964 284812 273970
rect 284760 273906 284812 273912
rect 284772 269113 284800 273906
rect 284574 269104 284630 269113
rect 284574 269039 284630 269048
rect 284758 269104 284814 269113
rect 284758 269039 284814 269048
rect 284588 259486 284616 269039
rect 284576 259480 284628 259486
rect 284576 259422 284628 259428
rect 284760 259480 284812 259486
rect 284760 259422 284812 259428
rect 284772 249898 284800 259422
rect 284668 249892 284720 249898
rect 284668 249834 284720 249840
rect 284760 249892 284812 249898
rect 284760 249834 284812 249840
rect 284680 249801 284708 249834
rect 284666 249792 284722 249801
rect 284666 249727 284722 249736
rect 284942 249792 284998 249801
rect 284942 249727 284998 249736
rect 284956 240174 284984 249727
rect 284760 240168 284812 240174
rect 284760 240110 284812 240116
rect 284944 240168 284996 240174
rect 284944 240110 284996 240116
rect 284772 222222 284800 240110
rect 284760 222216 284812 222222
rect 284760 222158 284812 222164
rect 284760 222080 284812 222086
rect 284760 222022 284812 222028
rect 284772 212566 284800 222022
rect 284760 212560 284812 212566
rect 284760 212502 284812 212508
rect 284944 212492 284996 212498
rect 284944 212434 284996 212440
rect 284956 201521 284984 212434
rect 284758 201512 284814 201521
rect 284758 201447 284814 201456
rect 284942 201512 284998 201521
rect 284942 201447 284998 201456
rect 284772 183598 284800 201447
rect 284760 183592 284812 183598
rect 284760 183534 284812 183540
rect 284760 183456 284812 183462
rect 284760 183398 284812 183404
rect 284772 180810 284800 183398
rect 284760 180804 284812 180810
rect 284760 180746 284812 180752
rect 284944 171148 284996 171154
rect 284944 171090 284996 171096
rect 284956 162926 284984 171090
rect 284760 162920 284812 162926
rect 284760 162862 284812 162868
rect 284944 162920 284996 162926
rect 284944 162862 284996 162868
rect 284772 135561 284800 162862
rect 284758 135552 284814 135561
rect 284758 135487 284814 135496
rect 284666 135280 284722 135289
rect 284666 135215 284722 135224
rect 284680 132462 284708 135215
rect 284668 132456 284720 132462
rect 284668 132398 284720 132404
rect 284668 126948 284720 126954
rect 284668 126890 284720 126896
rect 284680 122806 284708 126890
rect 284668 122800 284720 122806
rect 284668 122742 284720 122748
rect 284852 122800 284904 122806
rect 284852 122742 284904 122748
rect 284864 110922 284892 122742
rect 284772 110894 284892 110922
rect 284772 90234 284800 110894
rect 284760 90228 284812 90234
rect 284760 90170 284812 90176
rect 284760 85604 284812 85610
rect 284760 85546 284812 85552
rect 284772 84182 284800 85546
rect 284760 84176 284812 84182
rect 284760 84118 284812 84124
rect 284852 75812 284904 75818
rect 284852 75754 284904 75760
rect 284864 58002 284892 75754
rect 284760 57996 284812 58002
rect 284760 57938 284812 57944
rect 284852 57996 284904 58002
rect 284852 57938 284904 57944
rect 284772 53122 284800 57938
rect 284680 53094 284800 53122
rect 284680 44742 284708 53094
rect 284668 44736 284720 44742
rect 284668 44678 284720 44684
rect 284760 29028 284812 29034
rect 284760 28970 284812 28976
rect 284772 22114 284800 28970
rect 284772 22086 284892 22114
rect 284864 18086 284892 22086
rect 284852 18080 284904 18086
rect 284852 18022 284904 18028
rect 284668 18012 284720 18018
rect 284668 17954 284720 17960
rect 284680 13138 284708 17954
rect 284588 13110 284708 13138
rect 284482 8936 284538 8945
rect 284482 8871 284538 8880
rect 284588 7546 284616 13110
rect 284576 7540 284628 7546
rect 284576 7482 284628 7488
rect 284300 5432 284352 5438
rect 284300 5374 284352 5380
rect 283196 5364 283248 5370
rect 283196 5306 283248 5312
rect 283656 5296 283708 5302
rect 283656 5238 283708 5244
rect 282460 3936 282512 3942
rect 282460 3878 282512 3884
rect 281264 604 281316 610
rect 281264 546 281316 552
rect 281448 604 281500 610
rect 281448 546 281500 552
rect 281276 480 281304 546
rect 282472 480 282500 3878
rect 283668 480 283696 5238
rect 285600 4146 285628 337622
rect 285680 335640 285732 335646
rect 285680 335582 285732 335588
rect 285692 5506 285720 335582
rect 285770 202872 285826 202881
rect 285770 202807 285826 202816
rect 285784 198082 285812 202807
rect 285772 198076 285824 198082
rect 285772 198018 285824 198024
rect 285772 162852 285824 162858
rect 285772 162794 285824 162800
rect 285784 153241 285812 162794
rect 285770 153232 285826 153241
rect 285770 153167 285826 153176
rect 285876 9314 285904 340054
rect 285968 340054 286350 340082
rect 286612 340054 286810 340082
rect 287164 340054 287270 340082
rect 287348 340054 287822 340082
rect 287992 340054 288282 340082
rect 288544 340054 288742 340082
rect 289004 340054 289294 340082
rect 289464 340054 289754 340082
rect 289832 340054 290214 340082
rect 285968 335646 285996 340054
rect 286612 335646 286640 340054
rect 285956 335640 286008 335646
rect 285956 335582 286008 335588
rect 286048 335640 286100 335646
rect 286048 335582 286100 335588
rect 286600 335640 286652 335646
rect 286600 335582 286652 335588
rect 287060 335640 287112 335646
rect 287060 335582 287112 335588
rect 286060 321638 286088 335582
rect 286048 321632 286100 321638
rect 286048 321574 286100 321580
rect 285956 321564 286008 321570
rect 285956 321506 286008 321512
rect 285968 318782 285996 321506
rect 285956 318776 286008 318782
rect 285956 318718 286008 318724
rect 286140 318776 286192 318782
rect 286140 318718 286192 318724
rect 286152 313698 286180 318718
rect 286060 313670 286180 313698
rect 286060 299554 286088 313670
rect 285968 299526 286088 299554
rect 285968 298110 285996 299526
rect 285956 298104 286008 298110
rect 285956 298046 286008 298052
rect 285956 288448 286008 288454
rect 285956 288390 286008 288396
rect 285968 280158 285996 288390
rect 285956 280152 286008 280158
rect 285956 280094 286008 280100
rect 286140 280152 286192 280158
rect 286140 280094 286192 280100
rect 286152 279834 286180 280094
rect 286060 279806 286180 279834
rect 286060 261089 286088 279806
rect 286046 261080 286102 261089
rect 286046 261015 286102 261024
rect 285954 260944 286010 260953
rect 285954 260879 286010 260888
rect 285968 249830 285996 260879
rect 285956 249824 286008 249830
rect 286048 249824 286100 249830
rect 285956 249766 286008 249772
rect 286046 249792 286048 249801
rect 286100 249792 286102 249801
rect 286046 249727 286102 249736
rect 285954 249656 286010 249665
rect 285954 249591 286010 249600
rect 285968 245002 285996 249591
rect 285956 244996 286008 245002
rect 285956 244938 286008 244944
rect 285956 234524 286008 234530
rect 285956 234466 286008 234472
rect 285968 222193 285996 234466
rect 285954 222184 286010 222193
rect 285954 222119 286010 222128
rect 286138 222184 286194 222193
rect 286138 222119 286194 222128
rect 286152 220833 286180 222119
rect 285954 220824 286010 220833
rect 285954 220759 286010 220768
rect 286138 220824 286194 220833
rect 286138 220759 286194 220768
rect 285968 212242 285996 220759
rect 285968 212214 286180 212242
rect 286152 202910 286180 212214
rect 285956 202904 286008 202910
rect 285954 202872 285956 202881
rect 286140 202904 286192 202910
rect 286008 202872 286010 202881
rect 286140 202846 286192 202852
rect 285954 202807 286010 202816
rect 285956 198076 286008 198082
rect 285956 198018 286008 198024
rect 285968 183569 285996 198018
rect 285954 183560 286010 183569
rect 285954 183495 286010 183504
rect 285954 183424 286010 183433
rect 285954 183359 286010 183368
rect 285968 162858 285996 183359
rect 285956 162852 286008 162858
rect 285956 162794 286008 162800
rect 285954 153232 286010 153241
rect 285954 153167 285956 153176
rect 286008 153167 286010 153176
rect 286048 153196 286100 153202
rect 285956 153138 286008 153144
rect 286048 153138 286100 153144
rect 286060 144650 286088 153138
rect 286060 144622 286180 144650
rect 286152 135946 286180 144622
rect 285968 135918 286180 135946
rect 285968 113098 285996 135918
rect 285968 113070 286088 113098
rect 286060 103737 286088 113070
rect 286046 103728 286102 103737
rect 286046 103663 286102 103672
rect 285954 103592 286010 103601
rect 285954 103527 286010 103536
rect 285968 103494 285996 103527
rect 285956 103488 286008 103494
rect 285956 103430 286008 103436
rect 286140 93900 286192 93906
rect 286140 93842 286192 93848
rect 286152 85678 286180 93842
rect 286140 85672 286192 85678
rect 286140 85614 286192 85620
rect 286048 85604 286100 85610
rect 286048 85546 286100 85552
rect 286060 78538 286088 85546
rect 286048 78532 286100 78538
rect 286048 78474 286100 78480
rect 285956 66292 286008 66298
rect 285956 66234 286008 66240
rect 285968 58002 285996 66234
rect 285956 57996 286008 58002
rect 285956 57938 286008 57944
rect 286048 57996 286100 58002
rect 286048 57938 286100 57944
rect 286060 56574 286088 57938
rect 286048 56568 286100 56574
rect 286048 56510 286100 56516
rect 285956 46980 286008 46986
rect 285956 46922 286008 46928
rect 285968 46866 285996 46922
rect 285968 46838 286088 46866
rect 286060 37398 286088 46838
rect 286048 37392 286100 37398
rect 286048 37334 286100 37340
rect 285956 37324 286008 37330
rect 285956 37266 286008 37272
rect 285968 29034 285996 37266
rect 285956 29028 286008 29034
rect 285956 28970 286008 28976
rect 286048 29028 286100 29034
rect 286048 28970 286100 28976
rect 286060 27606 286088 28970
rect 286048 27600 286100 27606
rect 286048 27542 286100 27548
rect 285956 18012 286008 18018
rect 285956 17954 286008 17960
rect 285864 9308 285916 9314
rect 285864 9250 285916 9256
rect 285968 7478 285996 17954
rect 285956 7472 286008 7478
rect 285956 7414 286008 7420
rect 287072 7410 287100 335582
rect 287164 9382 287192 340054
rect 287348 11966 287376 340054
rect 287992 335646 288020 340054
rect 288256 337816 288308 337822
rect 288256 337758 288308 337764
rect 287980 335640 288032 335646
rect 287980 335582 288032 335588
rect 287336 11960 287388 11966
rect 287336 11902 287388 11908
rect 287152 9376 287204 9382
rect 287152 9318 287204 9324
rect 287060 7404 287112 7410
rect 287060 7346 287112 7352
rect 285680 5500 285732 5506
rect 285680 5442 285732 5448
rect 287152 5364 287204 5370
rect 287152 5306 287204 5312
rect 284760 4140 284812 4146
rect 284760 4082 284812 4088
rect 285588 4140 285640 4146
rect 285588 4082 285640 4088
rect 284772 480 284800 4082
rect 285956 3868 286008 3874
rect 285956 3810 286008 3816
rect 285968 480 285996 3810
rect 287164 480 287192 5306
rect 288268 626 288296 337758
rect 288440 335640 288492 335646
rect 288440 335582 288492 335588
rect 288346 16824 288402 16833
rect 288346 16759 288402 16768
rect 288360 16561 288388 16759
rect 288346 16552 288402 16561
rect 288346 16487 288402 16496
rect 288452 7342 288480 335582
rect 288544 10062 288572 340054
rect 289004 331242 289032 340054
rect 289464 335646 289492 340054
rect 289452 335640 289504 335646
rect 289452 335582 289504 335588
rect 289004 331214 289124 331242
rect 289096 328506 289124 331214
rect 288808 328500 288860 328506
rect 288808 328442 288860 328448
rect 289084 328500 289136 328506
rect 289084 328442 289136 328448
rect 288820 313954 288848 328442
rect 288624 313948 288676 313954
rect 288624 313890 288676 313896
rect 288808 313948 288860 313954
rect 288808 313890 288860 313896
rect 288636 299538 288664 313890
rect 288624 299532 288676 299538
rect 288624 299474 288676 299480
rect 288808 299532 288860 299538
rect 288808 299474 288860 299480
rect 288820 296698 288848 299474
rect 288728 296670 288848 296698
rect 288728 292602 288756 296670
rect 288716 292596 288768 292602
rect 288716 292538 288768 292544
rect 288808 292528 288860 292534
rect 288808 292470 288860 292476
rect 288820 280158 288848 292470
rect 288624 280152 288676 280158
rect 288624 280094 288676 280100
rect 288808 280152 288860 280158
rect 288808 280094 288860 280100
rect 288636 260914 288664 280094
rect 288624 260908 288676 260914
rect 288624 260850 288676 260856
rect 288808 260908 288860 260914
rect 288808 260850 288860 260856
rect 288820 253994 288848 260850
rect 288820 253966 288940 253994
rect 288912 238921 288940 253966
rect 288898 238912 288954 238921
rect 288898 238847 288954 238856
rect 289082 238504 289138 238513
rect 289082 238439 289138 238448
rect 289096 220862 289124 238439
rect 288900 220856 288952 220862
rect 288900 220798 288952 220804
rect 289084 220856 289136 220862
rect 289084 220798 289136 220804
rect 288912 212514 288940 220798
rect 288912 212486 289032 212514
rect 289004 205442 289032 212486
rect 288728 205414 289032 205442
rect 288728 193390 288756 205414
rect 288716 193384 288768 193390
rect 288716 193326 288768 193332
rect 288716 193248 288768 193254
rect 288716 193190 288768 193196
rect 288728 189038 288756 193190
rect 288716 189032 288768 189038
rect 288716 188974 288768 188980
rect 288900 179444 288952 179450
rect 288900 179386 288952 179392
rect 288912 161566 288940 179386
rect 288900 161560 288952 161566
rect 288900 161502 288952 161508
rect 288808 161424 288860 161430
rect 288808 161366 288860 161372
rect 288820 160070 288848 161366
rect 288716 160064 288768 160070
rect 288716 160006 288768 160012
rect 288808 160064 288860 160070
rect 288808 160006 288860 160012
rect 288728 155258 288756 160006
rect 288898 157448 288954 157457
rect 288898 157383 288900 157392
rect 288952 157383 288954 157392
rect 288900 157354 288952 157360
rect 288728 155230 288848 155258
rect 288820 142186 288848 155230
rect 288624 142180 288676 142186
rect 288624 142122 288676 142128
rect 288808 142180 288860 142186
rect 288808 142122 288860 142128
rect 288636 135674 288664 142122
rect 288636 135646 288848 135674
rect 288820 122874 288848 135646
rect 288808 122868 288860 122874
rect 288808 122810 288860 122816
rect 288808 121508 288860 121514
rect 288808 121450 288860 121456
rect 288820 119354 288848 121450
rect 288820 119326 288940 119354
rect 288912 104922 288940 119326
rect 288716 104916 288768 104922
rect 288716 104858 288768 104864
rect 288900 104916 288952 104922
rect 288900 104858 288952 104864
rect 288728 103494 288756 104858
rect 288716 103488 288768 103494
rect 288716 103430 288768 103436
rect 288808 103420 288860 103426
rect 288808 103362 288860 103368
rect 288820 75954 288848 103362
rect 288716 75948 288768 75954
rect 288716 75890 288768 75896
rect 288808 75948 288860 75954
rect 288808 75890 288860 75896
rect 288728 74526 288756 75890
rect 288716 74520 288768 74526
rect 288716 74462 288768 74468
rect 288992 74520 289044 74526
rect 288992 74462 289044 74468
rect 289004 48346 289032 74462
rect 288716 48340 288768 48346
rect 288716 48282 288768 48288
rect 288992 48340 289044 48346
rect 288992 48282 289044 48288
rect 288728 37262 288756 48282
rect 288716 37256 288768 37262
rect 288716 37198 288768 37204
rect 288808 27668 288860 27674
rect 288808 27610 288860 27616
rect 288820 26246 288848 27610
rect 288808 26240 288860 26246
rect 288808 26182 288860 26188
rect 288808 16652 288860 16658
rect 288808 16594 288860 16600
rect 288820 12034 288848 16594
rect 288808 12028 288860 12034
rect 288808 11970 288860 11976
rect 288532 10056 288584 10062
rect 288532 9998 288584 10004
rect 289832 9994 289860 340054
rect 290292 331242 290320 340190
rect 290464 337884 290516 337890
rect 290464 337826 290516 337832
rect 290108 331214 290320 331242
rect 290108 312610 290136 331214
rect 290108 312582 290320 312610
rect 290292 309074 290320 312582
rect 290200 309046 290320 309074
rect 290200 294642 290228 309046
rect 290004 294636 290056 294642
rect 290004 294578 290056 294584
rect 290188 294636 290240 294642
rect 290188 294578 290240 294584
rect 290016 289814 290044 294578
rect 290004 289808 290056 289814
rect 290004 289750 290056 289756
rect 290188 289808 290240 289814
rect 290188 289750 290240 289756
rect 290200 269142 290228 289750
rect 290096 269136 290148 269142
rect 290096 269078 290148 269084
rect 290188 269136 290240 269142
rect 290188 269078 290240 269084
rect 290108 251258 290136 269078
rect 290004 251252 290056 251258
rect 290004 251194 290056 251200
rect 290096 251252 290148 251258
rect 290096 251194 290148 251200
rect 290016 249762 290044 251194
rect 290004 249756 290056 249762
rect 290004 249698 290056 249704
rect 290188 249756 290240 249762
rect 290188 249698 290240 249704
rect 290200 240145 290228 249698
rect 290186 240136 290242 240145
rect 290186 240071 290242 240080
rect 290370 240136 290426 240145
rect 290370 240071 290426 240080
rect 290384 238746 290412 240071
rect 290372 238740 290424 238746
rect 290372 238682 290424 238688
rect 290372 230444 290424 230450
rect 290372 230386 290424 230392
rect 290384 220862 290412 230386
rect 290188 220856 290240 220862
rect 290188 220798 290240 220804
rect 290372 220856 290424 220862
rect 290372 220798 290424 220804
rect 290200 219434 290228 220798
rect 290188 219428 290240 219434
rect 290188 219370 290240 219376
rect 290188 212492 290240 212498
rect 290188 212434 290240 212440
rect 290200 209794 290228 212434
rect 290200 209766 290320 209794
rect 290292 201657 290320 209766
rect 290278 201648 290334 201657
rect 290278 201583 290334 201592
rect 290186 201512 290242 201521
rect 290186 201447 290242 201456
rect 290200 200122 290228 201447
rect 289912 200116 289964 200122
rect 289912 200058 289964 200064
rect 290188 200116 290240 200122
rect 290188 200058 290240 200064
rect 289924 190505 289952 200058
rect 289910 190496 289966 190505
rect 289910 190431 289966 190440
rect 290094 190496 290150 190505
rect 290094 190431 290150 190440
rect 290108 183546 290136 190431
rect 290016 183518 290136 183546
rect 290016 172689 290044 183518
rect 290002 172680 290058 172689
rect 290002 172615 290058 172624
rect 290002 172544 290058 172553
rect 290002 172479 290058 172488
rect 290016 161566 290044 172479
rect 290004 161560 290056 161566
rect 290004 161502 290056 161508
rect 290096 161492 290148 161498
rect 290096 161434 290148 161440
rect 290108 155258 290136 161434
rect 290108 155230 290320 155258
rect 290292 151722 290320 155230
rect 290200 151694 290320 151722
rect 290200 142186 290228 151694
rect 290096 142180 290148 142186
rect 290096 142122 290148 142128
rect 290188 142180 290240 142186
rect 290188 142122 290240 142128
rect 290108 132530 290136 142122
rect 290004 132524 290056 132530
rect 290004 132466 290056 132472
rect 290096 132524 290148 132530
rect 290096 132466 290148 132472
rect 290016 122806 290044 132466
rect 290004 122800 290056 122806
rect 290004 122742 290056 122748
rect 290004 113212 290056 113218
rect 290004 113154 290056 113160
rect 290016 95198 290044 113154
rect 290004 95192 290056 95198
rect 290004 95134 290056 95140
rect 290096 95192 290148 95198
rect 290096 95134 290148 95140
rect 290108 75954 290136 95134
rect 289912 75948 289964 75954
rect 289912 75890 289964 75896
rect 290096 75948 290148 75954
rect 290096 75890 290148 75896
rect 289924 75834 289952 75890
rect 289924 75806 290044 75834
rect 290016 12102 290044 75806
rect 290004 12096 290056 12102
rect 290004 12038 290056 12044
rect 289820 9988 289872 9994
rect 289820 9930 289872 9936
rect 288440 7336 288492 7342
rect 288440 7278 288492 7284
rect 289820 6520 289872 6526
rect 289820 6462 289872 6468
rect 288440 6452 288492 6458
rect 288440 6394 288492 6400
rect 288452 3330 288480 6394
rect 288532 6384 288584 6390
rect 288532 6326 288584 6332
rect 288440 3324 288492 3330
rect 288440 3266 288492 3272
rect 288544 3262 288572 6326
rect 289544 3800 289596 3806
rect 289544 3742 289596 3748
rect 288532 3256 288584 3262
rect 288532 3198 288584 3204
rect 288268 598 288388 626
rect 288360 480 288388 598
rect 289556 480 289584 3742
rect 289832 3398 289860 6462
rect 289820 3392 289872 3398
rect 289820 3334 289872 3340
rect 290476 3194 290504 337826
rect 291212 7274 291240 340068
rect 291304 340054 291686 340082
rect 291304 9926 291332 340054
rect 291764 335594 291792 340190
rect 291580 335566 291792 335594
rect 292592 340054 292698 340082
rect 292868 340054 293158 340082
rect 293328 340054 293710 340082
rect 293972 340054 294170 340082
rect 294248 340054 294630 340082
rect 291580 317422 291608 335566
rect 291568 317416 291620 317422
rect 291568 317358 291620 317364
rect 291660 317348 291712 317354
rect 291660 317290 291712 317296
rect 291672 287094 291700 317290
rect 291568 287088 291620 287094
rect 291568 287030 291620 287036
rect 291660 287088 291712 287094
rect 291660 287030 291712 287036
rect 291580 278866 291608 287030
rect 291568 278860 291620 278866
rect 291568 278802 291620 278808
rect 291752 278860 291804 278866
rect 291752 278802 291804 278808
rect 291764 269210 291792 278802
rect 291752 269204 291804 269210
rect 291752 269146 291804 269152
rect 291568 269068 291620 269074
rect 291568 269010 291620 269016
rect 291580 258233 291608 269010
rect 291566 258224 291622 258233
rect 291566 258159 291622 258168
rect 291474 258088 291530 258097
rect 291474 258023 291530 258032
rect 291488 248441 291516 258023
rect 291474 248432 291530 248441
rect 291474 248367 291530 248376
rect 291842 248432 291898 248441
rect 291842 248367 291898 248376
rect 291856 230194 291884 248367
rect 291856 230166 291976 230194
rect 291948 220862 291976 230166
rect 291660 220856 291712 220862
rect 291660 220798 291712 220804
rect 291936 220856 291988 220862
rect 291936 220798 291988 220804
rect 291672 219434 291700 220798
rect 291660 219428 291712 219434
rect 291660 219370 291712 219376
rect 291660 212492 291712 212498
rect 291660 212434 291712 212440
rect 291672 209794 291700 212434
rect 291672 209766 291792 209794
rect 291764 203130 291792 209766
rect 291764 203102 291884 203130
rect 291856 201657 291884 203102
rect 291842 201648 291898 201657
rect 291842 201583 291898 201592
rect 291658 201512 291714 201521
rect 291658 201447 291714 201456
rect 291672 200122 291700 201447
rect 291384 200116 291436 200122
rect 291384 200058 291436 200064
rect 291660 200116 291712 200122
rect 291660 200058 291712 200064
rect 291396 190505 291424 200058
rect 291382 190496 291438 190505
rect 291382 190431 291438 190440
rect 291566 190496 291622 190505
rect 291566 190431 291622 190440
rect 291580 188578 291608 190431
rect 291488 188550 291608 188578
rect 291488 188306 291516 188550
rect 291488 188278 291608 188306
rect 291580 183546 291608 188278
rect 291488 183518 291608 183546
rect 291488 172689 291516 183518
rect 291474 172680 291530 172689
rect 291474 172615 291530 172624
rect 291474 172544 291530 172553
rect 291474 172479 291530 172488
rect 291488 164914 291516 172479
rect 291396 164886 291516 164914
rect 291396 161362 291424 164886
rect 291384 161356 291436 161362
rect 291384 161298 291436 161304
rect 291568 161356 291620 161362
rect 291568 161298 291620 161304
rect 291580 160070 291608 161298
rect 291568 160064 291620 160070
rect 291568 160006 291620 160012
rect 291476 149116 291528 149122
rect 291476 149058 291528 149064
rect 291488 139398 291516 149058
rect 291476 139392 291528 139398
rect 291476 139334 291528 139340
rect 291660 121508 291712 121514
rect 291660 121450 291712 121456
rect 291672 117994 291700 121450
rect 291580 117966 291700 117994
rect 291580 104922 291608 117966
rect 291568 104916 291620 104922
rect 291568 104858 291620 104864
rect 291660 104916 291712 104922
rect 291660 104858 291712 104864
rect 291672 93974 291700 104858
rect 291660 93968 291712 93974
rect 291660 93910 291712 93916
rect 291752 93900 291804 93906
rect 291752 93842 291804 93848
rect 291764 93786 291792 93842
rect 291672 93758 291792 93786
rect 291672 85610 291700 93758
rect 291660 85604 291712 85610
rect 291660 85546 291712 85552
rect 291568 84244 291620 84250
rect 291568 84186 291620 84192
rect 291580 75954 291608 84186
rect 291384 75948 291436 75954
rect 291384 75890 291436 75896
rect 291568 75948 291620 75954
rect 291568 75890 291620 75896
rect 291396 75834 291424 75890
rect 291396 75806 291516 75834
rect 291488 12170 291516 75806
rect 291476 12164 291528 12170
rect 291476 12106 291528 12112
rect 291292 9920 291344 9926
rect 291292 9862 291344 9868
rect 291200 7268 291252 7274
rect 291200 7210 291252 7216
rect 292592 7206 292620 340054
rect 292764 335640 292816 335646
rect 292764 335582 292816 335588
rect 292776 12238 292804 335582
rect 292764 12232 292816 12238
rect 292764 12174 292816 12180
rect 292868 9858 292896 340054
rect 293328 335646 293356 340054
rect 293316 335640 293368 335646
rect 293316 335582 293368 335588
rect 292856 9852 292908 9858
rect 292856 9794 292908 9800
rect 292580 7200 292632 7206
rect 292580 7142 292632 7148
rect 293972 7138 294000 340054
rect 294248 335696 294276 340054
rect 294064 335668 294276 335696
rect 294064 9790 294092 335668
rect 294708 331242 294736 340190
rect 294248 331214 294736 331242
rect 295352 340054 295642 340082
rect 295720 340054 296102 340082
rect 296272 340054 296654 340082
rect 296732 340054 297114 340082
rect 297284 340054 297574 340082
rect 298126 340054 298232 340082
rect 294248 318850 294276 331214
rect 294236 318844 294288 318850
rect 294236 318786 294288 318792
rect 294328 318844 294380 318850
rect 294328 318786 294380 318792
rect 294340 312610 294368 318786
rect 294340 312582 294552 312610
rect 294524 309108 294552 312582
rect 294432 309080 294552 309108
rect 294432 304298 294460 309080
rect 294236 304292 294288 304298
rect 294236 304234 294288 304240
rect 294420 304292 294472 304298
rect 294420 304234 294472 304240
rect 294248 296698 294276 304234
rect 294248 296670 294368 296698
rect 294340 289882 294368 296670
rect 294328 289876 294380 289882
rect 294328 289818 294380 289824
rect 294236 287088 294288 287094
rect 294236 287030 294288 287036
rect 294248 277438 294276 287030
rect 294236 277432 294288 277438
rect 294236 277374 294288 277380
rect 294328 277432 294380 277438
rect 294328 277374 294380 277380
rect 294340 267782 294368 277374
rect 294144 267776 294196 267782
rect 294142 267744 294144 267753
rect 294328 267776 294380 267782
rect 294196 267744 294198 267753
rect 294328 267718 294380 267724
rect 294142 267679 294198 267688
rect 294234 267608 294290 267617
rect 294234 267543 294290 267552
rect 294248 241482 294276 267543
rect 295248 253224 295300 253230
rect 295248 253166 295300 253172
rect 295260 248441 295288 253166
rect 295246 248432 295302 248441
rect 295246 248367 295302 248376
rect 294248 241454 294368 241482
rect 294340 240106 294368 241454
rect 294328 240100 294380 240106
rect 294328 240042 294380 240048
rect 294420 240100 294472 240106
rect 294420 240042 294472 240048
rect 294432 220862 294460 240042
rect 294328 220856 294380 220862
rect 294328 220798 294380 220804
rect 294420 220856 294472 220862
rect 294420 220798 294472 220804
rect 294340 211138 294368 220798
rect 294236 211132 294288 211138
rect 294236 211074 294288 211080
rect 294328 211132 294380 211138
rect 294328 211074 294380 211080
rect 294248 198082 294276 211074
rect 294236 198076 294288 198082
rect 294236 198018 294288 198024
rect 294420 198076 294472 198082
rect 294420 198018 294472 198024
rect 294432 183598 294460 198018
rect 294236 183592 294288 183598
rect 294236 183534 294288 183540
rect 294420 183592 294472 183598
rect 294420 183534 294472 183540
rect 294248 178770 294276 183534
rect 294236 178764 294288 178770
rect 294236 178706 294288 178712
rect 294420 178764 294472 178770
rect 294420 178706 294472 178712
rect 294432 171086 294460 178706
rect 294420 171080 294472 171086
rect 294420 171022 294472 171028
rect 294420 161492 294472 161498
rect 294420 161434 294472 161440
rect 294432 160070 294460 161434
rect 294420 160064 294472 160070
rect 294420 160006 294472 160012
rect 294512 150476 294564 150482
rect 294512 150418 294564 150424
rect 294524 150346 294552 150418
rect 294512 150340 294564 150346
rect 294512 150282 294564 150288
rect 294236 140820 294288 140826
rect 294236 140762 294288 140768
rect 294248 140706 294276 140762
rect 294248 140678 294368 140706
rect 294340 109698 294368 140678
rect 294248 109670 294368 109698
rect 294248 100094 294276 109670
rect 294236 100088 294288 100094
rect 294236 100030 294288 100036
rect 294420 100088 294472 100094
rect 294420 100030 294472 100036
rect 294432 85610 294460 100030
rect 294236 85604 294288 85610
rect 294236 85546 294288 85552
rect 294420 85604 294472 85610
rect 294420 85546 294472 85552
rect 294248 64870 294276 85546
rect 294236 64864 294288 64870
rect 294236 64806 294288 64812
rect 294236 55276 294288 55282
rect 294236 55218 294288 55224
rect 294248 45558 294276 55218
rect 294236 45552 294288 45558
rect 294236 45494 294288 45500
rect 294420 45552 294472 45558
rect 294420 45494 294472 45500
rect 294432 20754 294460 45494
rect 295246 29608 295302 29617
rect 295246 29543 295302 29552
rect 295260 29345 295288 29543
rect 295246 29336 295302 29345
rect 295246 29271 295302 29280
rect 294248 20726 294460 20754
rect 294248 13326 294276 20726
rect 294236 13320 294288 13326
rect 294236 13262 294288 13268
rect 294052 9784 294104 9790
rect 294052 9726 294104 9732
rect 293960 7132 294012 7138
rect 293960 7074 294012 7080
rect 295352 7070 295380 340054
rect 295720 335696 295748 340054
rect 295444 335668 295748 335696
rect 295444 9722 295472 335668
rect 296272 335594 296300 340054
rect 295536 335566 296300 335594
rect 295536 328438 295564 335566
rect 295524 328432 295576 328438
rect 295524 328374 295576 328380
rect 295708 328432 295760 328438
rect 295708 328374 295760 328380
rect 295720 323490 295748 328374
rect 295628 323462 295748 323490
rect 295628 309262 295656 323462
rect 295616 309256 295668 309262
rect 295616 309198 295668 309204
rect 295524 309120 295576 309126
rect 295524 309062 295576 309068
rect 295536 292602 295564 309062
rect 295524 292596 295576 292602
rect 295524 292538 295576 292544
rect 295616 292528 295668 292534
rect 295616 292470 295668 292476
rect 295628 280226 295656 292470
rect 295524 280220 295576 280226
rect 295524 280162 295576 280168
rect 295616 280220 295668 280226
rect 295616 280162 295668 280168
rect 295536 267782 295564 280162
rect 295524 267776 295576 267782
rect 295800 267776 295852 267782
rect 295524 267718 295576 267724
rect 295720 267724 295800 267730
rect 295720 267718 295852 267724
rect 295720 267702 295840 267718
rect 295720 260914 295748 267702
rect 295708 260908 295760 260914
rect 295708 260850 295760 260856
rect 295800 260840 295852 260846
rect 295800 260782 295852 260788
rect 295812 258097 295840 260782
rect 295614 258088 295670 258097
rect 295614 258023 295670 258032
rect 295798 258088 295854 258097
rect 295798 258023 295854 258032
rect 295628 253230 295656 258023
rect 295616 253224 295668 253230
rect 295616 253166 295668 253172
rect 295522 248432 295578 248441
rect 295522 248367 295524 248376
rect 295576 248367 295578 248376
rect 295800 248396 295852 248402
rect 295524 248338 295576 248344
rect 295800 248338 295852 248344
rect 295812 238785 295840 248338
rect 295614 238776 295670 238785
rect 295614 238711 295616 238720
rect 295668 238711 295670 238720
rect 295798 238776 295854 238785
rect 295798 238711 295854 238720
rect 295616 238682 295668 238688
rect 295616 229152 295668 229158
rect 295616 229094 295668 229100
rect 295536 222222 295564 222253
rect 295628 222222 295656 229094
rect 295524 222216 295576 222222
rect 295616 222216 295668 222222
rect 295576 222164 295616 222170
rect 295524 222158 295668 222164
rect 295536 222142 295656 222158
rect 295536 202910 295564 202941
rect 295628 202910 295656 222142
rect 295524 202904 295576 202910
rect 295616 202904 295668 202910
rect 295576 202852 295616 202858
rect 295524 202846 295668 202852
rect 295536 202830 295656 202846
rect 295628 186386 295656 202830
rect 295616 186380 295668 186386
rect 295616 186322 295668 186328
rect 295524 186312 295576 186318
rect 295524 186254 295576 186260
rect 295536 178770 295564 186254
rect 295524 178764 295576 178770
rect 295524 178706 295576 178712
rect 295708 178764 295760 178770
rect 295708 178706 295760 178712
rect 295720 164218 295748 178706
rect 295524 164212 295576 164218
rect 295524 164154 295576 164160
rect 295708 164212 295760 164218
rect 295708 164154 295760 164160
rect 295536 132530 295564 164154
rect 295524 132524 295576 132530
rect 295524 132466 295576 132472
rect 295616 132524 295668 132530
rect 295616 132466 295668 132472
rect 295628 127650 295656 132466
rect 295628 127622 295840 127650
rect 295812 121446 295840 127622
rect 295800 121440 295852 121446
rect 295800 121382 295852 121388
rect 295524 111852 295576 111858
rect 295524 111794 295576 111800
rect 295536 101998 295564 111794
rect 295524 101992 295576 101998
rect 295524 101934 295576 101940
rect 295708 92540 295760 92546
rect 295708 92482 295760 92488
rect 295720 87038 295748 92482
rect 295708 87032 295760 87038
rect 295708 86974 295760 86980
rect 295708 86896 295760 86902
rect 295708 86838 295760 86844
rect 295720 75954 295748 86838
rect 295524 75948 295576 75954
rect 295524 75890 295576 75896
rect 295708 75948 295760 75954
rect 295708 75890 295760 75896
rect 295536 57050 295564 75890
rect 296626 64016 296682 64025
rect 296626 63951 296682 63960
rect 296640 63617 296668 63951
rect 296626 63608 296682 63617
rect 296626 63543 296682 63552
rect 295524 57044 295576 57050
rect 295524 56986 295576 56992
rect 295524 48340 295576 48346
rect 295524 48282 295576 48288
rect 295536 38690 295564 48282
rect 295524 38684 295576 38690
rect 295524 38626 295576 38632
rect 295616 38548 295668 38554
rect 295616 38490 295668 38496
rect 295628 29034 295656 38490
rect 296626 29472 296682 29481
rect 296626 29407 296682 29416
rect 296640 29345 296668 29407
rect 296626 29336 296682 29345
rect 296626 29271 296682 29280
rect 295524 29028 295576 29034
rect 295524 28970 295576 28976
rect 295616 29028 295668 29034
rect 295616 28970 295668 28976
rect 295536 27606 295564 28970
rect 295524 27600 295576 27606
rect 295524 27542 295576 27548
rect 295432 9716 295484 9722
rect 295432 9658 295484 9664
rect 295340 7064 295392 7070
rect 295340 7006 295392 7012
rect 296732 6730 296760 340054
rect 297284 335696 297312 340054
rect 297916 337204 297968 337210
rect 297916 337146 297968 337152
rect 296824 335668 297312 335696
rect 296824 328438 296852 335668
rect 296812 328432 296864 328438
rect 296812 328374 296864 328380
rect 296996 328432 297048 328438
rect 296996 328374 297048 328380
rect 297008 323490 297036 328374
rect 296916 323462 297036 323490
rect 296916 309262 296944 323462
rect 296904 309256 296956 309262
rect 296904 309198 296956 309204
rect 296812 309120 296864 309126
rect 296812 309062 296864 309068
rect 296824 292602 296852 309062
rect 296812 292596 296864 292602
rect 296812 292538 296864 292544
rect 296904 292528 296956 292534
rect 296904 292470 296956 292476
rect 296916 283014 296944 292470
rect 296904 283008 296956 283014
rect 296904 282950 296956 282956
rect 296812 282872 296864 282878
rect 296812 282814 296864 282820
rect 296824 269142 296852 282814
rect 296812 269136 296864 269142
rect 296812 269078 296864 269084
rect 297088 269136 297140 269142
rect 297088 269078 297140 269084
rect 297100 267730 297128 269078
rect 297008 267702 297128 267730
rect 297008 262954 297036 267702
rect 296812 262948 296864 262954
rect 296812 262890 296864 262896
rect 296996 262948 297048 262954
rect 296996 262890 297048 262896
rect 296824 258097 296852 262890
rect 296810 258088 296866 258097
rect 296810 258023 296866 258032
rect 296994 258088 297050 258097
rect 296994 258023 297050 258032
rect 297008 248470 297036 258023
rect 296904 248464 296956 248470
rect 296824 248412 296904 248418
rect 296824 248406 296956 248412
rect 296996 248464 297048 248470
rect 296996 248406 297048 248412
rect 296824 248390 296944 248406
rect 296824 239850 296852 248390
rect 296824 239822 296944 239850
rect 296824 202910 296852 202941
rect 296916 202910 296944 239822
rect 296812 202904 296864 202910
rect 296904 202904 296956 202910
rect 296864 202852 296904 202858
rect 296812 202846 296956 202852
rect 296824 202830 296944 202846
rect 296916 186454 296944 202830
rect 296904 186448 296956 186454
rect 296904 186390 296956 186396
rect 296812 186312 296864 186318
rect 296812 186254 296864 186260
rect 296824 178770 296852 186254
rect 296812 178764 296864 178770
rect 296812 178706 296864 178712
rect 296996 178764 297048 178770
rect 296996 178706 297048 178712
rect 297008 161498 297036 178706
rect 296996 161492 297048 161498
rect 296996 161434 297048 161440
rect 297088 161492 297140 161498
rect 297088 161434 297140 161440
rect 297100 151842 297128 161434
rect 296904 151836 296956 151842
rect 296904 151778 296956 151784
rect 297088 151836 297140 151842
rect 297088 151778 297140 151784
rect 296916 151745 296944 151778
rect 296902 151736 296958 151745
rect 296902 151671 296958 151680
rect 297178 151736 297234 151745
rect 297178 151671 297234 151680
rect 297192 142361 297220 151671
rect 297178 142352 297234 142361
rect 297178 142287 297234 142296
rect 296810 142216 296866 142225
rect 296810 142151 296866 142160
rect 296824 142118 296852 142151
rect 296812 142112 296864 142118
rect 296812 142054 296864 142060
rect 296904 132524 296956 132530
rect 296904 132466 296956 132472
rect 296916 122738 296944 132466
rect 296904 122732 296956 122738
rect 296904 122674 296956 122680
rect 296904 113212 296956 113218
rect 296904 113154 296956 113160
rect 296916 104922 296944 113154
rect 296812 104916 296864 104922
rect 296812 104858 296864 104864
rect 296904 104916 296956 104922
rect 296904 104858 296956 104864
rect 296824 95266 296852 104858
rect 296812 95260 296864 95266
rect 296812 95202 296864 95208
rect 296996 95124 297048 95130
rect 296996 95066 297048 95072
rect 297008 75954 297036 95066
rect 296812 75948 296864 75954
rect 296812 75890 296864 75896
rect 296996 75948 297048 75954
rect 296996 75890 297048 75896
rect 296824 66230 296852 75890
rect 296812 66224 296864 66230
rect 296812 66166 296864 66172
rect 296812 56228 296864 56234
rect 296812 56170 296864 56176
rect 296824 46850 296852 56170
rect 296812 46844 296864 46850
rect 296812 46786 296864 46792
rect 296904 43988 296956 43994
rect 296904 43930 296956 43936
rect 296916 13394 296944 43930
rect 296904 13388 296956 13394
rect 296904 13330 296956 13336
rect 296720 6724 296772 6730
rect 296720 6666 296772 6672
rect 297364 6724 297416 6730
rect 297364 6666 297416 6672
rect 295892 6656 295944 6662
rect 295892 6598 295944 6604
rect 294328 6316 294380 6322
rect 294328 6258 294380 6264
rect 290740 5432 290792 5438
rect 290740 5374 290792 5380
rect 290464 3188 290516 3194
rect 290464 3130 290516 3136
rect 290752 480 290780 5374
rect 291936 3256 291988 3262
rect 291936 3198 291988 3204
rect 291948 480 291976 3198
rect 293132 3052 293184 3058
rect 293132 2994 293184 3000
rect 293144 480 293172 2994
rect 294340 480 294368 6258
rect 295904 4146 295932 6598
rect 295892 4140 295944 4146
rect 295892 4082 295944 4088
rect 296720 4140 296772 4146
rect 296720 4082 296772 4088
rect 295524 3188 295576 3194
rect 295524 3130 295576 3136
rect 295536 480 295564 3130
rect 296732 480 296760 4082
rect 297376 4010 297404 6666
rect 297824 5500 297876 5506
rect 297824 5442 297876 5448
rect 297836 4026 297864 5442
rect 297928 4146 297956 337146
rect 298006 16824 298062 16833
rect 298006 16759 298062 16768
rect 298020 16561 298048 16759
rect 298006 16552 298062 16561
rect 298006 16487 298062 16496
rect 298204 12374 298232 340054
rect 298388 340054 298586 340082
rect 298664 340054 299046 340082
rect 298284 335640 298336 335646
rect 298284 335582 298336 335588
rect 298296 13462 298324 335582
rect 298284 13456 298336 13462
rect 298284 13398 298336 13404
rect 298192 12368 298244 12374
rect 298192 12310 298244 12316
rect 298388 6798 298416 340054
rect 298664 335646 298692 340054
rect 298652 335640 298704 335646
rect 298652 335582 298704 335588
rect 299584 331362 299612 340068
rect 299768 340054 300058 340082
rect 299768 331378 299796 340054
rect 300136 339130 300164 340190
rect 300044 339102 300164 339130
rect 300964 340054 301070 340082
rect 301240 340054 301530 340082
rect 301700 340054 301990 340082
rect 302344 340054 302542 340082
rect 302712 340054 303002 340082
rect 303080 340054 303462 340082
rect 303724 340054 303922 340082
rect 304184 340054 304474 340082
rect 304644 340054 304934 340082
rect 305104 340054 305394 340082
rect 305656 340054 305946 340082
rect 299572 331356 299624 331362
rect 299768 331350 299888 331378
rect 299572 331298 299624 331304
rect 299572 331084 299624 331090
rect 299572 331026 299624 331032
rect 299480 331016 299532 331022
rect 299480 330958 299532 330964
rect 299492 241466 299520 330958
rect 299480 241460 299532 241466
rect 299480 241402 299532 241408
rect 299480 231872 299532 231878
rect 299480 231814 299532 231820
rect 299492 222154 299520 231814
rect 299480 222148 299532 222154
rect 299480 222090 299532 222096
rect 299480 212560 299532 212566
rect 299480 212502 299532 212508
rect 299492 6866 299520 212502
rect 299584 12442 299612 331026
rect 299860 331022 299888 331350
rect 299848 331016 299900 331022
rect 299848 330958 299900 330964
rect 300044 330698 300072 339102
rect 300860 335640 300912 335646
rect 300860 335582 300912 335588
rect 299860 330670 300072 330698
rect 299860 317422 299888 330670
rect 299848 317416 299900 317422
rect 299848 317358 299900 317364
rect 299848 299532 299900 299538
rect 299848 299474 299900 299480
rect 299860 296682 299888 299474
rect 299848 296676 299900 296682
rect 299848 296618 299900 296624
rect 299940 296676 299992 296682
rect 299940 296618 299992 296624
rect 299952 270638 299980 296618
rect 299940 270632 299992 270638
rect 299940 270574 299992 270580
rect 299756 270564 299808 270570
rect 299756 270506 299808 270512
rect 299768 260658 299796 270506
rect 299768 260630 299888 260658
rect 299860 259434 299888 260630
rect 299768 259406 299888 259434
rect 299768 254538 299796 259406
rect 299768 254510 299888 254538
rect 299860 249801 299888 254510
rect 299846 249792 299902 249801
rect 299846 249727 299902 249736
rect 299938 249656 299994 249665
rect 299938 249591 299994 249600
rect 299952 231860 299980 249591
rect 299860 231832 299980 231860
rect 299860 222306 299888 231832
rect 299860 222278 299980 222306
rect 299952 211206 299980 222278
rect 299848 211200 299900 211206
rect 299848 211142 299900 211148
rect 299940 211200 299992 211206
rect 299940 211142 299992 211148
rect 299860 200297 299888 211142
rect 299846 200288 299902 200297
rect 299846 200223 299902 200232
rect 299754 200152 299810 200161
rect 299754 200087 299756 200096
rect 299808 200087 299810 200096
rect 299848 200116 299900 200122
rect 299756 200058 299808 200064
rect 299848 200058 299900 200064
rect 299860 190466 299888 200058
rect 299848 190460 299900 190466
rect 299848 190402 299900 190408
rect 299848 180872 299900 180878
rect 299848 180814 299900 180820
rect 299860 156618 299888 180814
rect 299860 156590 299980 156618
rect 299952 137426 299980 156590
rect 299756 137420 299808 137426
rect 299756 137362 299808 137368
rect 299940 137420 299992 137426
rect 299940 137362 299992 137368
rect 299768 125610 299796 137362
rect 299768 125582 299888 125610
rect 299860 114594 299888 125582
rect 299768 114566 299888 114594
rect 299768 109834 299796 114566
rect 299768 109806 299888 109834
rect 299860 77314 299888 109806
rect 299756 77308 299808 77314
rect 299756 77250 299808 77256
rect 299848 77308 299900 77314
rect 299848 77250 299900 77256
rect 299768 47002 299796 77250
rect 299768 46974 300072 47002
rect 300044 37398 300072 46974
rect 300032 37392 300084 37398
rect 300032 37334 300084 37340
rect 299848 18012 299900 18018
rect 299848 17954 299900 17960
rect 299860 13530 299888 17954
rect 299848 13524 299900 13530
rect 299848 13466 299900 13472
rect 299572 12436 299624 12442
rect 299572 12378 299624 12384
rect 299480 6860 299532 6866
rect 299480 6802 299532 6808
rect 298376 6792 298428 6798
rect 298376 6734 298428 6740
rect 298100 6588 298152 6594
rect 298100 6530 298152 6536
rect 297916 4140 297968 4146
rect 297916 4082 297968 4088
rect 298112 4078 298140 6530
rect 300872 6118 300900 335582
rect 300964 124166 300992 340054
rect 301240 335646 301268 340054
rect 301228 335640 301280 335646
rect 301228 335582 301280 335588
rect 301700 333334 301728 340054
rect 302240 335708 302292 335714
rect 302240 335650 302292 335656
rect 301044 333328 301096 333334
rect 301044 333270 301096 333276
rect 301688 333328 301740 333334
rect 301688 333270 301740 333276
rect 301056 306406 301084 333270
rect 301044 306400 301096 306406
rect 301228 306400 301280 306406
rect 301044 306342 301096 306348
rect 301226 306368 301228 306377
rect 301280 306368 301282 306377
rect 301226 306303 301282 306312
rect 301410 306368 301466 306377
rect 301410 306303 301466 306312
rect 301424 296818 301452 306303
rect 301044 296812 301096 296818
rect 301044 296754 301096 296760
rect 301412 296812 301464 296818
rect 301412 296754 301464 296760
rect 301056 296682 301084 296754
rect 301044 296676 301096 296682
rect 301044 296618 301096 296624
rect 301136 296676 301188 296682
rect 301136 296618 301188 296624
rect 301148 283778 301176 296618
rect 301148 283750 301268 283778
rect 301240 278798 301268 283750
rect 301044 278792 301096 278798
rect 301044 278734 301096 278740
rect 301228 278792 301280 278798
rect 301228 278734 301280 278740
rect 301056 273290 301084 278734
rect 301044 273284 301096 273290
rect 301044 273226 301096 273232
rect 301136 273216 301188 273222
rect 301136 273158 301188 273164
rect 301148 269090 301176 273158
rect 301148 269062 301268 269090
rect 301240 258058 301268 269062
rect 301228 258052 301280 258058
rect 301228 257994 301280 258000
rect 301412 258052 301464 258058
rect 301412 257994 301464 258000
rect 301424 248418 301452 257994
rect 301332 248390 301452 248418
rect 301332 240242 301360 248390
rect 301320 240236 301372 240242
rect 301320 240178 301372 240184
rect 301044 240100 301096 240106
rect 301044 240042 301096 240048
rect 301056 230518 301084 240042
rect 301044 230512 301096 230518
rect 301044 230454 301096 230460
rect 301228 230512 301280 230518
rect 301228 230454 301280 230460
rect 301240 222290 301268 230454
rect 301228 222284 301280 222290
rect 301228 222226 301280 222232
rect 301044 222148 301096 222154
rect 301044 222090 301096 222096
rect 301056 201482 301084 222090
rect 301044 201476 301096 201482
rect 301044 201418 301096 201424
rect 301136 201408 301188 201414
rect 301136 201350 301188 201356
rect 301148 188306 301176 201350
rect 301056 188278 301176 188306
rect 301056 182170 301084 188278
rect 301044 182164 301096 182170
rect 301044 182106 301096 182112
rect 301228 182164 301280 182170
rect 301228 182106 301280 182112
rect 301240 177154 301268 182106
rect 301148 177126 301268 177154
rect 301148 172514 301176 177126
rect 301044 172508 301096 172514
rect 301044 172450 301096 172456
rect 301136 172508 301188 172514
rect 301136 172450 301188 172456
rect 301056 156618 301084 172450
rect 301056 156590 301268 156618
rect 301240 154442 301268 156590
rect 301148 154414 301268 154442
rect 301148 144922 301176 154414
rect 301148 144894 301360 144922
rect 301332 143562 301360 144894
rect 301240 143534 301360 143562
rect 301240 142118 301268 143534
rect 301228 142112 301280 142118
rect 301228 142054 301280 142060
rect 301136 132524 301188 132530
rect 301136 132466 301188 132472
rect 300952 124160 301004 124166
rect 300952 124102 301004 124108
rect 300952 124024 301004 124030
rect 300952 123966 301004 123972
rect 300964 11694 300992 123966
rect 301148 122806 301176 132466
rect 301136 122800 301188 122806
rect 301136 122742 301188 122748
rect 301136 114436 301188 114442
rect 301136 114378 301188 114384
rect 301148 104854 301176 114378
rect 301136 104848 301188 104854
rect 301136 104790 301188 104796
rect 301320 104848 301372 104854
rect 301320 104790 301372 104796
rect 301332 96506 301360 104790
rect 301148 96478 301360 96506
rect 301148 93838 301176 96478
rect 301136 93832 301188 93838
rect 301136 93774 301188 93780
rect 301228 86896 301280 86902
rect 301228 86838 301280 86844
rect 301240 82822 301268 86838
rect 301228 82816 301280 82822
rect 301228 82758 301280 82764
rect 301228 73228 301280 73234
rect 301228 73170 301280 73176
rect 301240 69698 301268 73170
rect 301228 69692 301280 69698
rect 301228 69634 301280 69640
rect 301228 55140 301280 55146
rect 301228 55082 301280 55088
rect 301240 41970 301268 55082
rect 301240 41942 301360 41970
rect 301332 29102 301360 41942
rect 301320 29096 301372 29102
rect 301320 29038 301372 29044
rect 301228 28960 301280 28966
rect 301228 28902 301280 28908
rect 301240 27538 301268 28902
rect 301228 27532 301280 27538
rect 301228 27474 301280 27480
rect 301136 18012 301188 18018
rect 301136 17954 301188 17960
rect 301148 13598 301176 17954
rect 301136 13592 301188 13598
rect 301136 13534 301188 13540
rect 300952 11688 301004 11694
rect 300952 11630 301004 11636
rect 300860 6112 300912 6118
rect 300860 6054 300912 6060
rect 302252 6050 302280 335650
rect 302344 11626 302372 340054
rect 302712 335714 302740 340054
rect 302700 335708 302752 335714
rect 302700 335650 302752 335656
rect 303080 334762 303108 340054
rect 303160 337952 303212 337958
rect 303160 337894 303212 337900
rect 303068 334756 303120 334762
rect 303068 334698 303120 334704
rect 303172 334642 303200 337894
rect 303620 335640 303672 335646
rect 303620 335582 303672 335588
rect 302896 334614 303200 334642
rect 302516 328500 302568 328506
rect 302516 328442 302568 328448
rect 302528 327078 302556 328442
rect 302516 327072 302568 327078
rect 302516 327014 302568 327020
rect 302608 327072 302660 327078
rect 302608 327014 302660 327020
rect 302620 317506 302648 327014
rect 302528 317478 302648 317506
rect 302528 311250 302556 317478
rect 302528 311222 302740 311250
rect 302712 301594 302740 311222
rect 302528 301566 302740 301594
rect 302528 299418 302556 301566
rect 302528 299390 302648 299418
rect 302620 296698 302648 299390
rect 302528 296670 302648 296698
rect 302528 295322 302556 296670
rect 302516 295316 302568 295322
rect 302516 295258 302568 295264
rect 302700 295316 302752 295322
rect 302700 295258 302752 295264
rect 302712 285705 302740 295258
rect 302514 285696 302570 285705
rect 302514 285631 302570 285640
rect 302698 285696 302754 285705
rect 302698 285631 302754 285640
rect 302528 278798 302556 285631
rect 302516 278792 302568 278798
rect 302516 278734 302568 278740
rect 302608 278724 302660 278730
rect 302608 278666 302660 278672
rect 302620 276010 302648 278666
rect 302608 276004 302660 276010
rect 302608 275946 302660 275952
rect 302792 276004 302844 276010
rect 302792 275946 302844 275952
rect 302804 266393 302832 275946
rect 302514 266384 302570 266393
rect 302514 266319 302570 266328
rect 302790 266384 302846 266393
rect 302790 266319 302846 266328
rect 302528 258097 302556 266319
rect 302514 258088 302570 258097
rect 302514 258023 302570 258032
rect 302790 258088 302846 258097
rect 302790 258023 302846 258032
rect 302804 249830 302832 258023
rect 302700 249824 302752 249830
rect 302700 249766 302752 249772
rect 302792 249824 302844 249830
rect 302792 249766 302844 249772
rect 302712 231860 302740 249766
rect 302528 231832 302740 231860
rect 302528 222222 302556 231832
rect 302516 222216 302568 222222
rect 302516 222158 302568 222164
rect 302700 222216 302752 222222
rect 302700 222158 302752 222164
rect 302712 212650 302740 222158
rect 302712 212622 302832 212650
rect 302804 212378 302832 212622
rect 302620 212350 302832 212378
rect 302620 207806 302648 212350
rect 302608 207800 302660 207806
rect 302608 207742 302660 207748
rect 302608 202904 302660 202910
rect 302608 202846 302660 202852
rect 302620 196602 302648 202846
rect 302620 196574 302832 196602
rect 302804 190466 302832 196574
rect 302792 190460 302844 190466
rect 302792 190402 302844 190408
rect 302516 180872 302568 180878
rect 302516 180814 302568 180820
rect 302528 161498 302556 180814
rect 302516 161492 302568 161498
rect 302516 161434 302568 161440
rect 302608 161492 302660 161498
rect 302608 161434 302660 161440
rect 302620 154562 302648 161434
rect 302516 154556 302568 154562
rect 302516 154498 302568 154504
rect 302608 154556 302660 154562
rect 302608 154498 302660 154504
rect 302528 153202 302556 154498
rect 302424 153196 302476 153202
rect 302424 153138 302476 153144
rect 302516 153196 302568 153202
rect 302516 153138 302568 153144
rect 302436 143585 302464 153138
rect 302422 143576 302478 143585
rect 302422 143511 302478 143520
rect 302606 143576 302662 143585
rect 302606 143511 302662 143520
rect 302620 135250 302648 143511
rect 302516 135244 302568 135250
rect 302516 135186 302568 135192
rect 302608 135244 302660 135250
rect 302608 135186 302660 135192
rect 302528 133890 302556 135186
rect 302516 133884 302568 133890
rect 302516 133826 302568 133832
rect 302608 124228 302660 124234
rect 302608 124170 302660 124176
rect 302620 113218 302648 124170
rect 302424 113212 302476 113218
rect 302424 113154 302476 113160
rect 302608 113212 302660 113218
rect 302608 113154 302660 113160
rect 302436 104922 302464 113154
rect 302424 104916 302476 104922
rect 302424 104858 302476 104864
rect 302516 104916 302568 104922
rect 302516 104858 302568 104864
rect 302528 96694 302556 104858
rect 302516 96688 302568 96694
rect 302516 96630 302568 96636
rect 302608 96552 302660 96558
rect 302608 96494 302660 96500
rect 302620 82822 302648 96494
rect 302608 82816 302660 82822
rect 302608 82758 302660 82764
rect 302700 73228 302752 73234
rect 302700 73170 302752 73176
rect 302712 59566 302740 73170
rect 302700 59560 302752 59566
rect 302700 59502 302752 59508
rect 302516 46980 302568 46986
rect 302516 46922 302568 46928
rect 302528 42106 302556 46922
rect 302528 42078 302648 42106
rect 302620 19378 302648 42078
rect 302516 19372 302568 19378
rect 302516 19314 302568 19320
rect 302608 19372 302660 19378
rect 302608 19314 302660 19320
rect 302528 13666 302556 19314
rect 302516 13660 302568 13666
rect 302516 13602 302568 13608
rect 302332 11620 302384 11626
rect 302332 11562 302384 11568
rect 302240 6044 302292 6050
rect 302240 5986 302292 5992
rect 301412 4412 301464 4418
rect 301412 4354 301464 4360
rect 300308 4140 300360 4146
rect 300308 4082 300360 4088
rect 298100 4072 298152 4078
rect 297364 4004 297416 4010
rect 297836 3998 297956 4026
rect 298100 4014 298152 4020
rect 297364 3946 297416 3952
rect 297928 480 297956 3998
rect 299112 3392 299164 3398
rect 299112 3334 299164 3340
rect 299124 480 299152 3334
rect 300320 480 300348 4082
rect 301424 480 301452 4354
rect 302608 4072 302660 4078
rect 302608 4014 302660 4020
rect 302620 480 302648 4014
rect 302896 3398 302924 334614
rect 303632 5982 303660 335582
rect 303724 11558 303752 340054
rect 304184 335646 304212 340054
rect 304172 335640 304224 335646
rect 304172 335582 304224 335588
rect 304644 328506 304672 340054
rect 305000 333804 305052 333810
rect 305000 333746 305052 333752
rect 303896 328500 303948 328506
rect 303896 328442 303948 328448
rect 304632 328500 304684 328506
rect 304632 328442 304684 328448
rect 303908 311930 303936 328442
rect 303816 311902 303936 311930
rect 303816 311794 303844 311902
rect 303816 311766 303936 311794
rect 303908 292618 303936 311766
rect 303816 292590 303936 292618
rect 303816 292482 303844 292590
rect 303816 292454 303936 292482
rect 303908 196058 303936 292454
rect 303816 196030 303936 196058
rect 303816 195922 303844 196030
rect 303816 195894 303936 195922
rect 303908 176746 303936 195894
rect 303816 176718 303936 176746
rect 303816 176610 303844 176718
rect 303816 176582 303936 176610
rect 303908 138122 303936 176582
rect 303816 138094 303936 138122
rect 303816 137714 303844 138094
rect 303816 137686 303936 137714
rect 303908 118810 303936 137686
rect 303816 118782 303936 118810
rect 303816 118674 303844 118782
rect 303816 118646 303936 118674
rect 303908 80102 303936 118646
rect 304262 87408 304318 87417
rect 304262 87343 304318 87352
rect 304276 87009 304304 87343
rect 304262 87000 304318 87009
rect 304262 86935 304318 86944
rect 303896 80096 303948 80102
rect 303896 80038 303948 80044
rect 303896 79960 303948 79966
rect 303896 79902 303948 79908
rect 303908 77246 303936 79902
rect 303896 77240 303948 77246
rect 303896 77182 303948 77188
rect 303988 77240 304040 77246
rect 303988 77182 304040 77188
rect 304000 61418 304028 77182
rect 303908 61390 304028 61418
rect 303908 48414 303936 61390
rect 303896 48408 303948 48414
rect 303896 48350 303948 48356
rect 303896 48272 303948 48278
rect 303896 48214 303948 48220
rect 303908 42090 303936 48214
rect 303896 42084 303948 42090
rect 303896 42026 303948 42032
rect 303896 32428 303948 32434
rect 303896 32370 303948 32376
rect 303908 13734 303936 32370
rect 303896 13728 303948 13734
rect 303896 13670 303948 13676
rect 303712 11552 303764 11558
rect 303712 11494 303764 11500
rect 303620 5976 303672 5982
rect 303620 5918 303672 5924
rect 305012 5914 305040 333746
rect 305104 11490 305132 340054
rect 305656 333810 305684 340054
rect 306196 338020 306248 338026
rect 306196 337962 306248 337968
rect 305644 333804 305696 333810
rect 305644 333746 305696 333752
rect 305092 11484 305144 11490
rect 305092 11426 305144 11432
rect 305000 5908 305052 5914
rect 305000 5850 305052 5856
rect 305000 4344 305052 4350
rect 305000 4286 305052 4292
rect 302884 3392 302936 3398
rect 302884 3334 302936 3340
rect 303804 3324 303856 3330
rect 303804 3266 303856 3272
rect 303816 480 303844 3266
rect 305012 480 305040 4286
rect 306208 480 306236 337962
rect 306392 333282 306420 340068
rect 306668 340054 306866 340082
rect 307036 340054 307418 340082
rect 307878 340054 307984 340082
rect 306392 333254 306604 333282
rect 306472 333124 306524 333130
rect 306472 333066 306524 333072
rect 306288 157480 306340 157486
rect 306286 157448 306288 157457
rect 306340 157448 306342 157457
rect 306286 157383 306342 157392
rect 306286 110800 306342 110809
rect 306286 110735 306342 110744
rect 306300 110537 306328 110735
rect 306286 110528 306342 110537
rect 306286 110463 306342 110472
rect 306286 29200 306342 29209
rect 306286 29135 306342 29144
rect 306300 28937 306328 29135
rect 306286 28928 306342 28937
rect 306286 28863 306342 28872
rect 306484 11422 306512 333066
rect 306576 13802 306604 333254
rect 306668 333130 306696 340054
rect 306656 333124 306708 333130
rect 306656 333066 306708 333072
rect 307036 331242 307064 340054
rect 307760 335640 307812 335646
rect 307760 335582 307812 335588
rect 306760 331214 307064 331242
rect 306760 318850 306788 331214
rect 306748 318844 306800 318850
rect 306748 318786 306800 318792
rect 306840 318844 306892 318850
rect 306840 318786 306892 318792
rect 306852 311982 306880 318786
rect 306840 311976 306892 311982
rect 306840 311918 306892 311924
rect 306748 311840 306800 311846
rect 306748 311782 306800 311788
rect 306760 299538 306788 311782
rect 306748 299532 306800 299538
rect 306748 299474 306800 299480
rect 306840 299532 306892 299538
rect 306840 299474 306892 299480
rect 306852 296682 306880 299474
rect 306840 296676 306892 296682
rect 306840 296618 306892 296624
rect 306932 296676 306984 296682
rect 306932 296618 306984 296624
rect 306944 276010 306972 296618
rect 306656 276004 306708 276010
rect 306656 275946 306708 275952
rect 306932 276004 306984 276010
rect 306932 275946 306984 275952
rect 306668 266393 306696 275946
rect 306654 266384 306710 266393
rect 306654 266319 306710 266328
rect 306838 266384 306894 266393
rect 306838 266319 306894 266328
rect 306852 258058 306880 266319
rect 306840 258052 306892 258058
rect 306840 257994 306892 258000
rect 306748 248396 306800 248402
rect 306748 248338 306800 248344
rect 306760 238814 306788 248338
rect 306748 238808 306800 238814
rect 306748 238750 306800 238756
rect 306840 230512 306892 230518
rect 306840 230454 306892 230460
rect 306852 222306 306880 230454
rect 306852 222278 306972 222306
rect 306944 212548 306972 222278
rect 306852 212520 306972 212548
rect 306852 211138 306880 212520
rect 306656 211132 306708 211138
rect 306656 211074 306708 211080
rect 306840 211132 306892 211138
rect 306840 211074 306892 211080
rect 306668 209778 306696 211074
rect 306656 209772 306708 209778
rect 306656 209714 306708 209720
rect 306932 209772 306984 209778
rect 306932 209714 306984 209720
rect 306944 200161 306972 209714
rect 306746 200152 306802 200161
rect 306930 200152 306986 200161
rect 306746 200087 306748 200096
rect 306800 200087 306802 200096
rect 306840 200116 306892 200122
rect 306748 200058 306800 200064
rect 306930 200087 306986 200096
rect 306840 200058 306892 200064
rect 306852 190466 306880 200058
rect 306840 190460 306892 190466
rect 306840 190402 306892 190408
rect 306840 180872 306892 180878
rect 306840 180814 306892 180820
rect 306852 171086 306880 180814
rect 306840 171080 306892 171086
rect 306840 171022 306892 171028
rect 307024 171080 307076 171086
rect 307024 171022 307076 171028
rect 307036 161537 307064 171022
rect 306838 161528 306894 161537
rect 306838 161463 306894 161472
rect 307022 161528 307078 161537
rect 307022 161463 307078 161472
rect 306852 161430 306880 161463
rect 306840 161424 306892 161430
rect 306840 161366 306892 161372
rect 306932 151836 306984 151842
rect 306932 151778 306984 151784
rect 306944 137426 306972 151778
rect 306748 137420 306800 137426
rect 306748 137362 306800 137368
rect 306932 137420 306984 137426
rect 306932 137362 306984 137368
rect 306760 133890 306788 137362
rect 306748 133884 306800 133890
rect 306748 133826 306800 133832
rect 306840 124228 306892 124234
rect 306840 124170 306892 124176
rect 306852 122806 306880 124170
rect 306840 122800 306892 122806
rect 306840 122742 306892 122748
rect 306656 113212 306708 113218
rect 306656 113154 306708 113160
rect 306668 104922 306696 113154
rect 307666 110800 307722 110809
rect 307666 110735 307722 110744
rect 307680 110634 307708 110735
rect 307668 110628 307720 110634
rect 307668 110570 307720 110576
rect 306656 104916 306708 104922
rect 306656 104858 306708 104864
rect 306840 104916 306892 104922
rect 306840 104858 306892 104864
rect 306852 98734 306880 104858
rect 306840 98728 306892 98734
rect 306840 98670 306892 98676
rect 307024 98728 307076 98734
rect 307024 98670 307076 98676
rect 307036 93945 307064 98670
rect 306838 93936 306894 93945
rect 306760 93894 306838 93922
rect 306760 93838 306788 93894
rect 306838 93871 306894 93880
rect 307022 93936 307078 93945
rect 307022 93871 307078 93880
rect 306748 93832 306800 93838
rect 306748 93774 306800 93780
rect 306840 84244 306892 84250
rect 306840 84186 306892 84192
rect 306852 74594 306880 84186
rect 306748 74588 306800 74594
rect 306748 74530 306800 74536
rect 306840 74588 306892 74594
rect 306840 74530 306892 74536
rect 306760 46918 306788 74530
rect 306748 46912 306800 46918
rect 306748 46854 306800 46860
rect 306840 46844 306892 46850
rect 306840 46786 306892 46792
rect 306852 19378 306880 46786
rect 307666 28928 307722 28937
rect 307666 28863 307668 28872
rect 307720 28863 307722 28872
rect 307668 28834 307720 28840
rect 306748 19372 306800 19378
rect 306748 19314 306800 19320
rect 306840 19372 306892 19378
rect 306840 19314 306892 19320
rect 306564 13796 306616 13802
rect 306564 13738 306616 13744
rect 306472 11416 306524 11422
rect 306472 11358 306524 11364
rect 306760 9790 306788 19314
rect 306748 9784 306800 9790
rect 306748 9726 306800 9732
rect 306656 9716 306708 9722
rect 306656 9658 306708 9664
rect 306668 5846 306696 9658
rect 306656 5840 306708 5846
rect 306656 5782 306708 5788
rect 307772 5778 307800 335582
rect 307956 13054 307984 340054
rect 308048 340054 308338 340082
rect 308600 340054 308890 340082
rect 309244 340054 309350 340082
rect 309428 340054 309810 340082
rect 310072 340054 310362 340082
rect 310624 340054 310822 340082
rect 311084 340054 311282 340082
rect 311544 340054 311834 340082
rect 312004 340054 312294 340082
rect 307944 13048 307996 13054
rect 307944 12990 307996 12996
rect 308048 11354 308076 340054
rect 308600 335646 308628 340054
rect 308588 335640 308640 335646
rect 308588 335582 308640 335588
rect 309140 335640 309192 335646
rect 309140 335582 309192 335588
rect 309048 76288 309100 76294
rect 309046 76256 309048 76265
rect 309100 76256 309102 76265
rect 309046 76191 309102 76200
rect 308036 11348 308088 11354
rect 308036 11290 308088 11296
rect 307760 5772 307812 5778
rect 307760 5714 307812 5720
rect 309152 5710 309180 335582
rect 309244 9450 309272 340054
rect 309428 11286 309456 340054
rect 309784 337340 309836 337346
rect 309784 337282 309836 337288
rect 309416 11280 309468 11286
rect 309416 11222 309468 11228
rect 309232 9444 309284 9450
rect 309232 9386 309284 9392
rect 309140 5704 309192 5710
rect 309140 5646 309192 5652
rect 308588 4276 308640 4282
rect 308588 4218 308640 4224
rect 307390 3360 307446 3369
rect 307390 3295 307446 3304
rect 307404 480 307432 3295
rect 308600 480 308628 4218
rect 309796 4078 309824 337282
rect 310072 335646 310100 340054
rect 310060 335640 310112 335646
rect 310060 335582 310112 335588
rect 310520 335640 310572 335646
rect 310520 335582 310572 335588
rect 310532 5642 310560 335582
rect 310624 9518 310652 340054
rect 311084 331242 311112 340054
rect 311544 335646 311572 340054
rect 311532 335640 311584 335646
rect 311532 335582 311584 335588
rect 310808 331214 311112 331242
rect 310808 321638 310836 331214
rect 310796 321632 310848 321638
rect 310796 321574 310848 321580
rect 310888 321496 310940 321502
rect 310888 321438 310940 321444
rect 310900 311982 310928 321438
rect 310888 311976 310940 311982
rect 310888 311918 310940 311924
rect 310704 307896 310756 307902
rect 310704 307838 310756 307844
rect 310716 307766 310744 307838
rect 310704 307760 310756 307766
rect 310704 307702 310756 307708
rect 310888 298172 310940 298178
rect 310888 298114 310940 298120
rect 310900 293078 310928 298114
rect 310888 293072 310940 293078
rect 310888 293014 310940 293020
rect 310888 282804 310940 282810
rect 310888 282746 310940 282752
rect 310900 278730 310928 282746
rect 310888 278724 310940 278730
rect 310888 278666 310940 278672
rect 310888 263492 310940 263498
rect 310888 263434 310940 263440
rect 310900 256086 310928 263434
rect 310888 256080 310940 256086
rect 310888 256022 310940 256028
rect 310704 251320 310756 251326
rect 310704 251262 310756 251268
rect 310716 251190 310744 251262
rect 310704 251184 310756 251190
rect 310704 251126 310756 251132
rect 310888 241528 310940 241534
rect 310888 241470 310940 241476
rect 310900 234734 310928 241470
rect 310888 234728 310940 234734
rect 310888 234670 310940 234676
rect 310796 234592 310848 234598
rect 310796 234534 310848 234540
rect 310808 231810 310836 234534
rect 310796 231804 310848 231810
rect 310796 231746 310848 231752
rect 310888 222216 310940 222222
rect 310888 222158 310940 222164
rect 310900 215422 310928 222158
rect 310888 215416 310940 215422
rect 310888 215358 310940 215364
rect 310796 215280 310848 215286
rect 310796 215222 310848 215228
rect 310808 212498 310836 215222
rect 310796 212492 310848 212498
rect 310796 212434 310848 212440
rect 310888 202904 310940 202910
rect 310888 202846 310940 202852
rect 310900 196110 310928 202846
rect 310888 196104 310940 196110
rect 310888 196046 310940 196052
rect 310796 195968 310848 195974
rect 310796 195910 310848 195916
rect 310808 193225 310836 195910
rect 310794 193216 310850 193225
rect 310794 193151 310850 193160
rect 311070 193216 311126 193225
rect 311070 193151 311126 193160
rect 311084 183598 311112 193151
rect 310888 183592 310940 183598
rect 310888 183534 310940 183540
rect 311072 183592 311124 183598
rect 311072 183534 311124 183540
rect 310900 176798 310928 183534
rect 310888 176792 310940 176798
rect 310888 176734 310940 176740
rect 310796 176656 310848 176662
rect 310796 176598 310848 176604
rect 310808 167074 310836 176598
rect 310796 167068 310848 167074
rect 310796 167010 310848 167016
rect 310888 166932 310940 166938
rect 310888 166874 310940 166880
rect 310900 153377 310928 166874
rect 310886 153368 310942 153377
rect 310886 153303 310942 153312
rect 310794 153232 310850 153241
rect 310794 153167 310796 153176
rect 310848 153167 310850 153176
rect 310796 153138 310848 153144
rect 310796 147620 310848 147626
rect 310796 147562 310848 147568
rect 310808 143562 310836 147562
rect 310808 143534 310928 143562
rect 310900 138718 310928 143534
rect 310888 138712 310940 138718
rect 310888 138654 310940 138660
rect 310796 128308 310848 128314
rect 310796 128250 310848 128256
rect 310808 125610 310836 128250
rect 310808 125582 310928 125610
rect 310900 125526 310928 125582
rect 310888 125520 310940 125526
rect 310888 125462 310940 125468
rect 310796 116068 310848 116074
rect 310796 116010 310848 116016
rect 310808 115938 310836 116010
rect 310796 115932 310848 115938
rect 310796 115874 310848 115880
rect 310796 108996 310848 109002
rect 310796 108938 310848 108944
rect 310808 106298 310836 108938
rect 310808 106270 310928 106298
rect 310900 96830 310928 106270
rect 310888 96824 310940 96830
rect 310888 96766 310940 96772
rect 310796 96688 310848 96694
rect 310796 96630 310848 96636
rect 310808 91746 310836 96630
rect 310808 91718 310928 91746
rect 310900 77330 310928 91718
rect 310808 77302 310928 77330
rect 310808 67833 310836 77302
rect 310794 67824 310850 67833
rect 310794 67759 310850 67768
rect 310794 67688 310850 67697
rect 310794 67623 310850 67632
rect 310808 66230 310836 67623
rect 310796 66224 310848 66230
rect 310796 66166 310848 66172
rect 310796 60716 310848 60722
rect 310796 60658 310848 60664
rect 310808 56574 310836 60658
rect 310796 56568 310848 56574
rect 310796 56510 310848 56516
rect 310888 56568 310940 56574
rect 310888 56510 310940 56516
rect 310900 45558 310928 56510
rect 310888 45552 310940 45558
rect 310888 45494 310940 45500
rect 311072 45552 311124 45558
rect 311072 45494 311124 45500
rect 311084 27690 311112 45494
rect 310900 27662 311112 27690
rect 310900 26246 310928 27662
rect 310888 26240 310940 26246
rect 310888 26182 310940 26188
rect 310888 16652 310940 16658
rect 310888 16594 310940 16600
rect 310900 11218 310928 16594
rect 310888 11212 310940 11218
rect 310888 11154 310940 11160
rect 312004 9586 312032 340054
rect 312740 337278 312768 340068
rect 312728 337272 312780 337278
rect 312728 337214 312780 337220
rect 312544 337204 312596 337210
rect 312544 337146 312596 337152
rect 311992 9580 312044 9586
rect 311992 9522 312044 9528
rect 310612 9512 310664 9518
rect 310612 9454 310664 9460
rect 310520 5636 310572 5642
rect 310520 5578 310572 5584
rect 312082 4992 312138 5001
rect 312082 4927 312138 4936
rect 312096 4214 312124 4927
rect 312084 4208 312136 4214
rect 312084 4150 312136 4156
rect 312176 4208 312228 4214
rect 312176 4150 312228 4156
rect 309784 4072 309836 4078
rect 309784 4014 309836 4020
rect 310980 3392 311032 3398
rect 310980 3334 311032 3340
rect 309784 3120 309836 3126
rect 309784 3062 309836 3068
rect 309796 480 309824 3062
rect 310992 480 311020 3334
rect 312188 480 312216 4150
rect 312556 3058 312584 337146
rect 313292 5574 313320 340068
rect 313384 340054 313766 340082
rect 313384 9654 313412 340054
rect 314212 337142 314240 340068
rect 314778 340054 314884 340082
rect 314200 337136 314252 337142
rect 314200 337078 314252 337084
rect 314660 335640 314712 335646
rect 314660 335582 314712 335588
rect 314568 157480 314620 157486
rect 314566 157448 314568 157457
rect 314620 157448 314622 157457
rect 314566 157383 314622 157392
rect 313372 9648 313424 9654
rect 313372 9590 313424 9596
rect 313280 5568 313332 5574
rect 313280 5510 313332 5516
rect 314672 4865 314700 335582
rect 314856 12986 314884 340054
rect 314948 340054 315238 340082
rect 315408 340054 315698 340082
rect 314844 12980 314896 12986
rect 314844 12922 314896 12928
rect 314948 8906 314976 340054
rect 315408 335646 315436 340054
rect 316040 335708 316092 335714
rect 316040 335650 316092 335656
rect 315396 335640 315448 335646
rect 315396 335582 315448 335588
rect 315948 110628 316000 110634
rect 315948 110570 316000 110576
rect 315960 110537 315988 110570
rect 315946 110528 316002 110537
rect 315946 110463 316002 110472
rect 315946 28928 316002 28937
rect 315946 28863 315948 28872
rect 316000 28863 316002 28872
rect 315948 28834 316000 28840
rect 315946 16416 316002 16425
rect 315946 16351 316002 16360
rect 315960 16153 315988 16351
rect 315946 16144 316002 16153
rect 315946 16079 316002 16088
rect 314936 8900 314988 8906
rect 314936 8842 314988 8848
rect 315948 5024 316000 5030
rect 315946 4992 315948 5001
rect 316000 4992 316002 5001
rect 315946 4927 316002 4936
rect 314658 4856 314714 4865
rect 314658 4791 314714 4800
rect 316052 4758 316080 335650
rect 316132 335640 316184 335646
rect 316132 335582 316184 335588
rect 316144 8838 316172 335582
rect 316236 12918 316264 340068
rect 316328 340054 316710 340082
rect 316880 340054 317170 340082
rect 317616 340054 317722 340082
rect 317892 340054 318182 340082
rect 318352 340054 318642 340082
rect 318996 340054 319194 340082
rect 319272 340054 319654 340082
rect 319824 340054 320114 340082
rect 320284 340054 320666 340082
rect 320744 340054 321126 340082
rect 316328 335646 316356 340054
rect 316684 337136 316736 337142
rect 316684 337078 316736 337084
rect 316316 335640 316368 335646
rect 316316 335582 316368 335588
rect 316224 12912 316276 12918
rect 316224 12854 316276 12860
rect 316132 8832 316184 8838
rect 316132 8774 316184 8780
rect 316040 4752 316092 4758
rect 316040 4694 316092 4700
rect 314568 4072 314620 4078
rect 314568 4014 314620 4020
rect 313372 4004 313424 4010
rect 313372 3946 313424 3952
rect 312544 3052 312596 3058
rect 312544 2994 312596 3000
rect 313384 480 313412 3946
rect 314580 480 314608 4014
rect 316696 3262 316724 337078
rect 316880 335714 316908 340054
rect 316868 335708 316920 335714
rect 316868 335650 316920 335656
rect 317420 335640 317472 335646
rect 317420 335582 317472 335588
rect 317326 111072 317382 111081
rect 317326 111007 317382 111016
rect 317340 110537 317368 111007
rect 317326 110528 317382 110537
rect 317326 110463 317382 110472
rect 317328 76288 317380 76294
rect 317326 76256 317328 76265
rect 317380 76256 317382 76265
rect 317326 76191 317382 76200
rect 317326 29336 317382 29345
rect 317326 29271 317382 29280
rect 317340 28937 317368 29271
rect 317326 28928 317382 28937
rect 317326 28863 317382 28872
rect 317326 16688 317382 16697
rect 317326 16623 317382 16632
rect 317340 16425 317368 16623
rect 317326 16416 317382 16425
rect 317326 16351 317382 16360
rect 317432 4690 317460 335582
rect 317512 306400 317564 306406
rect 317512 306342 317564 306348
rect 317524 219434 317552 306342
rect 317512 219428 317564 219434
rect 317512 219370 317564 219376
rect 317512 209840 317564 209846
rect 317512 209782 317564 209788
rect 317524 200122 317552 209782
rect 317512 200116 317564 200122
rect 317512 200058 317564 200064
rect 317512 190528 317564 190534
rect 317512 190470 317564 190476
rect 317524 180810 317552 190470
rect 317512 180804 317564 180810
rect 317512 180746 317564 180752
rect 317512 142180 317564 142186
rect 317512 142122 317564 142128
rect 317524 137970 317552 142122
rect 317512 137964 317564 137970
rect 317512 137906 317564 137912
rect 317512 55276 317564 55282
rect 317512 55218 317564 55224
rect 317524 45558 317552 55218
rect 317512 45552 317564 45558
rect 317512 45494 317564 45500
rect 317512 31816 317564 31822
rect 317512 31758 317564 31764
rect 317524 8770 317552 31758
rect 317616 12850 317644 340054
rect 317892 335628 317920 340054
rect 318352 335646 318380 340054
rect 318800 335708 318852 335714
rect 318800 335650 318852 335656
rect 317708 335600 317920 335628
rect 318340 335640 318392 335646
rect 317708 306406 317736 335600
rect 318340 335582 318392 335588
rect 317696 306400 317748 306406
rect 317696 306342 317748 306348
rect 317696 219428 317748 219434
rect 317696 219370 317748 219376
rect 317708 209846 317736 219370
rect 317696 209840 317748 209846
rect 317696 209782 317748 209788
rect 317696 200116 317748 200122
rect 317696 200058 317748 200064
rect 317708 190534 317736 200058
rect 317696 190528 317748 190534
rect 317696 190470 317748 190476
rect 317696 180804 317748 180810
rect 317696 180746 317748 180752
rect 317708 142186 317736 180746
rect 317696 142180 317748 142186
rect 317696 142122 317748 142128
rect 317788 137964 317840 137970
rect 317788 137906 317840 137912
rect 317800 128330 317828 137906
rect 317708 128302 317828 128330
rect 317708 106282 317736 128302
rect 317696 106276 317748 106282
rect 317696 106218 317748 106224
rect 317880 106276 317932 106282
rect 317880 106218 317932 106224
rect 317892 96642 317920 106218
rect 317800 96626 317920 96642
rect 317788 96620 317920 96626
rect 317840 96614 317920 96620
rect 317788 96562 317840 96568
rect 317800 96531 317828 96562
rect 317788 89684 317840 89690
rect 317788 89626 317840 89632
rect 317800 86986 317828 89626
rect 317800 86958 317920 86986
rect 317892 86902 317920 86958
rect 317696 86896 317748 86902
rect 317696 86838 317748 86844
rect 317880 86896 317932 86902
rect 317880 86838 317932 86844
rect 317708 55282 317736 86838
rect 318706 76256 318762 76265
rect 318706 76191 318762 76200
rect 318720 75993 318748 76191
rect 318706 75984 318762 75993
rect 318706 75919 318762 75928
rect 317696 55276 317748 55282
rect 317696 55218 317748 55224
rect 317696 45552 317748 45558
rect 317696 45494 317748 45500
rect 317708 31822 317736 45494
rect 317696 31816 317748 31822
rect 317696 31758 317748 31764
rect 317604 12844 317656 12850
rect 317604 12786 317656 12792
rect 317512 8764 317564 8770
rect 317512 8706 317564 8712
rect 318708 4752 318760 4758
rect 318708 4694 318760 4700
rect 317420 4684 317472 4690
rect 317420 4626 317472 4632
rect 318720 3466 318748 4694
rect 318812 4622 318840 335650
rect 318892 335640 318944 335646
rect 318892 335582 318944 335588
rect 318904 8702 318932 335582
rect 318996 12782 319024 340054
rect 319272 335646 319300 340054
rect 319444 337000 319496 337006
rect 319444 336942 319496 336948
rect 319260 335640 319312 335646
rect 319260 335582 319312 335588
rect 318984 12776 319036 12782
rect 318984 12718 319036 12724
rect 318892 8696 318944 8702
rect 318892 8638 318944 8644
rect 318800 4616 318852 4622
rect 318800 4558 318852 4564
rect 318708 3460 318760 3466
rect 318708 3402 318760 3408
rect 316684 3256 316736 3262
rect 316684 3198 316736 3204
rect 318064 3256 318116 3262
rect 318064 3198 318116 3204
rect 315764 3052 315816 3058
rect 315764 2994 315816 3000
rect 315776 480 315804 2994
rect 316960 2984 317012 2990
rect 316960 2926 317012 2932
rect 316972 480 317000 2926
rect 318076 480 318104 3198
rect 319456 3194 319484 336942
rect 319824 335714 319852 340054
rect 319812 335708 319864 335714
rect 319812 335650 319864 335656
rect 320180 335640 320232 335646
rect 320180 335582 320232 335588
rect 320192 8634 320220 335582
rect 320284 12714 320312 340054
rect 320744 335646 320772 340054
rect 320732 335640 320784 335646
rect 320732 335582 320784 335588
rect 321468 329180 321520 329186
rect 321468 329122 321520 329128
rect 320272 12708 320324 12714
rect 320272 12650 320324 12656
rect 320180 8628 320232 8634
rect 320180 8570 320232 8576
rect 320364 4480 320416 4486
rect 320364 4422 320416 4428
rect 320376 3534 320404 4422
rect 321480 3534 321508 329122
rect 321572 4690 321600 340068
rect 321756 340054 322138 340082
rect 322216 340054 322598 340082
rect 322952 340054 323058 340082
rect 323136 340054 323518 340082
rect 323688 340054 324070 340082
rect 324332 340054 324530 340082
rect 324700 340054 324990 340082
rect 321652 335640 321704 335646
rect 321652 335582 321704 335588
rect 321664 8566 321692 335582
rect 321756 12646 321784 340054
rect 322216 335646 322244 340054
rect 322204 335640 322256 335646
rect 322204 335582 322256 335588
rect 322202 29336 322258 29345
rect 322202 29271 322258 29280
rect 322216 29073 322244 29271
rect 322202 29064 322258 29073
rect 322202 28999 322258 29008
rect 322202 16688 322258 16697
rect 322202 16623 322258 16632
rect 322216 16425 322244 16623
rect 322202 16416 322258 16425
rect 322202 16351 322258 16360
rect 321744 12640 321796 12646
rect 321744 12582 321796 12588
rect 321652 8560 321704 8566
rect 321652 8502 321704 8508
rect 321560 4684 321612 4690
rect 321560 4626 321612 4632
rect 322952 4622 322980 340054
rect 323136 12578 323164 340054
rect 323688 328506 323716 340054
rect 323308 328500 323360 328506
rect 323308 328442 323360 328448
rect 323676 328500 323728 328506
rect 323676 328442 323728 328448
rect 323320 311982 323348 328442
rect 323308 311976 323360 311982
rect 323308 311918 323360 311924
rect 323216 311908 323268 311914
rect 323216 311850 323268 311856
rect 323228 304314 323256 311850
rect 323228 304286 323440 304314
rect 323412 302138 323440 304286
rect 323320 302110 323440 302138
rect 323320 299470 323348 302110
rect 323308 299464 323360 299470
rect 323308 299406 323360 299412
rect 323308 288448 323360 288454
rect 323360 288396 323440 288402
rect 323308 288390 323440 288396
rect 323320 288374 323440 288390
rect 323412 283626 323440 288374
rect 323400 283620 323452 283626
rect 323400 283562 323452 283568
rect 323492 278792 323544 278798
rect 323490 278760 323492 278769
rect 323544 278760 323546 278769
rect 323490 278695 323546 278704
rect 323674 278760 323730 278769
rect 323674 278695 323730 278704
rect 323688 270314 323716 278695
rect 323504 270286 323716 270314
rect 323504 260982 323532 270286
rect 323400 260976 323452 260982
rect 323400 260918 323452 260924
rect 323492 260976 323544 260982
rect 323492 260918 323544 260924
rect 323412 259457 323440 260918
rect 323214 259448 323270 259457
rect 323214 259383 323270 259392
rect 323398 259448 323454 259457
rect 323398 259383 323454 259392
rect 323228 249830 323256 259383
rect 323216 249824 323268 249830
rect 323216 249766 323268 249772
rect 323492 249824 323544 249830
rect 323492 249766 323544 249772
rect 323504 241602 323532 249766
rect 323492 241596 323544 241602
rect 323492 241538 323544 241544
rect 323400 241528 323452 241534
rect 323400 241470 323452 241476
rect 323412 236722 323440 241470
rect 323412 236694 323532 236722
rect 323504 231878 323532 236694
rect 323308 231872 323360 231878
rect 323308 231814 323360 231820
rect 323492 231872 323544 231878
rect 323492 231814 323544 231820
rect 323320 227066 323348 231814
rect 323320 227038 323532 227066
rect 323504 224890 323532 227038
rect 323412 224862 323532 224890
rect 323412 217410 323440 224862
rect 323412 217382 323532 217410
rect 323504 212566 323532 217382
rect 323308 212560 323360 212566
rect 323308 212502 323360 212508
rect 323492 212560 323544 212566
rect 323492 212502 323544 212508
rect 323320 205698 323348 212502
rect 323308 205692 323360 205698
rect 323308 205634 323360 205640
rect 323400 205556 323452 205562
rect 323400 205498 323452 205504
rect 323412 198098 323440 205498
rect 323412 198070 323532 198098
rect 323504 193254 323532 198070
rect 323308 193248 323360 193254
rect 323306 193216 323308 193225
rect 323492 193248 323544 193254
rect 323360 193216 323362 193225
rect 323306 193151 323362 193160
rect 323490 193216 323492 193225
rect 323544 193216 323546 193225
rect 323490 193151 323546 193160
rect 323504 186266 323532 193151
rect 323412 186238 323532 186266
rect 323412 178786 323440 186238
rect 323412 178758 323532 178786
rect 323504 173942 323532 178758
rect 323308 173936 323360 173942
rect 323308 173878 323360 173884
rect 323492 173936 323544 173942
rect 323492 173878 323544 173884
rect 323320 169402 323348 173878
rect 323320 169374 323440 169402
rect 323412 157434 323440 169374
rect 323412 157406 323532 157434
rect 323504 157298 323532 157406
rect 323412 157270 323532 157298
rect 323412 144906 323440 157270
rect 323308 144900 323360 144906
rect 323308 144842 323360 144848
rect 323400 144900 323452 144906
rect 323400 144842 323452 144848
rect 323320 143546 323348 144842
rect 323308 143540 323360 143546
rect 323308 143482 323360 143488
rect 323492 143540 323544 143546
rect 323492 143482 323544 143488
rect 323504 128330 323532 143482
rect 323412 128302 323532 128330
rect 323412 125594 323440 128302
rect 323216 125588 323268 125594
rect 323216 125530 323268 125536
rect 323400 125588 323452 125594
rect 323400 125530 323452 125536
rect 323228 118674 323256 125530
rect 323228 118646 323348 118674
rect 323320 106298 323348 118646
rect 323320 106270 323440 106298
rect 323412 99482 323440 106270
rect 323400 99476 323452 99482
rect 323400 99418 323452 99424
rect 323400 99340 323452 99346
rect 323400 99282 323452 99288
rect 323412 77314 323440 99282
rect 323400 77308 323452 77314
rect 323400 77250 323452 77256
rect 323400 75948 323452 75954
rect 323400 75890 323452 75896
rect 323412 67658 323440 75890
rect 323308 67652 323360 67658
rect 323308 67594 323360 67600
rect 323400 67652 323452 67658
rect 323400 67594 323452 67600
rect 323320 66230 323348 67594
rect 323308 66224 323360 66230
rect 323308 66166 323360 66172
rect 323308 48340 323360 48346
rect 323308 48282 323360 48288
rect 323320 46918 323348 48282
rect 323308 46912 323360 46918
rect 323308 46854 323360 46860
rect 323308 37324 323360 37330
rect 323308 37266 323360 37272
rect 323320 34354 323348 37266
rect 323320 34326 323440 34354
rect 323412 28966 323440 34326
rect 323216 28960 323268 28966
rect 323216 28902 323268 28908
rect 323400 28960 323452 28966
rect 323400 28902 323452 28908
rect 323228 19394 323256 28902
rect 323228 19366 323348 19394
rect 323124 12572 323176 12578
rect 323124 12514 323176 12520
rect 323320 12510 323348 19366
rect 323308 12504 323360 12510
rect 323308 12446 323360 12452
rect 323124 12436 323176 12442
rect 323124 12378 323176 12384
rect 323136 8498 323164 12378
rect 323124 8492 323176 8498
rect 323124 8434 323176 8440
rect 324332 4758 324360 340054
rect 324700 335730 324728 340054
rect 324424 335702 324728 335730
rect 324424 7614 324452 335702
rect 325068 328506 325096 340190
rect 325712 340054 326002 340082
rect 326080 340054 326462 340082
rect 326632 340054 327014 340082
rect 327092 340054 327474 340082
rect 324688 328500 324740 328506
rect 324688 328442 324740 328448
rect 325056 328500 325108 328506
rect 325056 328442 325108 328448
rect 324700 311930 324728 328442
rect 324608 311902 324728 311930
rect 324608 304314 324636 311902
rect 324516 304286 324636 304314
rect 324516 302138 324544 304286
rect 324516 302110 324728 302138
rect 324700 299470 324728 302110
rect 324688 299464 324740 299470
rect 324688 299406 324740 299412
rect 324688 289876 324740 289882
rect 324688 289818 324740 289824
rect 324700 285002 324728 289818
rect 324700 284974 324820 285002
rect 324792 269142 324820 284974
rect 324596 269136 324648 269142
rect 324596 269078 324648 269084
rect 324780 269136 324832 269142
rect 324780 269078 324832 269084
rect 324608 260846 324636 269078
rect 324596 260840 324648 260846
rect 324596 260782 324648 260788
rect 324688 260772 324740 260778
rect 324688 260714 324740 260720
rect 324700 259418 324728 260714
rect 324688 259412 324740 259418
rect 324688 259354 324740 259360
rect 324780 259412 324832 259418
rect 324780 259354 324832 259360
rect 324792 231878 324820 259354
rect 324688 231872 324740 231878
rect 324688 231814 324740 231820
rect 324780 231872 324832 231878
rect 324780 231814 324832 231820
rect 324700 222222 324728 231814
rect 324688 222216 324740 222222
rect 324688 222158 324740 222164
rect 324780 222216 324832 222222
rect 324780 222158 324832 222164
rect 324792 212566 324820 222158
rect 324688 212560 324740 212566
rect 324688 212502 324740 212508
rect 324780 212560 324832 212566
rect 324780 212502 324832 212508
rect 324700 202910 324728 212502
rect 324596 202904 324648 202910
rect 324596 202846 324648 202852
rect 324688 202904 324740 202910
rect 324688 202846 324740 202852
rect 324608 193254 324636 202846
rect 324596 193248 324648 193254
rect 324596 193190 324648 193196
rect 324688 193248 324740 193254
rect 324688 193190 324740 193196
rect 324700 191826 324728 193190
rect 324688 191820 324740 191826
rect 324688 191762 324740 191768
rect 324872 191820 324924 191826
rect 324872 191762 324924 191768
rect 324884 182209 324912 191762
rect 324502 182200 324558 182209
rect 324502 182135 324504 182144
rect 324556 182135 324558 182144
rect 324870 182200 324926 182209
rect 324870 182135 324926 182144
rect 324504 182106 324556 182112
rect 324688 182096 324740 182102
rect 324688 182038 324740 182044
rect 324700 164234 324728 182038
rect 324608 164206 324728 164234
rect 324608 157434 324636 164206
rect 324516 157406 324636 157434
rect 324516 157298 324544 157406
rect 324516 157270 324636 157298
rect 324608 144906 324636 157270
rect 324596 144900 324648 144906
rect 324596 144842 324648 144848
rect 324780 144900 324832 144906
rect 324780 144842 324832 144848
rect 324792 139890 324820 144842
rect 324700 139862 324820 139890
rect 324700 128466 324728 139862
rect 324700 128438 324820 128466
rect 324792 125633 324820 128438
rect 324594 125624 324650 125633
rect 324594 125559 324596 125568
rect 324648 125559 324650 125568
rect 324778 125624 324834 125633
rect 324778 125559 324780 125568
rect 324596 125530 324648 125536
rect 324832 125559 324834 125568
rect 324780 125530 324832 125536
rect 324792 120578 324820 125530
rect 324700 120550 324820 120578
rect 324700 109698 324728 120550
rect 324516 109670 324728 109698
rect 324516 106264 324544 109670
rect 324516 106236 324636 106264
rect 324608 104825 324636 106236
rect 324594 104816 324650 104825
rect 324594 104751 324650 104760
rect 324778 104680 324834 104689
rect 324778 104615 324834 104624
rect 324792 95198 324820 104615
rect 324596 95192 324648 95198
rect 324596 95134 324648 95140
rect 324780 95192 324832 95198
rect 324780 95134 324832 95140
rect 324608 90420 324636 95134
rect 324608 90392 324728 90420
rect 324700 85542 324728 90392
rect 324688 85536 324740 85542
rect 324688 85478 324740 85484
rect 324596 75948 324648 75954
rect 324596 75890 324648 75896
rect 324608 72486 324636 75890
rect 324596 72480 324648 72486
rect 324596 72422 324648 72428
rect 324780 72480 324832 72486
rect 324780 72422 324832 72428
rect 324792 66230 324820 72422
rect 324780 66224 324832 66230
rect 324780 66166 324832 66172
rect 324688 56636 324740 56642
rect 324688 56578 324740 56584
rect 324700 48346 324728 56578
rect 324688 48340 324740 48346
rect 324688 48282 324740 48288
rect 324780 48340 324832 48346
rect 324780 48282 324832 48288
rect 324792 46918 324820 48282
rect 324780 46912 324832 46918
rect 324780 46854 324832 46860
rect 324688 37324 324740 37330
rect 324688 37266 324740 37272
rect 324700 18018 324728 37266
rect 324504 18012 324556 18018
rect 324504 17954 324556 17960
rect 324688 18012 324740 18018
rect 324688 17954 324740 17960
rect 324516 8430 324544 17954
rect 324504 8424 324556 8430
rect 324504 8366 324556 8372
rect 324412 7608 324464 7614
rect 324412 7550 324464 7556
rect 325608 5024 325660 5030
rect 325608 4966 325660 4972
rect 324320 4752 324372 4758
rect 324320 4694 324372 4700
rect 324228 4684 324280 4690
rect 324228 4626 324280 4632
rect 322940 4616 322992 4622
rect 322940 4558 322992 4564
rect 322848 4548 322900 4554
rect 322848 4490 322900 4496
rect 322860 3670 322888 4490
rect 322848 3664 322900 3670
rect 322848 3606 322900 3612
rect 320364 3528 320416 3534
rect 320364 3470 320416 3476
rect 320456 3528 320508 3534
rect 320456 3470 320508 3476
rect 321468 3528 321520 3534
rect 321468 3470 321520 3476
rect 324044 3528 324096 3534
rect 324044 3470 324096 3476
rect 319444 3188 319496 3194
rect 319444 3130 319496 3136
rect 319260 2916 319312 2922
rect 319260 2858 319312 2864
rect 319272 480 319300 2858
rect 320468 480 320496 3470
rect 321652 3460 321704 3466
rect 321652 3402 321704 3408
rect 321664 480 321692 3402
rect 322848 2916 322900 2922
rect 322848 2858 322900 2864
rect 322860 480 322888 2858
rect 324056 480 324084 3470
rect 324240 3058 324268 4626
rect 325620 3942 325648 4966
rect 325712 4894 325740 340054
rect 326080 335594 326108 340054
rect 325804 335566 326108 335594
rect 325804 7682 325832 335566
rect 326632 333334 326660 340054
rect 325884 333328 325936 333334
rect 325884 333270 325936 333276
rect 326620 333328 326672 333334
rect 326620 333270 326672 333276
rect 325896 328522 325924 333270
rect 325896 328494 326016 328522
rect 325988 317422 326016 328494
rect 325976 317416 326028 317422
rect 325976 317358 326028 317364
rect 325884 307828 325936 307834
rect 325884 307770 325936 307776
rect 325896 299470 325924 307770
rect 325884 299464 325936 299470
rect 325884 299406 325936 299412
rect 325976 299396 326028 299402
rect 325976 299338 326028 299344
rect 325988 298110 326016 299338
rect 325976 298104 326028 298110
rect 325976 298046 326028 298052
rect 326068 298104 326120 298110
rect 326068 298046 326120 298052
rect 326080 275210 326108 298046
rect 325988 275182 326108 275210
rect 325988 270502 326016 275182
rect 325976 270496 326028 270502
rect 325976 270438 326028 270444
rect 326068 270496 326120 270502
rect 326068 270438 326120 270444
rect 326080 255898 326108 270438
rect 325988 255870 326108 255898
rect 325988 251190 326016 255870
rect 325976 251184 326028 251190
rect 325976 251126 326028 251132
rect 326068 251184 326120 251190
rect 326068 251126 326120 251132
rect 326080 236586 326108 251126
rect 325988 236558 326108 236586
rect 325988 231849 326016 236558
rect 325974 231840 326030 231849
rect 325974 231775 326030 231784
rect 326066 231704 326122 231713
rect 326066 231639 326122 231648
rect 326080 217274 326108 231639
rect 325988 217246 326108 217274
rect 325988 212514 326016 217246
rect 325896 212486 326016 212514
rect 325896 202881 325924 212486
rect 325882 202872 325938 202881
rect 325882 202807 325938 202816
rect 325974 202736 326030 202745
rect 325974 202671 326030 202680
rect 325988 188442 326016 202671
rect 325896 188414 326016 188442
rect 325896 183569 325924 188414
rect 325882 183560 325938 183569
rect 325882 183495 325938 183504
rect 326066 183560 326122 183569
rect 326066 183495 326122 183504
rect 326080 182170 326108 183495
rect 326068 182164 326120 182170
rect 326068 182106 326120 182112
rect 326252 182164 326304 182170
rect 326252 182106 326304 182112
rect 326264 172553 326292 182106
rect 325974 172544 326030 172553
rect 325974 172479 326030 172488
rect 326250 172544 326306 172553
rect 326250 172479 326306 172488
rect 325988 166410 326016 172479
rect 325896 166382 326016 166410
rect 325896 162858 325924 166382
rect 325884 162852 325936 162858
rect 325884 162794 325936 162800
rect 326160 162852 326212 162858
rect 326160 162794 326212 162800
rect 326172 153241 326200 162794
rect 325974 153232 326030 153241
rect 325974 153167 326030 153176
rect 326158 153232 326214 153241
rect 326158 153167 326214 153176
rect 325988 145081 326016 153167
rect 325974 145072 326030 145081
rect 325974 145007 326030 145016
rect 325882 144936 325938 144945
rect 325882 144871 325884 144880
rect 325936 144871 325938 144880
rect 325884 144842 325936 144848
rect 325976 144832 326028 144838
rect 325976 144774 326028 144780
rect 325988 143546 326016 144774
rect 325976 143540 326028 143546
rect 325976 143482 326028 143488
rect 325976 132524 326028 132530
rect 325976 132466 326028 132472
rect 325988 118046 326016 132466
rect 325976 118040 326028 118046
rect 325976 117982 326028 117988
rect 325884 104916 325936 104922
rect 325884 104858 325936 104864
rect 325896 100042 325924 104858
rect 325896 100014 326016 100042
rect 325988 95334 326016 100014
rect 325976 95328 326028 95334
rect 325976 95270 326028 95276
rect 326068 95260 326120 95266
rect 326068 95202 326120 95208
rect 326080 87038 326108 95202
rect 326068 87032 326120 87038
rect 326068 86974 326120 86980
rect 325976 86964 326028 86970
rect 325976 86906 326028 86912
rect 325988 70514 326016 86906
rect 325976 70508 326028 70514
rect 325976 70450 326028 70456
rect 325884 70372 325936 70378
rect 325884 70314 325936 70320
rect 325896 58070 325924 70314
rect 325884 58064 325936 58070
rect 325884 58006 325936 58012
rect 325884 57928 325936 57934
rect 325884 57870 325936 57876
rect 325896 48278 325924 57870
rect 325884 48272 325936 48278
rect 325884 48214 325936 48220
rect 325976 48204 326028 48210
rect 325976 48146 326028 48152
rect 325988 46918 326016 48146
rect 325976 46912 326028 46918
rect 325976 46854 326028 46860
rect 326068 46912 326120 46918
rect 326068 46854 326120 46860
rect 326080 26058 326108 46854
rect 325988 26030 326108 26058
rect 325988 12510 326016 26030
rect 325976 12504 326028 12510
rect 325976 12446 326028 12452
rect 325884 12436 325936 12442
rect 325884 12378 325936 12384
rect 325896 8974 325924 12378
rect 325884 8968 325936 8974
rect 325884 8910 325936 8916
rect 325792 7676 325844 7682
rect 325792 7618 325844 7624
rect 327092 5574 327120 340054
rect 327552 339130 327580 340190
rect 328486 340054 328684 340082
rect 327460 339102 327580 339130
rect 327460 327146 327488 339102
rect 327724 336796 327776 336802
rect 327724 336738 327776 336744
rect 327264 327140 327316 327146
rect 327264 327082 327316 327088
rect 327448 327140 327500 327146
rect 327448 327082 327500 327088
rect 327276 309126 327304 327082
rect 327172 309120 327224 309126
rect 327172 309062 327224 309068
rect 327264 309120 327316 309126
rect 327264 309062 327316 309068
rect 327184 307766 327212 309062
rect 327172 307760 327224 307766
rect 327172 307702 327224 307708
rect 327264 298172 327316 298178
rect 327264 298114 327316 298120
rect 327276 289814 327304 298114
rect 327264 289808 327316 289814
rect 327264 289750 327316 289756
rect 327264 283620 327316 283626
rect 327264 283562 327316 283568
rect 327276 263702 327304 283562
rect 327264 263696 327316 263702
rect 327264 263638 327316 263644
rect 327172 263560 327224 263566
rect 327172 263502 327224 263508
rect 327184 251258 327212 263502
rect 327172 251252 327224 251258
rect 327172 251194 327224 251200
rect 327264 251252 327316 251258
rect 327264 251194 327316 251200
rect 327276 246378 327304 251194
rect 327276 246350 327396 246378
rect 327368 230518 327396 246350
rect 327172 230512 327224 230518
rect 327172 230454 327224 230460
rect 327356 230512 327408 230518
rect 327356 230454 327408 230460
rect 327184 220674 327212 230454
rect 327184 220646 327304 220674
rect 327276 207754 327304 220646
rect 327276 207726 327396 207754
rect 327368 197962 327396 207726
rect 327276 197934 327396 197962
rect 327276 186454 327304 197934
rect 327264 186448 327316 186454
rect 327264 186390 327316 186396
rect 327172 186312 327224 186318
rect 327172 186254 327224 186260
rect 327184 173942 327212 186254
rect 327172 173936 327224 173942
rect 327172 173878 327224 173884
rect 327264 173936 327316 173942
rect 327264 173878 327316 173884
rect 327276 164234 327304 173878
rect 327184 164206 327304 164234
rect 327184 157418 327212 164206
rect 327172 157412 327224 157418
rect 327172 157354 327224 157360
rect 327264 157276 327316 157282
rect 327264 157218 327316 157224
rect 327276 149818 327304 157218
rect 327276 149790 327396 149818
rect 327368 144945 327396 149790
rect 327170 144936 327226 144945
rect 327170 144871 327172 144880
rect 327224 144871 327226 144880
rect 327354 144936 327410 144945
rect 327354 144871 327356 144880
rect 327172 144842 327224 144848
rect 327408 144871 327410 144880
rect 327356 144842 327408 144848
rect 327368 137850 327396 144842
rect 327276 137822 327396 137850
rect 327276 135250 327304 137822
rect 327264 135244 327316 135250
rect 327264 135186 327316 135192
rect 327172 129736 327224 129742
rect 327172 129678 327224 129684
rect 327184 125594 327212 129678
rect 327172 125588 327224 125594
rect 327172 125530 327224 125536
rect 327356 125588 327408 125594
rect 327356 125530 327408 125536
rect 327368 117858 327396 125530
rect 327368 117830 327488 117858
rect 327460 113257 327488 117830
rect 327262 113248 327318 113257
rect 327262 113183 327318 113192
rect 327446 113248 327502 113257
rect 327446 113183 327502 113192
rect 327276 113150 327304 113183
rect 327264 113144 327316 113150
rect 327264 113086 327316 113092
rect 327172 103556 327224 103562
rect 327172 103498 327224 103504
rect 327184 103465 327212 103498
rect 327170 103456 327226 103465
rect 327170 103391 327226 103400
rect 327446 103320 327502 103329
rect 327446 103255 327502 103264
rect 327460 90438 327488 103255
rect 327264 90432 327316 90438
rect 327264 90374 327316 90380
rect 327448 90432 327500 90438
rect 327448 90374 327500 90380
rect 327276 72298 327304 90374
rect 327184 72270 327304 72298
rect 327184 58002 327212 72270
rect 327172 57996 327224 58002
rect 327172 57938 327224 57944
rect 327264 57860 327316 57866
rect 327264 57802 327316 57808
rect 327276 53122 327304 57802
rect 327184 53094 327304 53122
rect 327184 48278 327212 53094
rect 327172 48272 327224 48278
rect 327172 48214 327224 48220
rect 327356 48272 327408 48278
rect 327356 48214 327408 48220
rect 327368 46918 327396 48214
rect 327356 46912 327408 46918
rect 327356 46854 327408 46860
rect 327356 38548 327408 38554
rect 327356 38490 327408 38496
rect 327368 29034 327396 38490
rect 327172 29028 327224 29034
rect 327172 28970 327224 28976
rect 327356 29028 327408 29034
rect 327356 28970 327408 28976
rect 327184 18034 327212 28970
rect 327184 18006 327304 18034
rect 327276 17950 327304 18006
rect 327264 17944 327316 17950
rect 327264 17886 327316 17892
rect 327264 9648 327316 9654
rect 327264 9590 327316 9596
rect 327276 8344 327304 9590
rect 327184 8316 327304 8344
rect 327184 7002 327212 8316
rect 327172 6996 327224 7002
rect 327172 6938 327224 6944
rect 327080 5568 327132 5574
rect 327080 5510 327132 5516
rect 325700 4888 325752 4894
rect 325700 4830 325752 4836
rect 327080 4888 327132 4894
rect 327080 4830 327132 4836
rect 326528 4684 326580 4690
rect 326528 4626 326580 4632
rect 325608 3936 325660 3942
rect 325608 3878 325660 3884
rect 326436 3936 326488 3942
rect 326436 3878 326488 3884
rect 325240 3188 325292 3194
rect 325240 3130 325292 3136
rect 324228 3052 324280 3058
rect 324228 2994 324280 3000
rect 325252 480 325280 3130
rect 326448 480 326476 3878
rect 326540 3670 326568 4626
rect 326528 3664 326580 3670
rect 326528 3606 326580 3612
rect 327092 2922 327120 4830
rect 327632 3732 327684 3738
rect 327632 3674 327684 3680
rect 327080 2916 327132 2922
rect 327080 2858 327132 2864
rect 327644 480 327672 3674
rect 327736 3602 327764 336738
rect 328552 334552 328604 334558
rect 328552 334494 328604 334500
rect 328458 110936 328514 110945
rect 328458 110871 328514 110880
rect 328472 110673 328500 110871
rect 328458 110664 328514 110673
rect 328458 110599 328514 110608
rect 328274 16824 328330 16833
rect 328274 16759 328330 16768
rect 328288 16561 328316 16759
rect 328274 16552 328330 16561
rect 328274 16487 328330 16496
rect 328564 7750 328592 334494
rect 328656 9042 328684 340054
rect 328748 340054 328946 340082
rect 329024 340054 329406 340082
rect 329958 340054 330064 340082
rect 328644 9036 328696 9042
rect 328644 8978 328696 8984
rect 328552 7744 328604 7750
rect 328552 7686 328604 7692
rect 328748 4962 328776 340054
rect 329024 334558 329052 340054
rect 329840 335640 329892 335646
rect 329840 335582 329892 335588
rect 329012 334552 329064 334558
rect 329012 334494 329064 334500
rect 329852 5098 329880 335582
rect 329930 248432 329986 248441
rect 329930 248367 329986 248376
rect 329944 244254 329972 248367
rect 329932 244248 329984 244254
rect 329932 244190 329984 244196
rect 329930 220824 329986 220833
rect 329930 220759 329986 220768
rect 329944 202910 329972 220759
rect 329932 202904 329984 202910
rect 329930 202872 329932 202881
rect 329984 202872 329986 202881
rect 329930 202807 329986 202816
rect 329944 198082 329972 202807
rect 329932 198076 329984 198082
rect 329932 198018 329984 198024
rect 329932 162852 329984 162858
rect 329932 162794 329984 162800
rect 329944 153241 329972 162794
rect 329930 153232 329986 153241
rect 329930 153167 329986 153176
rect 329932 56636 329984 56642
rect 329932 56578 329984 56584
rect 329944 48385 329972 56578
rect 329930 48376 329986 48385
rect 329930 48311 329986 48320
rect 330036 9110 330064 340054
rect 330128 340054 330418 340082
rect 330588 340054 330878 340082
rect 330128 335646 330156 340054
rect 330588 336734 330616 340054
rect 330576 336728 330628 336734
rect 330576 336670 330628 336676
rect 331416 336122 331444 340068
rect 331508 340054 331890 340082
rect 331968 340054 332350 340082
rect 332796 340054 332902 340082
rect 333072 340054 333362 340082
rect 333440 340054 333822 340082
rect 334176 340054 334374 340082
rect 334544 340054 334834 340082
rect 334912 340054 335294 340082
rect 335464 340054 335846 340082
rect 336016 340054 336306 340082
rect 331404 336116 331456 336122
rect 331404 336058 331456 336064
rect 331508 335918 331536 340054
rect 331220 335912 331272 335918
rect 331220 335854 331272 335860
rect 331496 335912 331548 335918
rect 331496 335854 331548 335860
rect 330116 335640 330168 335646
rect 330116 335582 330168 335588
rect 330208 327208 330260 327214
rect 330208 327150 330260 327156
rect 330220 298178 330248 327150
rect 330116 298172 330168 298178
rect 330116 298114 330168 298120
rect 330208 298172 330260 298178
rect 330208 298114 330260 298120
rect 330128 296721 330156 298114
rect 330114 296712 330170 296721
rect 330114 296647 330170 296656
rect 330666 296712 330722 296721
rect 330666 296647 330722 296656
rect 330680 287094 330708 296647
rect 330484 287088 330536 287094
rect 330484 287030 330536 287036
rect 330668 287088 330720 287094
rect 330668 287030 330720 287036
rect 330220 278798 330248 278829
rect 330496 278798 330524 287030
rect 330208 278792 330260 278798
rect 330128 278740 330208 278746
rect 330128 278734 330260 278740
rect 330484 278792 330536 278798
rect 330484 278734 330536 278740
rect 330128 278718 330248 278734
rect 330128 273902 330156 278718
rect 330116 273896 330168 273902
rect 330116 273838 330168 273844
rect 330208 269136 330260 269142
rect 330206 269104 330208 269113
rect 330260 269104 330262 269113
rect 330206 269039 330262 269048
rect 330390 269104 330446 269113
rect 330390 269039 330446 269048
rect 330404 259486 330432 269039
rect 330116 259480 330168 259486
rect 330116 259422 330168 259428
rect 330392 259480 330444 259486
rect 330392 259422 330444 259428
rect 330128 258058 330156 259422
rect 330116 258052 330168 258058
rect 330116 257994 330168 258000
rect 330300 258052 330352 258058
rect 330300 257994 330352 258000
rect 330312 248441 330340 257994
rect 330298 248432 330354 248441
rect 330298 248367 330354 248376
rect 330208 244248 330260 244254
rect 330208 244190 330260 244196
rect 330220 227066 330248 244190
rect 330128 227038 330248 227066
rect 330128 222170 330156 227038
rect 330128 222142 330248 222170
rect 330220 220833 330248 222142
rect 330206 220824 330262 220833
rect 330206 220759 330262 220768
rect 330116 202904 330168 202910
rect 330114 202872 330116 202881
rect 330168 202872 330170 202881
rect 330114 202807 330170 202816
rect 330116 198076 330168 198082
rect 330116 198018 330168 198024
rect 330128 186998 330156 198018
rect 330116 186992 330168 186998
rect 330116 186934 330168 186940
rect 330300 186992 330352 186998
rect 330300 186934 330352 186940
rect 330312 182209 330340 186934
rect 330114 182200 330170 182209
rect 330114 182135 330170 182144
rect 330298 182200 330354 182209
rect 330298 182135 330354 182144
rect 330128 172514 330156 182135
rect 330116 172508 330168 172514
rect 330116 172450 330168 172456
rect 330300 172508 330352 172514
rect 330300 172450 330352 172456
rect 330312 162897 330340 172450
rect 330114 162888 330170 162897
rect 330114 162823 330116 162832
rect 330168 162823 330170 162832
rect 330298 162888 330354 162897
rect 330298 162823 330354 162832
rect 330116 162794 330168 162800
rect 330206 153232 330262 153241
rect 330206 153167 330262 153176
rect 330220 147642 330248 153167
rect 330128 147614 330248 147642
rect 330128 143546 330156 147614
rect 330116 143540 330168 143546
rect 330116 143482 330168 143488
rect 330208 138712 330260 138718
rect 330208 138654 330260 138660
rect 330220 125746 330248 138654
rect 330220 125718 330340 125746
rect 330312 124234 330340 125718
rect 330116 124228 330168 124234
rect 330116 124170 330168 124176
rect 330300 124228 330352 124234
rect 330300 124170 330352 124176
rect 330128 122806 330156 124170
rect 330116 122800 330168 122806
rect 330116 122742 330168 122748
rect 330116 113212 330168 113218
rect 330116 113154 330168 113160
rect 330128 103442 330156 113154
rect 330128 103414 330248 103442
rect 330220 98734 330248 103414
rect 330208 98728 330260 98734
rect 330208 98670 330260 98676
rect 330208 86964 330260 86970
rect 330208 86906 330260 86912
rect 330220 80730 330248 86906
rect 330128 80702 330248 80730
rect 330128 77194 330156 80702
rect 330128 77166 330340 77194
rect 330312 67658 330340 77166
rect 330116 67652 330168 67658
rect 330116 67594 330168 67600
rect 330300 67652 330352 67658
rect 330300 67594 330352 67600
rect 330128 66230 330156 67594
rect 330116 66224 330168 66230
rect 330116 66166 330168 66172
rect 330114 48376 330170 48385
rect 330114 48311 330170 48320
rect 330128 46918 330156 48311
rect 330116 46912 330168 46918
rect 330116 46854 330168 46860
rect 330116 37324 330168 37330
rect 330116 37266 330168 37272
rect 330128 28914 330156 37266
rect 330128 28886 330248 28914
rect 330220 27606 330248 28886
rect 330208 27600 330260 27606
rect 330208 27542 330260 27548
rect 330116 9716 330168 9722
rect 330116 9658 330168 9664
rect 330024 9104 330076 9110
rect 330024 9046 330076 9052
rect 330128 7818 330156 9658
rect 330116 7812 330168 7818
rect 330116 7754 330168 7760
rect 331232 5166 331260 335854
rect 331968 335510 331996 340054
rect 332692 335708 332744 335714
rect 332692 335650 332744 335656
rect 332600 335640 332652 335646
rect 332600 335582 332652 335588
rect 331312 335504 331364 335510
rect 331312 335446 331364 335452
rect 331956 335504 332008 335510
rect 331956 335446 332008 335452
rect 331324 86970 331352 335446
rect 331404 327140 331456 327146
rect 331404 327082 331456 327088
rect 331416 280158 331444 327082
rect 331404 280152 331456 280158
rect 331404 280094 331456 280100
rect 331404 270564 331456 270570
rect 331404 270506 331456 270512
rect 331416 241466 331444 270506
rect 331404 241460 331456 241466
rect 331404 241402 331456 241408
rect 331404 231872 331456 231878
rect 331404 231814 331456 231820
rect 331416 222193 331444 231814
rect 331402 222184 331458 222193
rect 331402 222119 331458 222128
rect 331586 222184 331642 222193
rect 331586 222119 331642 222128
rect 331600 212566 331628 222119
rect 331404 212560 331456 212566
rect 331404 212502 331456 212508
rect 331588 212560 331640 212566
rect 331588 212502 331640 212508
rect 331416 202881 331444 212502
rect 331402 202872 331458 202881
rect 331402 202807 331458 202816
rect 331586 202872 331642 202881
rect 331586 202807 331642 202816
rect 331600 193254 331628 202807
rect 331404 193248 331456 193254
rect 331404 193190 331456 193196
rect 331588 193248 331640 193254
rect 331588 193190 331640 193196
rect 331416 183569 331444 193190
rect 331402 183560 331458 183569
rect 331402 183495 331458 183504
rect 331586 183560 331642 183569
rect 331586 183495 331642 183504
rect 331600 173942 331628 183495
rect 331404 173936 331456 173942
rect 331404 173878 331456 173884
rect 331588 173936 331640 173942
rect 331588 173878 331640 173884
rect 331416 86970 331444 173878
rect 331312 86964 331364 86970
rect 331312 86906 331364 86912
rect 331404 86964 331456 86970
rect 331404 86906 331456 86912
rect 331312 86828 331364 86834
rect 331312 86770 331364 86776
rect 331404 86828 331456 86834
rect 331404 86770 331456 86776
rect 331324 7886 331352 86770
rect 331416 8362 331444 86770
rect 331862 29608 331918 29617
rect 331862 29543 331918 29552
rect 331876 29345 331904 29543
rect 331862 29336 331918 29345
rect 331862 29271 331918 29280
rect 331404 8356 331456 8362
rect 331404 8298 331456 8304
rect 331312 7880 331364 7886
rect 331312 7822 331364 7828
rect 332612 5234 332640 335582
rect 332704 7954 332732 335650
rect 332796 9178 332824 340054
rect 333072 335646 333100 340054
rect 333244 337272 333296 337278
rect 333244 337214 333296 337220
rect 333060 335640 333112 335646
rect 333060 335582 333112 335588
rect 332784 9172 332836 9178
rect 332784 9114 332836 9120
rect 332692 7948 332744 7954
rect 332692 7890 332744 7896
rect 332600 5228 332652 5234
rect 332600 5170 332652 5176
rect 331220 5160 331272 5166
rect 331220 5102 331272 5108
rect 329840 5092 329892 5098
rect 329840 5034 329892 5040
rect 328736 4956 328788 4962
rect 328736 4898 328788 4904
rect 328460 4820 328512 4826
rect 328460 4762 328512 4768
rect 328472 3942 328500 4762
rect 328460 3936 328512 3942
rect 328460 3878 328512 3884
rect 328828 3936 328880 3942
rect 328828 3878 328880 3884
rect 327724 3596 327776 3602
rect 327724 3538 327776 3544
rect 328840 480 328868 3878
rect 333256 3874 333284 337214
rect 333440 335714 333468 340054
rect 333428 335708 333480 335714
rect 333428 335650 333480 335656
rect 334072 335708 334124 335714
rect 334072 335650 334124 335656
rect 333980 335640 334032 335646
rect 333980 335582 334032 335588
rect 333612 4956 333664 4962
rect 333612 4898 333664 4904
rect 332416 3868 332468 3874
rect 332416 3810 332468 3816
rect 333244 3868 333296 3874
rect 333244 3810 333296 3816
rect 331312 3664 331364 3670
rect 331312 3606 331364 3612
rect 331324 3210 331352 3606
rect 331232 3182 331352 3210
rect 330024 2848 330076 2854
rect 330024 2790 330076 2796
rect 330036 480 330064 2790
rect 331232 480 331260 3182
rect 332428 480 332456 3810
rect 333624 480 333652 4898
rect 333992 4622 334020 335582
rect 334084 8022 334112 335650
rect 334176 9246 334204 340054
rect 334544 335646 334572 340054
rect 334912 335714 334940 340054
rect 335268 337068 335320 337074
rect 335268 337010 335320 337016
rect 334900 335708 334952 335714
rect 334900 335650 334952 335656
rect 334532 335640 334584 335646
rect 334532 335582 334584 335588
rect 334164 9240 334216 9246
rect 334164 9182 334216 9188
rect 334072 8016 334124 8022
rect 334072 7958 334124 7964
rect 333980 4616 334032 4622
rect 333980 4558 334032 4564
rect 335280 3874 335308 337010
rect 335360 334212 335412 334218
rect 335360 334154 335412 334160
rect 335372 4486 335400 334154
rect 335464 6662 335492 340054
rect 336016 334218 336044 340054
rect 336096 337680 336148 337686
rect 336096 337622 336148 337628
rect 336004 334212 336056 334218
rect 336004 334154 336056 334160
rect 336108 334098 336136 337622
rect 336016 334070 336136 334098
rect 335452 6656 335504 6662
rect 335452 6598 335504 6604
rect 335360 4480 335412 4486
rect 335360 4422 335412 4428
rect 334716 3868 334768 3874
rect 334716 3810 334768 3816
rect 335268 3868 335320 3874
rect 335268 3810 335320 3816
rect 334728 480 334756 3810
rect 336016 3074 336044 334070
rect 336752 332042 336780 340068
rect 336844 340054 337318 340082
rect 336740 332036 336792 332042
rect 336740 331978 336792 331984
rect 336844 331362 336872 340054
rect 337396 335594 337424 340190
rect 338238 340054 338344 340082
rect 337120 335566 337424 335594
rect 338120 335640 338172 335646
rect 338120 335582 338172 335588
rect 336924 332036 336976 332042
rect 336924 331978 336976 331984
rect 336832 331356 336884 331362
rect 336832 331298 336884 331304
rect 336832 331220 336884 331226
rect 336832 331162 336884 331168
rect 336844 77382 336872 331162
rect 336936 87242 336964 331978
rect 337120 331208 337148 335566
rect 337120 331180 337240 331208
rect 337212 321638 337240 331180
rect 337200 321632 337252 321638
rect 337200 321574 337252 321580
rect 337200 320884 337252 320890
rect 337200 320826 337252 320832
rect 337212 317422 337240 320826
rect 337200 317416 337252 317422
rect 337200 317358 337252 317364
rect 337200 311772 337252 311778
rect 337200 311714 337252 311720
rect 337212 307766 337240 311714
rect 337200 307760 337252 307766
rect 337200 307702 337252 307708
rect 337292 298172 337344 298178
rect 337292 298114 337344 298120
rect 337304 292602 337332 298114
rect 337108 292596 337160 292602
rect 337108 292538 337160 292544
rect 337292 292596 337344 292602
rect 337292 292538 337344 292544
rect 337120 287065 337148 292538
rect 337106 287056 337162 287065
rect 337106 286991 337162 287000
rect 337290 287056 337346 287065
rect 337290 286991 337346 287000
rect 337304 285666 337332 286991
rect 337292 285660 337344 285666
rect 337292 285602 337344 285608
rect 337200 276072 337252 276078
rect 337200 276014 337252 276020
rect 337212 266354 337240 276014
rect 337016 266348 337068 266354
rect 337016 266290 337068 266296
rect 337200 266348 337252 266354
rect 337200 266290 337252 266296
rect 337028 256737 337056 266290
rect 337014 256728 337070 256737
rect 337014 256663 337070 256672
rect 337198 256728 337254 256737
rect 337198 256663 337254 256672
rect 337212 254046 337240 256663
rect 337200 254040 337252 254046
rect 337200 253982 337252 253988
rect 337108 247172 337160 247178
rect 337108 247114 337160 247120
rect 337120 247042 337148 247114
rect 337108 247036 337160 247042
rect 337108 246978 337160 246984
rect 337108 244248 337160 244254
rect 337108 244190 337160 244196
rect 337120 237402 337148 244190
rect 337120 237374 337240 237402
rect 337212 231674 337240 237374
rect 337200 231668 337252 231674
rect 337200 231610 337252 231616
rect 337292 220856 337344 220862
rect 337292 220798 337344 220804
rect 337304 212634 337332 220798
rect 337292 212628 337344 212634
rect 337292 212570 337344 212576
rect 337200 212492 337252 212498
rect 337200 212434 337252 212440
rect 337212 211138 337240 212434
rect 337200 211132 337252 211138
rect 337200 211074 337252 211080
rect 337384 211132 337436 211138
rect 337384 211074 337436 211080
rect 337396 201521 337424 211074
rect 337106 201512 337162 201521
rect 337106 201447 337162 201456
rect 337382 201512 337438 201521
rect 337382 201447 337438 201456
rect 337120 193390 337148 201447
rect 337108 193384 337160 193390
rect 337108 193326 337160 193332
rect 337108 193248 337160 193254
rect 337108 193190 337160 193196
rect 337120 188578 337148 193190
rect 337120 188550 337424 188578
rect 337396 173942 337424 188550
rect 337108 173936 337160 173942
rect 337108 173878 337160 173884
rect 337384 173936 337436 173942
rect 337384 173878 337436 173884
rect 337120 172514 337148 173878
rect 337108 172508 337160 172514
rect 337108 172450 337160 172456
rect 337108 164212 337160 164218
rect 337108 164154 337160 164160
rect 337120 162874 337148 164154
rect 337120 162846 337240 162874
rect 337212 154562 337240 162846
rect 337200 154556 337252 154562
rect 337200 154498 337252 154504
rect 337292 152380 337344 152386
rect 337292 152322 337344 152328
rect 337304 135289 337332 152322
rect 337106 135280 337162 135289
rect 337106 135215 337162 135224
rect 337290 135280 337346 135289
rect 337290 135215 337346 135224
rect 337120 133890 337148 135215
rect 337108 133884 337160 133890
rect 337108 133826 337160 133832
rect 337200 124228 337252 124234
rect 337200 124170 337252 124176
rect 337212 122806 337240 124170
rect 337200 122800 337252 122806
rect 337200 122742 337252 122748
rect 337200 118040 337252 118046
rect 337200 117982 337252 117988
rect 337212 109698 337240 117982
rect 337120 109670 337240 109698
rect 337120 103494 337148 109670
rect 337108 103488 337160 103494
rect 337108 103430 337160 103436
rect 337200 93900 337252 93906
rect 337200 93842 337252 93848
rect 337212 90438 337240 93842
rect 337016 90432 337068 90438
rect 337016 90374 337068 90380
rect 337200 90432 337252 90438
rect 337200 90374 337252 90380
rect 336924 87236 336976 87242
rect 336924 87178 336976 87184
rect 336924 87032 336976 87038
rect 336924 86974 336976 86980
rect 336936 77382 336964 86974
rect 337028 84182 337056 90374
rect 337016 84176 337068 84182
rect 337016 84118 337068 84124
rect 336832 77376 336884 77382
rect 336832 77318 336884 77324
rect 336924 77376 336976 77382
rect 336924 77318 336976 77324
rect 336832 77240 336884 77246
rect 336832 77182 336884 77188
rect 336924 77240 336976 77246
rect 336924 77182 336976 77188
rect 336740 16720 336792 16726
rect 336738 16688 336740 16697
rect 336792 16688 336794 16697
rect 336738 16623 336794 16632
rect 336844 6730 336872 77182
rect 336936 8090 336964 77182
rect 337200 66292 337252 66298
rect 337200 66234 337252 66240
rect 337212 60874 337240 66234
rect 337212 60846 337332 60874
rect 337304 58834 337332 60846
rect 337212 58806 337332 58834
rect 337212 50946 337240 58806
rect 337120 50918 337240 50946
rect 337120 41154 337148 50918
rect 337120 41126 337240 41154
rect 337212 24342 337240 41126
rect 337200 24336 337252 24342
rect 337200 24278 337252 24284
rect 337108 19372 337160 19378
rect 337108 19314 337160 19320
rect 337120 12510 337148 19314
rect 337108 12504 337160 12510
rect 337108 12446 337160 12452
rect 337016 12436 337068 12442
rect 337016 12378 337068 12384
rect 336924 8084 336976 8090
rect 336924 8026 336976 8032
rect 336832 6724 336884 6730
rect 336832 6666 336884 6672
rect 337028 4554 337056 12378
rect 337108 5092 337160 5098
rect 337108 5034 337160 5040
rect 337016 4548 337068 4554
rect 337016 4490 337068 4496
rect 335924 3058 336044 3074
rect 335912 3052 336044 3058
rect 335964 3046 336044 3052
rect 336096 3052 336148 3058
rect 335912 2994 335964 3000
rect 336096 2994 336148 3000
rect 336108 2938 336136 2994
rect 335924 2910 336136 2938
rect 335924 480 335952 2910
rect 337120 480 337148 5034
rect 338132 5030 338160 335582
rect 338210 16960 338266 16969
rect 338210 16895 338266 16904
rect 338224 16726 338252 16895
rect 338212 16720 338264 16726
rect 338212 16662 338264 16668
rect 338316 8158 338344 340054
rect 338408 340054 338790 340082
rect 338960 340054 339250 340082
rect 339604 340054 339710 340082
rect 338304 8152 338356 8158
rect 338304 8094 338356 8100
rect 338408 6594 338436 340054
rect 338960 335646 338988 340054
rect 338948 335640 339000 335646
rect 338948 335582 339000 335588
rect 338856 328500 338908 328506
rect 338856 328442 338908 328448
rect 338868 311930 338896 328442
rect 338776 311902 338896 311930
rect 338776 311794 338804 311902
rect 338776 311766 338896 311794
rect 338868 302258 338896 311766
rect 338856 302252 338908 302258
rect 338856 302194 338908 302200
rect 338948 302116 339000 302122
rect 338948 302058 339000 302064
rect 338960 299470 338988 302058
rect 338948 299464 339000 299470
rect 338948 299406 339000 299412
rect 338856 299396 338908 299402
rect 338856 299338 338908 299344
rect 338868 280158 338896 299338
rect 338856 280152 338908 280158
rect 338856 280094 338908 280100
rect 338856 270564 338908 270570
rect 338856 270506 338908 270512
rect 338868 260846 338896 270506
rect 338856 260840 338908 260846
rect 338856 260782 338908 260788
rect 338856 251252 338908 251258
rect 338856 251194 338908 251200
rect 338868 241505 338896 251194
rect 338670 241496 338726 241505
rect 338670 241431 338726 241440
rect 338854 241496 338910 241505
rect 338854 241431 338910 241440
rect 338684 231878 338712 241431
rect 338672 231872 338724 231878
rect 338672 231814 338724 231820
rect 338856 231872 338908 231878
rect 338856 231814 338908 231820
rect 338868 222193 338896 231814
rect 338670 222184 338726 222193
rect 338670 222119 338726 222128
rect 338854 222184 338910 222193
rect 338854 222119 338910 222128
rect 338684 212566 338712 222119
rect 338672 212560 338724 212566
rect 338672 212502 338724 212508
rect 338856 212560 338908 212566
rect 338856 212502 338908 212508
rect 338868 202881 338896 212502
rect 338670 202872 338726 202881
rect 338670 202807 338726 202816
rect 338854 202872 338910 202881
rect 338854 202807 338910 202816
rect 338684 193254 338712 202807
rect 338672 193248 338724 193254
rect 338672 193190 338724 193196
rect 338856 193248 338908 193254
rect 338856 193190 338908 193196
rect 338868 176662 338896 193190
rect 338856 176656 338908 176662
rect 338856 176598 338908 176604
rect 338856 176520 338908 176526
rect 338856 176462 338908 176468
rect 338868 154737 338896 176462
rect 338854 154728 338910 154737
rect 339604 154698 339632 340054
rect 340248 337414 340276 340068
rect 340236 337408 340288 337414
rect 340236 337350 340288 337356
rect 340340 328506 340368 340190
rect 340984 340054 341182 340082
rect 340788 337408 340840 337414
rect 340788 337350 340840 337356
rect 339776 328500 339828 328506
rect 339776 328442 339828 328448
rect 340328 328500 340380 328506
rect 340328 328442 340380 328448
rect 339788 311930 339816 328442
rect 339696 311902 339816 311930
rect 339696 311794 339724 311902
rect 339696 311766 339816 311794
rect 339788 282962 339816 311766
rect 339696 282934 339816 282962
rect 339696 282826 339724 282934
rect 339696 282798 339816 282826
rect 339788 263650 339816 282798
rect 339696 263622 339816 263650
rect 339696 263514 339724 263622
rect 339696 263486 339816 263514
rect 339788 244338 339816 263486
rect 339696 244310 339816 244338
rect 339696 244202 339724 244310
rect 339696 244174 339816 244202
rect 339788 225026 339816 244174
rect 339696 224998 339816 225026
rect 339696 224890 339724 224998
rect 339696 224862 339816 224890
rect 339788 205714 339816 224862
rect 339696 205686 339816 205714
rect 339696 205578 339724 205686
rect 339696 205550 339816 205578
rect 339788 188426 339816 205550
rect 339776 188420 339828 188426
rect 339776 188362 339828 188368
rect 339868 183592 339920 183598
rect 339868 183534 339920 183540
rect 339880 173942 339908 183534
rect 339684 173936 339736 173942
rect 339684 173878 339736 173884
rect 339868 173936 339920 173942
rect 339868 173878 339920 173884
rect 339696 156618 339724 173878
rect 339696 156590 339816 156618
rect 338854 154663 338910 154672
rect 339592 154692 339644 154698
rect 339592 154634 339644 154640
rect 338854 154592 338910 154601
rect 338854 154527 338910 154536
rect 339592 154556 339644 154562
rect 338868 147694 338896 154527
rect 339592 154498 339644 154504
rect 338856 147688 338908 147694
rect 338856 147630 338908 147636
rect 338948 147620 339000 147626
rect 338948 147562 339000 147568
rect 338776 138038 338804 138069
rect 338960 138038 338988 147562
rect 338764 138032 338816 138038
rect 338948 138032 339000 138038
rect 338816 137980 338896 137986
rect 338764 137974 338896 137980
rect 338948 137974 339000 137980
rect 338776 137958 338896 137974
rect 338868 99498 338896 137958
rect 338776 99470 338896 99498
rect 338776 99362 338804 99470
rect 338776 99334 338896 99362
rect 338868 80102 338896 99334
rect 338856 80096 338908 80102
rect 338856 80038 338908 80044
rect 338856 79960 338908 79966
rect 338856 79902 338908 79908
rect 338868 60874 338896 79902
rect 338868 60846 338988 60874
rect 338960 58834 338988 60846
rect 338868 58806 338988 58834
rect 338868 51762 338896 58806
rect 338868 51734 338988 51762
rect 338960 46918 338988 51734
rect 338488 46912 338540 46918
rect 338488 46854 338540 46860
rect 338948 46912 339000 46918
rect 338948 46854 339000 46860
rect 338500 45558 338528 46854
rect 338488 45552 338540 45558
rect 338488 45494 338540 45500
rect 338672 27668 338724 27674
rect 338672 27610 338724 27616
rect 338684 19378 338712 27610
rect 338672 19372 338724 19378
rect 338672 19314 338724 19320
rect 338856 19372 338908 19378
rect 338856 19314 338908 19320
rect 338868 14498 338896 19314
rect 338776 14470 338896 14498
rect 338396 6588 338448 6594
rect 338396 6530 338448 6536
rect 338120 5024 338172 5030
rect 338120 4966 338172 4972
rect 338776 3874 338804 14470
rect 339604 8226 339632 154498
rect 339788 151858 339816 156590
rect 339788 151830 339908 151858
rect 339880 151774 339908 151830
rect 339868 151768 339920 151774
rect 339868 151710 339920 151716
rect 339776 142180 339828 142186
rect 339776 142122 339828 142128
rect 339788 99498 339816 142122
rect 339696 99470 339816 99498
rect 339696 95198 339724 99470
rect 339684 95192 339736 95198
rect 339684 95134 339736 95140
rect 339776 77308 339828 77314
rect 339776 77250 339828 77256
rect 339788 56658 339816 77250
rect 339696 56630 339816 56658
rect 339696 56574 339724 56630
rect 339684 56568 339736 56574
rect 339684 56510 339736 56516
rect 339960 46980 340012 46986
rect 339960 46922 340012 46928
rect 339972 37330 340000 46922
rect 339776 37324 339828 37330
rect 339776 37266 339828 37272
rect 339960 37324 340012 37330
rect 339960 37266 340012 37272
rect 339788 12458 339816 37266
rect 339696 12430 339816 12458
rect 339592 8220 339644 8226
rect 339592 8162 339644 8168
rect 339696 6526 339724 12430
rect 339684 6520 339736 6526
rect 339684 6462 339736 6468
rect 338764 3868 338816 3874
rect 338764 3810 338816 3816
rect 338304 3732 338356 3738
rect 338304 3674 338356 3680
rect 338316 480 338344 3674
rect 340800 3330 340828 337350
rect 340984 8294 341012 340054
rect 341628 337550 341656 340068
rect 341720 340054 342194 340082
rect 342364 340054 342654 340082
rect 341616 337544 341668 337550
rect 341616 337486 341668 337492
rect 341720 335578 341748 340054
rect 341800 337204 341852 337210
rect 341800 337146 341852 337152
rect 341708 335572 341760 335578
rect 341708 335514 341760 335520
rect 341812 335458 341840 337146
rect 341536 335430 341840 335458
rect 341432 328500 341484 328506
rect 341432 328442 341484 328448
rect 341444 321638 341472 328442
rect 341432 321632 341484 321638
rect 341432 321574 341484 321580
rect 341432 318844 341484 318850
rect 341432 318786 341484 318792
rect 341444 311914 341472 318786
rect 341248 311908 341300 311914
rect 341248 311850 341300 311856
rect 341432 311908 341484 311914
rect 341432 311850 341484 311856
rect 341260 309126 341288 311850
rect 341248 309120 341300 309126
rect 341248 309062 341300 309068
rect 341156 299532 341208 299538
rect 341156 299474 341208 299480
rect 341168 299418 341196 299474
rect 341168 299390 341288 299418
rect 341260 292618 341288 299390
rect 341168 292590 341288 292618
rect 341168 282946 341196 292590
rect 341156 282940 341208 282946
rect 341156 282882 341208 282888
rect 341156 280220 341208 280226
rect 341156 280162 341208 280168
rect 341168 280106 341196 280162
rect 341168 280078 341380 280106
rect 341352 273170 341380 280078
rect 341168 273142 341380 273170
rect 341168 270586 341196 273142
rect 341168 270558 341288 270586
rect 341260 270502 341288 270558
rect 341248 270496 341300 270502
rect 341248 270438 341300 270444
rect 341432 270496 341484 270502
rect 341432 270438 341484 270444
rect 341444 260953 341472 270438
rect 341062 260944 341118 260953
rect 341062 260879 341118 260888
rect 341430 260944 341486 260953
rect 341430 260879 341486 260888
rect 341076 260846 341104 260879
rect 341064 260840 341116 260846
rect 341064 260782 341116 260788
rect 341064 253768 341116 253774
rect 341064 253710 341116 253716
rect 341076 231878 341104 253710
rect 341064 231872 341116 231878
rect 341064 231814 341116 231820
rect 341156 231872 341208 231878
rect 341156 231814 341208 231820
rect 341168 225010 341196 231814
rect 341156 225004 341208 225010
rect 341156 224946 341208 224952
rect 341064 222216 341116 222222
rect 341064 222158 341116 222164
rect 341076 215234 341104 222158
rect 341076 215206 341288 215234
rect 341260 209778 341288 215206
rect 341248 209772 341300 209778
rect 341248 209714 341300 209720
rect 341340 209772 341392 209778
rect 341340 209714 341392 209720
rect 341352 198762 341380 209714
rect 341248 198756 341300 198762
rect 341248 198698 341300 198704
rect 341340 198756 341392 198762
rect 341340 198698 341392 198704
rect 341260 189038 341288 198698
rect 341248 189032 341300 189038
rect 341248 188974 341300 188980
rect 341432 189032 341484 189038
rect 341432 188974 341484 188980
rect 341444 179489 341472 188974
rect 341246 179480 341302 179489
rect 341246 179415 341302 179424
rect 341430 179480 341486 179489
rect 341430 179415 341486 179424
rect 341260 179382 341288 179415
rect 341248 179376 341300 179382
rect 341248 179318 341300 179324
rect 341248 169788 341300 169794
rect 341248 169730 341300 169736
rect 341260 160070 341288 169730
rect 341248 160064 341300 160070
rect 341248 160006 341300 160012
rect 341248 143404 341300 143410
rect 341248 143346 341300 143352
rect 341260 132569 341288 143346
rect 341062 132560 341118 132569
rect 341062 132495 341118 132504
rect 341246 132560 341302 132569
rect 341246 132495 341302 132504
rect 341076 123978 341104 132495
rect 341076 123950 341288 123978
rect 341260 122754 341288 123950
rect 341168 122726 341288 122754
rect 341168 118130 341196 122726
rect 341168 118102 341288 118130
rect 341260 104938 341288 118102
rect 341168 104910 341288 104938
rect 341168 103494 341196 104910
rect 341156 103488 341208 103494
rect 341156 103430 341208 103436
rect 341064 77308 341116 77314
rect 341064 77250 341116 77256
rect 341076 77178 341104 77250
rect 341064 77172 341116 77178
rect 341064 77114 341116 77120
rect 341156 70304 341208 70310
rect 341156 70246 341208 70252
rect 341168 60722 341196 70246
rect 341156 60716 341208 60722
rect 341156 60658 341208 60664
rect 341340 60716 341392 60722
rect 341340 60658 341392 60664
rect 341352 57934 341380 60658
rect 341340 57928 341392 57934
rect 341340 57870 341392 57876
rect 341432 50924 341484 50930
rect 341432 50866 341484 50872
rect 341444 41478 341472 50866
rect 341432 41472 341484 41478
rect 341432 41414 341484 41420
rect 341432 38616 341484 38622
rect 341432 38558 341484 38564
rect 341444 29034 341472 38558
rect 341156 29028 341208 29034
rect 341156 28970 341208 28976
rect 341432 29028 341484 29034
rect 341432 28970 341484 28976
rect 341168 24154 341196 28970
rect 341168 24126 341288 24154
rect 340972 8288 341024 8294
rect 340972 8230 341024 8236
rect 341260 6458 341288 24126
rect 341248 6452 341300 6458
rect 341248 6394 341300 6400
rect 341536 3874 341564 335430
rect 342364 6186 342392 340054
rect 342904 337136 342956 337142
rect 342904 337078 342956 337084
rect 342352 6180 342404 6186
rect 342352 6122 342404 6128
rect 342916 4146 342944 337078
rect 343100 336802 343128 340068
rect 343088 336796 343140 336802
rect 343088 336738 343140 336744
rect 343652 6390 343680 340068
rect 344112 337482 344140 340068
rect 344572 337686 344600 340068
rect 345138 340054 345244 340082
rect 344560 337680 344612 337686
rect 344560 337622 344612 337628
rect 344376 337544 344428 337550
rect 344376 337486 344428 337492
rect 344100 337476 344152 337482
rect 344100 337418 344152 337424
rect 344284 336864 344336 336870
rect 344284 336806 344336 336812
rect 343640 6384 343692 6390
rect 343640 6326 343692 6332
rect 344296 4146 344324 336806
rect 342904 4140 342956 4146
rect 342904 4082 342956 4088
rect 343640 4140 343692 4146
rect 343640 4082 343692 4088
rect 344284 4140 344336 4146
rect 344284 4082 344336 4088
rect 341524 3868 341576 3874
rect 341524 3810 341576 3816
rect 341892 3868 341944 3874
rect 341892 3810 341944 3816
rect 341156 3392 341208 3398
rect 340892 3340 341156 3346
rect 340892 3334 341208 3340
rect 339500 3324 339552 3330
rect 339500 3266 339552 3272
rect 340788 3324 340840 3330
rect 340788 3266 340840 3272
rect 340892 3318 341196 3334
rect 339512 480 339540 3266
rect 340892 3210 340920 3318
rect 340708 3182 340920 3210
rect 340708 480 340736 3182
rect 341904 480 341932 3810
rect 343088 3800 343140 3806
rect 343088 3742 343140 3748
rect 343100 480 343128 3742
rect 343652 2854 343680 4082
rect 344388 2990 344416 337486
rect 345216 6254 345244 340054
rect 345584 337618 345612 340068
rect 345676 340054 346058 340082
rect 345572 337612 345624 337618
rect 345572 337554 345624 337560
rect 345676 336954 345704 340054
rect 345492 336938 345704 336954
rect 345480 336932 345704 336938
rect 345532 336926 345704 336932
rect 345940 336932 345992 336938
rect 345480 336874 345532 336880
rect 345940 336874 345992 336880
rect 345952 331242 345980 336874
rect 345676 331214 345980 331242
rect 345204 6248 345256 6254
rect 345204 6190 345256 6196
rect 345676 3126 345704 331214
rect 346596 5302 346624 340068
rect 347056 337890 347084 340068
rect 347044 337884 347096 337890
rect 347044 337826 347096 337832
rect 347516 328574 347544 340068
rect 347976 340054 348082 340082
rect 347504 328568 347556 328574
rect 347504 328510 347556 328516
rect 347976 5370 348004 340054
rect 348424 337884 348476 337890
rect 348424 337826 348476 337832
rect 347964 5364 348016 5370
rect 347964 5306 348016 5312
rect 346584 5296 346636 5302
rect 346584 5238 346636 5244
rect 347872 4140 347924 4146
rect 347872 4082 347924 4088
rect 345664 3120 345716 3126
rect 345664 3062 345716 3068
rect 346676 3120 346728 3126
rect 346676 3062 346728 3068
rect 344376 2984 344428 2990
rect 344376 2926 344428 2932
rect 345480 2984 345532 2990
rect 345480 2926 345532 2932
rect 344560 2916 344612 2922
rect 344560 2858 344612 2864
rect 343640 2848 343692 2854
rect 344572 2802 344600 2858
rect 343640 2790 343692 2796
rect 344296 2774 344600 2802
rect 344296 480 344324 2774
rect 345492 480 345520 2926
rect 346688 480 346716 3062
rect 347884 480 347912 4082
rect 348436 3330 348464 337826
rect 348528 337754 348556 340068
rect 348516 337748 348568 337754
rect 348516 337690 348568 337696
rect 348988 337210 349016 340068
rect 349356 340054 349554 340082
rect 349068 337476 349120 337482
rect 349068 337418 349120 337424
rect 348976 337204 349028 337210
rect 348976 337146 349028 337152
rect 349080 4146 349108 337418
rect 349356 5438 349384 340054
rect 350000 337686 350028 340068
rect 350184 340054 350474 340082
rect 350644 340054 351026 340082
rect 349988 337680 350040 337686
rect 349988 337622 350040 337628
rect 350184 337618 350212 340054
rect 350172 337612 350224 337618
rect 350172 337554 350224 337560
rect 350644 6322 350672 340054
rect 351184 337612 351236 337618
rect 351184 337554 351236 337560
rect 350632 6316 350684 6322
rect 350632 6258 350684 6264
rect 349344 5432 349396 5438
rect 349344 5374 349396 5380
rect 349068 4140 349120 4146
rect 349068 4082 349120 4088
rect 350632 4072 350684 4078
rect 350632 4014 350684 4020
rect 350540 4004 350592 4010
rect 350540 3946 350592 3952
rect 350552 3482 350580 3946
rect 350644 3913 350672 4014
rect 350630 3904 350686 3913
rect 350630 3839 350686 3848
rect 350552 3454 350672 3482
rect 350540 3392 350592 3398
rect 350540 3334 350592 3340
rect 348424 3324 348476 3330
rect 348424 3266 348476 3272
rect 348976 3324 349028 3330
rect 348976 3266 349028 3272
rect 348988 1714 349016 3266
rect 350264 3256 350316 3262
rect 350264 3198 350316 3204
rect 348988 1686 349108 1714
rect 349080 480 349108 1686
rect 350276 480 350304 3198
rect 350552 3194 350580 3334
rect 350644 3194 350672 3454
rect 350540 3188 350592 3194
rect 350540 3130 350592 3136
rect 350632 3188 350684 3194
rect 350632 3130 350684 3136
rect 351196 2990 351224 337554
rect 351472 336802 351500 340068
rect 351932 337822 351960 340068
rect 352116 340054 352498 340082
rect 351920 337816 351972 337822
rect 351920 337758 351972 337764
rect 351828 337544 351880 337550
rect 351828 337486 351880 337492
rect 351460 336796 351512 336802
rect 351460 336738 351512 336744
rect 351840 4146 351868 337486
rect 352116 5506 352144 340054
rect 352944 337958 352972 340068
rect 352932 337952 352984 337958
rect 352932 337894 352984 337900
rect 353404 337006 353432 340068
rect 353496 340054 353970 340082
rect 353392 337000 353444 337006
rect 353392 336942 353444 336948
rect 352564 336796 352616 336802
rect 352564 336738 352616 336744
rect 352104 5500 352156 5506
rect 352104 5442 352156 5448
rect 352576 4486 352604 336738
rect 353496 4554 353524 340054
rect 354416 338094 354444 340068
rect 354404 338088 354456 338094
rect 354404 338030 354456 338036
rect 354876 337686 354904 340068
rect 354968 340054 355442 340082
rect 354864 337680 354916 337686
rect 354864 337622 354916 337628
rect 353484 4548 353536 4554
rect 353484 4490 353536 4496
rect 352564 4480 352616 4486
rect 352564 4422 352616 4428
rect 354968 4350 354996 340054
rect 355888 338026 355916 340068
rect 356256 340054 356362 340082
rect 356624 340054 356914 340082
rect 355876 338020 355928 338026
rect 355876 337962 355928 337968
rect 355324 337952 355376 337958
rect 355324 337894 355376 337900
rect 355336 4418 355364 337894
rect 355968 337136 356020 337142
rect 355968 337078 356020 337084
rect 355324 4412 355376 4418
rect 355324 4354 355376 4360
rect 354956 4344 355008 4350
rect 354956 4286 355008 4292
rect 351368 4140 351420 4146
rect 351368 4082 351420 4088
rect 351828 4140 351880 4146
rect 351828 4082 351880 4088
rect 352564 4140 352616 4146
rect 352564 4082 352616 4088
rect 351184 2984 351236 2990
rect 351184 2926 351236 2932
rect 351380 480 351408 4082
rect 352576 480 352604 4082
rect 354126 4040 354182 4049
rect 354126 3975 354182 3984
rect 354140 3942 354168 3975
rect 354128 3936 354180 3942
rect 354220 3936 354272 3942
rect 354128 3878 354180 3884
rect 354218 3904 354220 3913
rect 354272 3904 354274 3913
rect 354218 3839 354274 3848
rect 353668 3392 353720 3398
rect 353668 3334 353720 3340
rect 353760 3392 353812 3398
rect 353760 3334 353812 3340
rect 353680 3097 353708 3334
rect 353666 3088 353722 3097
rect 353666 3023 353722 3032
rect 353772 480 353800 3334
rect 355980 2990 356008 337078
rect 356152 335640 356204 335646
rect 356152 335582 356204 335588
rect 356164 4282 356192 335582
rect 356152 4276 356204 4282
rect 356152 4218 356204 4224
rect 356256 3369 356284 340054
rect 356624 335646 356652 340054
rect 356704 337680 356756 337686
rect 356704 337622 356756 337628
rect 356612 335640 356664 335646
rect 356612 335582 356664 335588
rect 356242 3360 356298 3369
rect 356242 3295 356298 3304
rect 356716 2990 356744 337622
rect 357360 336870 357388 340068
rect 357348 336864 357400 336870
rect 357348 336806 357400 336812
rect 357820 336802 357848 340068
rect 358004 340054 358386 340082
rect 358846 340054 358952 340082
rect 357808 336796 357860 336802
rect 357808 336738 357860 336744
rect 358004 331906 358032 340054
rect 358084 338088 358136 338094
rect 358084 338030 358136 338036
rect 357348 331900 357400 331906
rect 357348 331842 357400 331848
rect 357992 331900 358044 331906
rect 357992 331842 358044 331848
rect 357360 327162 357388 331842
rect 357360 327134 357480 327162
rect 357452 327078 357480 327134
rect 357440 327072 357492 327078
rect 357440 327014 357492 327020
rect 357532 317484 357584 317490
rect 357532 317426 357584 317432
rect 357544 311930 357572 317426
rect 357544 311902 357848 311930
rect 357820 309126 357848 311902
rect 357808 309120 357860 309126
rect 357808 309062 357860 309068
rect 357900 299532 357952 299538
rect 357900 299474 357952 299480
rect 357912 292602 357940 299474
rect 357440 292596 357492 292602
rect 357440 292538 357492 292544
rect 357900 292596 357952 292602
rect 357900 292538 357952 292544
rect 357452 289814 357480 292538
rect 357440 289808 357492 289814
rect 357440 289750 357492 289756
rect 357716 280220 357768 280226
rect 357716 280162 357768 280168
rect 357728 273290 357756 280162
rect 357440 273284 357492 273290
rect 357440 273226 357492 273232
rect 357716 273284 357768 273290
rect 357716 273226 357768 273232
rect 357452 263616 357480 273226
rect 357452 263588 357664 263616
rect 357636 263514 357664 263588
rect 357544 263486 357664 263514
rect 357544 259418 357572 263486
rect 357532 259412 357584 259418
rect 357532 259354 357584 259360
rect 357716 249824 357768 249830
rect 357716 249766 357768 249772
rect 357728 244202 357756 249766
rect 357636 244174 357756 244202
rect 357636 241482 357664 244174
rect 357636 241454 357756 241482
rect 357728 224890 357756 241454
rect 357636 224862 357756 224890
rect 357636 220833 357664 224862
rect 357438 220824 357494 220833
rect 357438 220759 357494 220768
rect 357622 220824 357678 220833
rect 357622 220759 357678 220768
rect 357452 211177 357480 220759
rect 357438 211168 357494 211177
rect 357438 211103 357494 211112
rect 357714 211168 357770 211177
rect 357714 211103 357770 211112
rect 357728 205578 357756 211103
rect 357636 205550 357756 205578
rect 357636 196058 357664 205550
rect 357544 196030 357664 196058
rect 357544 195974 357572 196030
rect 357532 195968 357584 195974
rect 357532 195910 357584 195916
rect 357716 195968 357768 195974
rect 357716 195910 357768 195916
rect 357728 193225 357756 195910
rect 357714 193216 357770 193225
rect 357714 193151 357770 193160
rect 357898 193216 357954 193225
rect 357898 193151 357954 193160
rect 357912 173942 357940 193151
rect 357624 173936 357676 173942
rect 357624 173878 357676 173884
rect 357900 173936 357952 173942
rect 357900 173878 357952 173884
rect 357636 164393 357664 173878
rect 357622 164384 357678 164393
rect 357622 164319 357678 164328
rect 357530 164248 357586 164257
rect 357530 164183 357586 164192
rect 357544 162858 357572 164183
rect 357532 162852 357584 162858
rect 357532 162794 357584 162800
rect 357808 162852 357860 162858
rect 357808 162794 357860 162800
rect 357820 144974 357848 162794
rect 357532 144968 357584 144974
rect 357532 144910 357584 144916
rect 357808 144968 357860 144974
rect 357808 144910 357860 144916
rect 357544 143546 357572 144910
rect 357256 143540 357308 143546
rect 357256 143482 357308 143488
rect 357532 143540 357584 143546
rect 357532 143482 357584 143488
rect 357268 133929 357296 143482
rect 357254 133920 357310 133929
rect 357254 133855 357310 133864
rect 357438 133920 357494 133929
rect 357438 133855 357494 133864
rect 357452 130370 357480 133855
rect 357452 130342 357572 130370
rect 357544 118794 357572 130342
rect 357532 118788 357584 118794
rect 357532 118730 357584 118736
rect 357440 118652 357492 118658
rect 357440 118594 357492 118600
rect 357452 111058 357480 118594
rect 357452 111030 357572 111058
rect 357544 106282 357572 111030
rect 357532 106276 357584 106282
rect 357532 106218 357584 106224
rect 357624 106276 357676 106282
rect 357624 106218 357676 106224
rect 357636 104854 357664 106218
rect 357624 104848 357676 104854
rect 357624 104790 357676 104796
rect 357624 95260 357676 95266
rect 357624 95202 357676 95208
rect 357636 89842 357664 95202
rect 357636 89814 357756 89842
rect 357728 89706 357756 89814
rect 357544 89678 357756 89706
rect 357544 85542 357572 89678
rect 357532 85536 357584 85542
rect 357532 85478 357584 85484
rect 357624 75948 357676 75954
rect 357624 75890 357676 75896
rect 357636 60738 357664 75890
rect 357636 60710 357756 60738
rect 357728 50946 357756 60710
rect 357636 50918 357756 50946
rect 357636 41426 357664 50918
rect 357636 41398 357756 41426
rect 357728 31770 357756 41398
rect 357544 31742 357756 31770
rect 357544 31634 357572 31742
rect 357544 31606 357664 31634
rect 357636 28966 357664 31606
rect 357624 28960 357676 28966
rect 357624 28902 357676 28908
rect 357808 28960 357860 28966
rect 357808 28902 357860 28908
rect 357820 4214 357848 28902
rect 357808 4208 357860 4214
rect 357808 4150 357860 4156
rect 358096 4078 358124 338030
rect 358728 337816 358780 337822
rect 358728 337758 358780 337764
rect 358740 309126 358768 337758
rect 358728 309120 358780 309126
rect 358728 309062 358780 309068
rect 358728 299532 358780 299538
rect 358728 299474 358780 299480
rect 358740 298110 358768 299474
rect 358728 298104 358780 298110
rect 358728 298046 358780 298052
rect 358728 288448 358780 288454
rect 358728 288390 358780 288396
rect 358740 280362 358768 288390
rect 358728 280356 358780 280362
rect 358728 280298 358780 280304
rect 358728 280220 358780 280226
rect 358728 280162 358780 280168
rect 358740 278769 358768 280162
rect 358542 278760 358598 278769
rect 358542 278695 358598 278704
rect 358726 278760 358782 278769
rect 358726 278695 358782 278704
rect 358556 269142 358584 278695
rect 358544 269136 358596 269142
rect 358544 269078 358596 269084
rect 358728 269136 358780 269142
rect 358728 269078 358780 269084
rect 358740 259457 358768 269078
rect 358542 259448 358598 259457
rect 358542 259383 358598 259392
rect 358726 259448 358782 259457
rect 358726 259383 358782 259392
rect 358556 249830 358584 259383
rect 358544 249824 358596 249830
rect 358544 249766 358596 249772
rect 358728 249824 358780 249830
rect 358728 249766 358780 249772
rect 358740 240145 358768 249766
rect 358542 240136 358598 240145
rect 358542 240071 358598 240080
rect 358726 240136 358782 240145
rect 358726 240071 358782 240080
rect 358556 230518 358584 240071
rect 358544 230512 358596 230518
rect 358544 230454 358596 230460
rect 358728 230512 358780 230518
rect 358728 230454 358780 230460
rect 358740 220833 358768 230454
rect 358542 220824 358598 220833
rect 358542 220759 358598 220768
rect 358726 220824 358782 220833
rect 358726 220759 358782 220768
rect 358556 211177 358584 220759
rect 358542 211168 358598 211177
rect 358542 211103 358598 211112
rect 358726 211168 358782 211177
rect 358726 211103 358782 211112
rect 358740 196602 358768 211103
rect 358740 196574 358860 196602
rect 358832 191826 358860 196574
rect 358544 191820 358596 191826
rect 358544 191762 358596 191768
rect 358820 191820 358872 191826
rect 358820 191762 358872 191768
rect 358556 182209 358584 191762
rect 358542 182200 358598 182209
rect 358542 182135 358598 182144
rect 358726 182200 358782 182209
rect 358726 182135 358782 182144
rect 358740 182034 358768 182135
rect 358728 182028 358780 182034
rect 358728 181970 358780 181976
rect 358820 173868 358872 173874
rect 358820 173810 358872 173816
rect 358832 164286 358860 173810
rect 358728 164280 358780 164286
rect 358728 164222 358780 164228
rect 358820 164280 358872 164286
rect 358820 164222 358872 164228
rect 358740 162858 358768 164222
rect 358728 162852 358780 162858
rect 358728 162794 358780 162800
rect 358728 154556 358780 154562
rect 358728 154498 358780 154504
rect 358740 153218 358768 154498
rect 358740 153190 358860 153218
rect 358832 144974 358860 153190
rect 358728 144968 358780 144974
rect 358728 144910 358780 144916
rect 358820 144968 358872 144974
rect 358820 144910 358872 144916
rect 358740 143546 358768 144910
rect 358728 143540 358780 143546
rect 358728 143482 358780 143488
rect 358728 135244 358780 135250
rect 358728 135186 358780 135192
rect 358740 133906 358768 135186
rect 358740 133878 358860 133906
rect 358832 125662 358860 133878
rect 358728 125656 358780 125662
rect 358728 125598 358780 125604
rect 358820 125656 358872 125662
rect 358820 125598 358872 125604
rect 358740 124166 358768 125598
rect 358728 124160 358780 124166
rect 358728 124102 358780 124108
rect 358728 114572 358780 114578
rect 358728 114514 358780 114520
rect 358740 106593 358768 114514
rect 358726 106584 358782 106593
rect 358726 106519 358782 106528
rect 358726 106312 358782 106321
rect 358726 106247 358782 106256
rect 358740 104854 358768 106247
rect 358728 104848 358780 104854
rect 358728 104790 358780 104796
rect 358820 95260 358872 95266
rect 358820 95202 358872 95208
rect 358832 95146 358860 95202
rect 358648 95118 358860 95146
rect 358648 85610 358676 95118
rect 358544 85604 358596 85610
rect 358544 85546 358596 85552
rect 358636 85604 358688 85610
rect 358636 85546 358688 85552
rect 358556 75954 358584 85546
rect 358544 75948 358596 75954
rect 358544 75890 358596 75896
rect 358728 75948 358780 75954
rect 358728 75890 358780 75896
rect 358740 66178 358768 75890
rect 358740 66150 358860 66178
rect 358832 56642 358860 66150
rect 358728 56636 358780 56642
rect 358728 56578 358780 56584
rect 358820 56636 358872 56642
rect 358820 56578 358872 56584
rect 358740 48346 358768 56578
rect 358728 48340 358780 48346
rect 358728 48282 358780 48288
rect 358728 46980 358780 46986
rect 358728 46922 358780 46928
rect 358740 46866 358768 46922
rect 358740 46838 358860 46866
rect 358832 37330 358860 46838
rect 358728 37324 358780 37330
rect 358728 37266 358780 37272
rect 358820 37324 358872 37330
rect 358820 37266 358872 37272
rect 358740 27690 358768 37266
rect 358648 27662 358768 27690
rect 358648 27606 358676 27662
rect 358636 27600 358688 27606
rect 358636 27542 358688 27548
rect 358544 9716 358596 9722
rect 358544 9658 358596 9664
rect 357440 4072 357492 4078
rect 357440 4014 357492 4020
rect 358084 4072 358136 4078
rect 358176 4072 358228 4078
rect 358084 4014 358136 4020
rect 358174 4040 358176 4049
rect 358228 4040 358230 4049
rect 357452 3346 357480 4014
rect 358174 3975 358230 3984
rect 357268 3318 357480 3346
rect 357268 3262 357296 3318
rect 357256 3256 357308 3262
rect 357256 3198 357308 3204
rect 357348 3256 357400 3262
rect 357348 3198 357400 3204
rect 356794 3088 356850 3097
rect 356794 3023 356850 3032
rect 356808 2990 356836 3023
rect 354956 2984 355008 2990
rect 354956 2926 355008 2932
rect 355968 2984 356020 2990
rect 355968 2926 356020 2932
rect 356060 2984 356112 2990
rect 356060 2926 356112 2932
rect 356704 2984 356756 2990
rect 356704 2926 356756 2932
rect 356796 2984 356848 2990
rect 356796 2926 356848 2932
rect 354968 480 354996 2926
rect 356072 2854 356100 2926
rect 356060 2848 356112 2854
rect 356060 2790 356112 2796
rect 356152 2848 356204 2854
rect 356152 2790 356204 2796
rect 356164 480 356192 2790
rect 357360 480 357388 3198
rect 358556 480 358584 9658
rect 358924 3194 358952 340054
rect 359108 340054 359306 340082
rect 359384 340054 359766 340082
rect 359004 335640 359056 335646
rect 359004 335582 359056 335588
rect 359016 4758 359044 335582
rect 359004 4752 359056 4758
rect 359004 4694 359056 4700
rect 359108 3942 359136 340054
rect 359384 335646 359412 340054
rect 359464 337204 359516 337210
rect 359464 337146 359516 337152
rect 359372 335640 359424 335646
rect 359372 335582 359424 335588
rect 359096 3936 359148 3942
rect 359096 3878 359148 3884
rect 358912 3188 358964 3194
rect 358912 3130 358964 3136
rect 359476 2990 359504 337146
rect 360304 336938 360332 340068
rect 360764 337686 360792 340068
rect 360948 340054 361238 340082
rect 360752 337680 360804 337686
rect 360752 337622 360804 337628
rect 360292 336932 360344 336938
rect 360292 336874 360344 336880
rect 360948 327321 360976 340054
rect 361776 337346 361804 340068
rect 361868 340054 362250 340082
rect 362328 340054 362710 340082
rect 363156 340054 363262 340082
rect 361764 337340 361816 337346
rect 361764 337282 361816 337288
rect 361672 333328 361724 333334
rect 361672 333270 361724 333276
rect 360934 327312 360990 327321
rect 360934 327247 360990 327256
rect 360474 327176 360530 327185
rect 360474 327111 360530 327120
rect 360488 327078 360516 327111
rect 360476 327072 360528 327078
rect 360476 327014 360528 327020
rect 360384 317484 360436 317490
rect 360384 317426 360436 317432
rect 360396 311930 360424 317426
rect 360304 311902 360424 311930
rect 360304 311794 360332 311902
rect 360304 311766 360424 311794
rect 360396 302274 360424 311766
rect 360396 302246 360516 302274
rect 360488 282946 360516 302246
rect 360292 282940 360344 282946
rect 360292 282882 360344 282888
rect 360476 282940 360528 282946
rect 360476 282882 360528 282888
rect 360304 282826 360332 282882
rect 360304 282798 360424 282826
rect 360396 273306 360424 282798
rect 360396 273278 360516 273306
rect 360488 263634 360516 273278
rect 360292 263628 360344 263634
rect 360292 263570 360344 263576
rect 360476 263628 360528 263634
rect 360476 263570 360528 263576
rect 360304 263514 360332 263570
rect 360304 263486 360424 263514
rect 360396 253994 360424 263486
rect 360396 253966 360516 253994
rect 360488 244322 360516 253966
rect 360292 244316 360344 244322
rect 360292 244258 360344 244264
rect 360476 244316 360528 244322
rect 360476 244258 360528 244264
rect 360304 244202 360332 244258
rect 360304 244174 360424 244202
rect 360396 234682 360424 244174
rect 360396 234654 360516 234682
rect 360488 225010 360516 234654
rect 360292 225004 360344 225010
rect 360292 224946 360344 224952
rect 360476 225004 360528 225010
rect 360476 224946 360528 224952
rect 360304 224890 360332 224946
rect 360304 224862 360424 224890
rect 360396 215370 360424 224862
rect 360396 215342 360516 215370
rect 360488 205698 360516 215342
rect 360292 205692 360344 205698
rect 360292 205634 360344 205640
rect 360476 205692 360528 205698
rect 360476 205634 360528 205640
rect 360304 205578 360332 205634
rect 360304 205550 360424 205578
rect 360396 196058 360424 205550
rect 360396 196030 360516 196058
rect 360488 173942 360516 196030
rect 360476 173936 360528 173942
rect 360476 173878 360528 173884
rect 360568 173936 360620 173942
rect 360568 173878 360620 173884
rect 360580 166954 360608 173878
rect 360396 166926 360608 166954
rect 360106 157584 360162 157593
rect 360290 157584 360346 157593
rect 360162 157542 360290 157570
rect 360106 157519 360162 157528
rect 360290 157519 360346 157528
rect 360396 157434 360424 166926
rect 360304 157406 360424 157434
rect 360304 157298 360332 157406
rect 360304 157270 360424 157298
rect 360396 144922 360424 157270
rect 360304 144894 360424 144922
rect 360304 143546 360332 144894
rect 360292 143540 360344 143546
rect 360292 143482 360344 143488
rect 360384 137964 360436 137970
rect 360384 137906 360436 137912
rect 360396 118726 360424 137906
rect 360384 118720 360436 118726
rect 360384 118662 360436 118668
rect 360476 118652 360528 118658
rect 360476 118594 360528 118600
rect 360488 106298 360516 118594
rect 360396 106270 360516 106298
rect 360396 96801 360424 106270
rect 360382 96792 360438 96801
rect 360382 96727 360438 96736
rect 360290 96656 360346 96665
rect 360290 96591 360292 96600
rect 360344 96591 360346 96600
rect 360384 96620 360436 96626
rect 360292 96562 360344 96568
rect 360384 96562 360436 96568
rect 360396 86970 360424 96562
rect 360384 86964 360436 86970
rect 360384 86906 360436 86912
rect 360200 77308 360252 77314
rect 360200 77250 360252 77256
rect 360212 72434 360240 77250
rect 360212 72406 360332 72434
rect 360198 63880 360254 63889
rect 360198 63815 360254 63824
rect 360106 63744 360162 63753
rect 360212 63730 360240 63815
rect 360162 63702 360240 63730
rect 360106 63679 360162 63688
rect 360304 60722 360332 72406
rect 360292 60716 360344 60722
rect 360292 60658 360344 60664
rect 360476 60716 360528 60722
rect 360476 60658 360528 60664
rect 360488 57934 360516 60658
rect 360384 57928 360436 57934
rect 360384 57870 360436 57876
rect 360476 57928 360528 57934
rect 360476 57870 360528 57876
rect 360396 41426 360424 57870
rect 360304 41410 360424 41426
rect 360292 41404 360424 41410
rect 360344 41398 360424 41404
rect 360476 41404 360528 41410
rect 360292 41346 360344 41352
rect 360476 41346 360528 41352
rect 360106 40216 360162 40225
rect 360290 40216 360346 40225
rect 360162 40174 360290 40202
rect 360106 40151 360162 40160
rect 360290 40151 360346 40160
rect 360488 31822 360516 41346
rect 360476 31816 360528 31822
rect 360476 31758 360528 31764
rect 360292 31748 360344 31754
rect 360292 31690 360344 31696
rect 360304 28914 360332 31690
rect 360304 28886 360424 28914
rect 360396 12458 360424 28886
rect 360396 12430 360516 12458
rect 360488 4690 360516 12430
rect 361684 4894 361712 333270
rect 361672 4888 361724 4894
rect 361672 4830 361724 4836
rect 360476 4684 360528 4690
rect 360476 4626 360528 4632
rect 360936 4140 360988 4146
rect 360936 4082 360988 4088
rect 359740 3936 359792 3942
rect 359740 3878 359792 3884
rect 359464 2984 359516 2990
rect 359464 2926 359516 2932
rect 359752 480 359780 3878
rect 360948 480 360976 4082
rect 361868 3466 361896 340054
rect 362224 336864 362276 336870
rect 362224 336806 362276 336812
rect 362236 4078 362264 336806
rect 362328 333334 362356 340054
rect 362868 337816 362920 337822
rect 362868 337758 362920 337764
rect 362316 333328 362368 333334
rect 362316 333270 362368 333276
rect 362224 4072 362276 4078
rect 362224 4014 362276 4020
rect 361856 3460 361908 3466
rect 361856 3402 361908 3408
rect 362880 3330 362908 337758
rect 363052 335640 363104 335646
rect 363052 335582 363104 335588
rect 363064 4826 363092 335582
rect 363052 4820 363104 4826
rect 363052 4762 363104 4768
rect 363156 3534 363184 340054
rect 363708 337210 363736 340068
rect 363800 340054 364182 340082
rect 363696 337204 363748 337210
rect 363696 337146 363748 337152
rect 363604 336796 363656 336802
rect 363604 336738 363656 336744
rect 363328 4140 363380 4146
rect 363328 4082 363380 4088
rect 363144 3528 363196 3534
rect 363144 3470 363196 3476
rect 362132 3324 362184 3330
rect 362132 3266 362184 3272
rect 362868 3324 362920 3330
rect 362868 3266 362920 3272
rect 362144 480 362172 3266
rect 363340 480 363368 4082
rect 363616 3602 363644 336738
rect 363800 335646 363828 340054
rect 364248 338020 364300 338026
rect 364248 337962 364300 337968
rect 363788 335640 363840 335646
rect 363788 335582 363840 335588
rect 364260 4146 364288 337962
rect 364720 336802 364748 340068
rect 365180 336870 365208 340068
rect 365640 337890 365668 340068
rect 365824 340054 366206 340082
rect 365628 337884 365680 337890
rect 365628 337826 365680 337832
rect 365168 336864 365220 336870
rect 365168 336806 365220 336812
rect 364708 336796 364760 336802
rect 364708 336738 364760 336744
rect 364248 4140 364300 4146
rect 364248 4082 364300 4088
rect 365824 3670 365852 340054
rect 366652 337210 366680 340068
rect 367126 340054 367232 340082
rect 366916 337612 366968 337618
rect 366916 337554 366968 337560
rect 366640 337204 366692 337210
rect 366640 337146 366692 337152
rect 366822 183560 366878 183569
rect 366822 183495 366878 183504
rect 366836 174010 366864 183495
rect 366928 174078 366956 337554
rect 367008 337340 367060 337346
rect 367008 337282 367060 337288
rect 367020 241505 367048 337282
rect 367006 241496 367062 241505
rect 367006 241431 367062 241440
rect 367006 231976 367062 231985
rect 367006 231911 367062 231920
rect 367020 193186 367048 231911
rect 367008 193180 367060 193186
rect 367008 193122 367060 193128
rect 367008 183592 367060 183598
rect 367006 183560 367008 183569
rect 367060 183560 367062 183569
rect 367006 183495 367062 183504
rect 366916 174072 366968 174078
rect 366916 174014 366968 174020
rect 366824 174004 366876 174010
rect 366824 173946 366876 173952
rect 367008 174004 367060 174010
rect 367008 173946 367060 173952
rect 366916 173936 366968 173942
rect 367020 173913 367048 173946
rect 366916 173878 366968 173884
rect 367006 173904 367062 173913
rect 366928 19310 366956 173878
rect 367006 173839 367062 173848
rect 367006 164248 367062 164257
rect 367006 164183 367062 164192
rect 367020 154562 367048 164183
rect 367008 154556 367060 154562
rect 367008 154498 367060 154504
rect 367008 144968 367060 144974
rect 367008 144910 367060 144916
rect 367020 125594 367048 144910
rect 367008 125588 367060 125594
rect 367008 125530 367060 125536
rect 367008 116068 367060 116074
rect 367008 116010 367060 116016
rect 367020 115938 367048 116010
rect 367008 115932 367060 115938
rect 367008 115874 367060 115880
rect 367008 106344 367060 106350
rect 367008 106286 367060 106292
rect 367020 96801 367048 106286
rect 367006 96792 367062 96801
rect 367006 96727 367062 96736
rect 367006 96656 367062 96665
rect 367006 96591 367008 96600
rect 367060 96591 367062 96600
rect 367008 96562 367060 96568
rect 367008 87032 367060 87038
rect 367008 86974 367060 86980
rect 367020 77450 367048 86974
rect 367008 77444 367060 77450
rect 367008 77386 367060 77392
rect 367008 77308 367060 77314
rect 367008 77250 367060 77256
rect 367020 57934 367048 77250
rect 367008 57928 367060 57934
rect 367008 57870 367060 57876
rect 367008 48340 367060 48346
rect 367008 48282 367060 48288
rect 367020 38622 367048 48282
rect 367008 38616 367060 38622
rect 367008 38558 367060 38564
rect 367008 29096 367060 29102
rect 367100 29096 367152 29102
rect 367008 29038 367060 29044
rect 367098 29064 367100 29073
rect 367152 29064 367154 29073
rect 367020 28966 367048 29038
rect 367098 28999 367154 29008
rect 367008 28960 367060 28966
rect 367008 28902 367060 28908
rect 367008 19372 367060 19378
rect 367008 19314 367060 19320
rect 366916 19304 366968 19310
rect 366916 19246 366968 19252
rect 367020 19242 367048 19314
rect 366824 19236 366876 19242
rect 366824 19178 366876 19184
rect 367008 19236 367060 19242
rect 367008 19178 367060 19184
rect 365812 3664 365864 3670
rect 365812 3606 365864 3612
rect 363604 3596 363656 3602
rect 363604 3538 363656 3544
rect 365720 3596 365772 3602
rect 365720 3538 365772 3544
rect 364524 3324 364576 3330
rect 364524 3266 364576 3272
rect 364536 480 364564 3266
rect 365732 480 365760 3538
rect 366836 2938 366864 19178
rect 366916 12368 366968 12374
rect 366916 12310 366968 12316
rect 366928 3602 366956 12310
rect 367204 4962 367232 340054
rect 367664 337074 367692 340068
rect 367940 340054 368138 340082
rect 367652 337068 367704 337074
rect 367652 337010 367704 337016
rect 367940 335646 367968 340054
rect 367284 335640 367336 335646
rect 367284 335582 367336 335588
rect 367928 335640 367980 335646
rect 367928 335582 367980 335588
rect 367192 4956 367244 4962
rect 367192 4898 367244 4904
rect 366916 3596 366968 3602
rect 366916 3538 366968 3544
rect 367296 3194 367324 335582
rect 368584 5098 368612 340068
rect 368676 340054 369150 340082
rect 368572 5092 368624 5098
rect 368572 5034 368624 5040
rect 368676 3806 368704 340054
rect 369596 337754 369624 340068
rect 370056 337958 370084 340068
rect 370148 340054 370622 340082
rect 370044 337952 370096 337958
rect 370044 337894 370096 337900
rect 369584 337748 369636 337754
rect 369584 337690 369636 337696
rect 369768 337408 369820 337414
rect 369768 337350 369820 337356
rect 369124 337136 369176 337142
rect 369124 337078 369176 337084
rect 368664 3800 368716 3806
rect 368664 3742 368716 3748
rect 369136 3534 369164 337078
rect 369780 4146 369808 337350
rect 369216 4140 369268 4146
rect 369216 4082 369268 4088
rect 369768 4140 369820 4146
rect 369768 4082 369820 4088
rect 369124 3528 369176 3534
rect 369124 3470 369176 3476
rect 368020 3460 368072 3466
rect 368020 3402 368072 3408
rect 367284 3188 367336 3194
rect 367284 3130 367336 3136
rect 366836 2910 366956 2938
rect 366928 480 366956 2910
rect 368032 480 368060 3402
rect 369228 480 369256 4082
rect 370148 3874 370176 340054
rect 371068 337142 371096 340068
rect 371528 338094 371556 340068
rect 371516 338088 371568 338094
rect 371516 338030 371568 338036
rect 371148 337952 371200 337958
rect 371148 337894 371200 337900
rect 371056 337136 371108 337142
rect 371056 337078 371108 337084
rect 370504 336796 370556 336802
rect 370504 336738 370556 336744
rect 370412 4140 370464 4146
rect 370412 4082 370464 4088
rect 370136 3868 370188 3874
rect 370136 3810 370188 3816
rect 370424 480 370452 4082
rect 370516 3126 370544 336738
rect 371160 4146 371188 337894
rect 372080 337482 372108 340068
rect 372068 337476 372120 337482
rect 372068 337418 372120 337424
rect 372540 336802 372568 340068
rect 373000 337278 373028 340068
rect 373276 340054 373566 340082
rect 374026 340054 374132 340082
rect 372988 337272 373040 337278
rect 372988 337214 373040 337220
rect 372528 336796 372580 336802
rect 372528 336738 372580 336744
rect 373276 328506 373304 340054
rect 373908 337544 373960 337550
rect 373908 337486 373960 337492
rect 372712 328500 372764 328506
rect 372712 328442 372764 328448
rect 373264 328500 373316 328506
rect 373264 328442 373316 328448
rect 372724 311930 372752 328442
rect 372632 311902 372752 311930
rect 372632 311794 372660 311902
rect 372632 311766 372752 311794
rect 372724 299470 372752 311766
rect 372712 299464 372764 299470
rect 372712 299406 372764 299412
rect 372712 289876 372764 289882
rect 372712 289818 372764 289824
rect 372724 280158 372752 289818
rect 372712 280152 372764 280158
rect 372712 280094 372764 280100
rect 372712 270564 372764 270570
rect 372712 270506 372764 270512
rect 372724 260846 372752 270506
rect 372712 260840 372764 260846
rect 372712 260782 372764 260788
rect 372712 251252 372764 251258
rect 372712 251194 372764 251200
rect 372724 241505 372752 251194
rect 372526 241496 372582 241505
rect 372526 241431 372582 241440
rect 372710 241496 372766 241505
rect 372710 241431 372766 241440
rect 372540 231878 372568 241431
rect 372528 231872 372580 231878
rect 372528 231814 372580 231820
rect 372712 231872 372764 231878
rect 372712 231814 372764 231820
rect 372724 222193 372752 231814
rect 372526 222184 372582 222193
rect 372526 222119 372582 222128
rect 372710 222184 372766 222193
rect 372710 222119 372766 222128
rect 372540 212566 372568 222119
rect 372528 212560 372580 212566
rect 372528 212502 372580 212508
rect 372712 212560 372764 212566
rect 372712 212502 372764 212508
rect 372724 202881 372752 212502
rect 372526 202872 372582 202881
rect 372526 202807 372582 202816
rect 372710 202872 372766 202881
rect 372710 202807 372766 202816
rect 372540 193254 372568 202807
rect 372528 193248 372580 193254
rect 372528 193190 372580 193196
rect 372712 193248 372764 193254
rect 372712 193190 372764 193196
rect 372724 183569 372752 193190
rect 372526 183560 372582 183569
rect 372526 183495 372582 183504
rect 372710 183560 372766 183569
rect 372710 183495 372766 183504
rect 372540 173942 372568 183495
rect 372528 173936 372580 173942
rect 372528 173878 372580 173884
rect 372804 173936 372856 173942
rect 372804 173878 372856 173884
rect 372816 164218 372844 173878
rect 372804 164212 372856 164218
rect 372804 164154 372856 164160
rect 372804 159316 372856 159322
rect 372804 159258 372856 159264
rect 372816 138174 372844 159258
rect 372804 138168 372856 138174
rect 372804 138110 372856 138116
rect 372712 135312 372764 135318
rect 372712 135254 372764 135260
rect 372724 125594 372752 135254
rect 372712 125588 372764 125594
rect 372712 125530 372764 125536
rect 372712 116000 372764 116006
rect 372712 115942 372764 115948
rect 372724 99498 372752 115942
rect 372632 99470 372752 99498
rect 372632 99362 372660 99470
rect 372632 99334 372752 99362
rect 372724 91746 372752 99334
rect 372540 91718 372752 91746
rect 372540 86986 372568 91718
rect 372448 86958 372568 86986
rect 372448 79966 372476 86958
rect 372436 79960 372488 79966
rect 372436 79902 372488 79908
rect 372804 79960 372856 79966
rect 372804 79902 372856 79908
rect 372816 75886 372844 79902
rect 372804 75880 372856 75886
rect 372804 75822 372856 75828
rect 372712 66292 372764 66298
rect 372712 66234 372764 66240
rect 372724 51082 372752 66234
rect 372632 51054 372752 51082
rect 372632 50946 372660 51054
rect 372632 50918 372752 50946
rect 372724 31890 372752 50918
rect 372712 31884 372764 31890
rect 372712 31826 372764 31832
rect 372712 29028 372764 29034
rect 372712 28970 372764 28976
rect 372724 22098 372752 28970
rect 372712 22092 372764 22098
rect 372712 22034 372764 22040
rect 372804 22024 372856 22030
rect 372804 21966 372856 21972
rect 371148 4140 371200 4146
rect 371148 4082 371200 4088
rect 372816 4026 372844 21966
rect 372724 3998 372844 4026
rect 372724 3738 372752 3998
rect 373920 3874 373948 337486
rect 374104 3942 374132 340054
rect 374472 337482 374500 340068
rect 374460 337476 374512 337482
rect 374460 337418 374512 337424
rect 374564 336734 374592 340190
rect 375498 340054 375696 340082
rect 375288 337544 375340 337550
rect 375288 337486 375340 337492
rect 374552 336728 374604 336734
rect 374552 336670 374604 336676
rect 374460 327140 374512 327146
rect 374460 327082 374512 327088
rect 374472 318850 374500 327082
rect 374368 318844 374420 318850
rect 374368 318786 374420 318792
rect 374460 318844 374512 318850
rect 374460 318786 374512 318792
rect 374380 311982 374408 318786
rect 374368 311976 374420 311982
rect 374368 311918 374420 311924
rect 374460 311772 374512 311778
rect 374460 311714 374512 311720
rect 374472 307766 374500 311714
rect 374460 307760 374512 307766
rect 374460 307702 374512 307708
rect 374368 289876 374420 289882
rect 374368 289818 374420 289824
rect 374380 273222 374408 289818
rect 374368 273216 374420 273222
rect 374368 273158 374420 273164
rect 374368 273080 374420 273086
rect 374368 273022 374420 273028
rect 374380 253910 374408 273022
rect 374368 253904 374420 253910
rect 374368 253846 374420 253852
rect 374368 253768 374420 253774
rect 374368 253710 374420 253716
rect 374380 234598 374408 253710
rect 374368 234592 374420 234598
rect 374368 234534 374420 234540
rect 374368 234456 374420 234462
rect 374368 234398 374420 234404
rect 374380 215286 374408 234398
rect 374368 215280 374420 215286
rect 374368 215222 374420 215228
rect 374368 215144 374420 215150
rect 374368 215086 374420 215092
rect 374380 195974 374408 215086
rect 374368 195968 374420 195974
rect 374368 195910 374420 195916
rect 374368 195832 374420 195838
rect 374368 195774 374420 195780
rect 374380 176662 374408 195774
rect 374368 176656 374420 176662
rect 374368 176598 374420 176604
rect 374368 176520 374420 176526
rect 374368 176462 374420 176468
rect 374380 157350 374408 176462
rect 374368 157344 374420 157350
rect 374368 157286 374420 157292
rect 374368 157208 374420 157214
rect 374368 157150 374420 157156
rect 374380 114753 374408 157150
rect 374366 114744 374422 114753
rect 374366 114679 374422 114688
rect 374274 114608 374330 114617
rect 374330 114566 374408 114594
rect 374274 114543 374330 114552
rect 374380 114510 374408 114566
rect 374368 114504 374420 114510
rect 374368 114446 374420 114452
rect 374368 104984 374420 104990
rect 374368 104926 374420 104932
rect 374380 104854 374408 104926
rect 374368 104848 374420 104854
rect 374368 104790 374420 104796
rect 374368 99340 374420 99346
rect 374368 99282 374420 99288
rect 374380 60738 374408 99282
rect 374288 60710 374408 60738
rect 374288 60602 374316 60710
rect 374288 60574 374408 60602
rect 374380 41426 374408 60574
rect 374288 41398 374408 41426
rect 374288 41290 374316 41398
rect 374288 41262 374408 41290
rect 374380 22166 374408 41262
rect 374368 22160 374420 22166
rect 374368 22102 374420 22108
rect 374368 22024 374420 22030
rect 374368 21966 374420 21972
rect 374092 3936 374144 3942
rect 374092 3878 374144 3884
rect 372804 3868 372856 3874
rect 372804 3810 372856 3816
rect 373908 3868 373960 3874
rect 373908 3810 373960 3816
rect 372712 3732 372764 3738
rect 372712 3674 372764 3680
rect 371608 3596 371660 3602
rect 371608 3538 371660 3544
rect 370504 3120 370556 3126
rect 370504 3062 370556 3068
rect 371620 480 371648 3538
rect 372816 480 372844 3810
rect 374000 3800 374052 3806
rect 374000 3742 374052 3748
rect 374012 480 374040 3742
rect 374380 2990 374408 21966
rect 375300 3806 375328 337486
rect 375288 3800 375340 3806
rect 375288 3742 375340 3748
rect 375196 3664 375248 3670
rect 375196 3606 375248 3612
rect 374368 2984 374420 2990
rect 374368 2926 374420 2932
rect 375208 480 375236 3606
rect 375668 3398 375696 340054
rect 375944 337754 375972 340068
rect 376036 340054 376510 340082
rect 375932 337748 375984 337754
rect 375932 337690 375984 337696
rect 376036 336954 376064 340054
rect 376668 338088 376720 338094
rect 376588 338048 376668 338076
rect 376588 337686 376616 338048
rect 376668 338030 376720 338036
rect 376758 338056 376814 338065
rect 376758 337991 376760 338000
rect 376812 337991 376814 338000
rect 376760 337962 376812 337968
rect 376576 337680 376628 337686
rect 376576 337622 376628 337628
rect 375852 336926 376064 336954
rect 375852 336734 375880 336926
rect 376956 336802 376984 340068
rect 377416 337890 377444 340068
rect 377508 340054 377890 340082
rect 377404 337884 377456 337890
rect 377404 337826 377456 337832
rect 376024 336796 376076 336802
rect 376024 336738 376076 336744
rect 376944 336796 376996 336802
rect 376944 336738 376996 336744
rect 375840 336728 375892 336734
rect 375840 336670 375892 336676
rect 375932 327140 375984 327146
rect 375932 327082 375984 327088
rect 375944 318850 375972 327082
rect 375840 318844 375892 318850
rect 375840 318786 375892 318792
rect 375932 318844 375984 318850
rect 375932 318786 375984 318792
rect 375852 317422 375880 318786
rect 375840 317416 375892 317422
rect 375840 317358 375892 317364
rect 375840 307828 375892 307834
rect 375840 307770 375892 307776
rect 375852 299554 375880 307770
rect 375852 299526 375972 299554
rect 375944 299470 375972 299526
rect 375932 299464 375984 299470
rect 375932 299406 375984 299412
rect 375840 289876 375892 289882
rect 375840 289818 375892 289824
rect 375852 273222 375880 289818
rect 375840 273216 375892 273222
rect 375840 273158 375892 273164
rect 375840 273080 375892 273086
rect 375840 273022 375892 273028
rect 375852 253910 375880 273022
rect 375840 253904 375892 253910
rect 375840 253846 375892 253852
rect 375840 253768 375892 253774
rect 375840 253710 375892 253716
rect 375852 234598 375880 253710
rect 375840 234592 375892 234598
rect 375840 234534 375892 234540
rect 375840 234456 375892 234462
rect 375840 234398 375892 234404
rect 375852 215286 375880 234398
rect 375840 215280 375892 215286
rect 375840 215222 375892 215228
rect 375840 215144 375892 215150
rect 375840 215086 375892 215092
rect 375852 195974 375880 215086
rect 375840 195968 375892 195974
rect 375840 195910 375892 195916
rect 375840 195832 375892 195838
rect 375840 195774 375892 195780
rect 375852 176662 375880 195774
rect 375840 176656 375892 176662
rect 375840 176598 375892 176604
rect 375840 176520 375892 176526
rect 375840 176462 375892 176468
rect 375852 157350 375880 176462
rect 375840 157344 375892 157350
rect 375840 157286 375892 157292
rect 375840 157208 375892 157214
rect 375840 157150 375892 157156
rect 375852 153202 375880 157150
rect 375840 153196 375892 153202
rect 375840 153138 375892 153144
rect 375840 143608 375892 143614
rect 375840 143550 375892 143556
rect 375852 133890 375880 143550
rect 375840 133884 375892 133890
rect 375840 133826 375892 133832
rect 375840 124228 375892 124234
rect 375840 124170 375892 124176
rect 375852 114510 375880 124170
rect 375840 114504 375892 114510
rect 375840 114446 375892 114452
rect 375840 104984 375892 104990
rect 375840 104926 375892 104932
rect 375852 104854 375880 104926
rect 375840 104848 375892 104854
rect 375840 104790 375892 104796
rect 375840 95260 375892 95266
rect 375840 95202 375892 95208
rect 375852 60738 375880 95202
rect 375760 60710 375880 60738
rect 375760 60602 375788 60710
rect 375760 60574 375880 60602
rect 375852 41426 375880 60574
rect 375760 41398 375880 41426
rect 375760 41290 375788 41398
rect 375760 41262 375880 41290
rect 375852 28966 375880 41262
rect 375840 28960 375892 28966
rect 375840 28902 375892 28908
rect 375840 19372 375892 19378
rect 375840 19314 375892 19320
rect 375656 3392 375708 3398
rect 375656 3334 375708 3340
rect 375852 2854 375880 19314
rect 376036 3262 376064 336738
rect 377508 335594 377536 340054
rect 378048 337000 378100 337006
rect 378048 336942 378100 336948
rect 377680 336796 377732 336802
rect 377680 336738 377732 336744
rect 377140 335566 377536 335594
rect 377140 323610 377168 335566
rect 377692 335458 377720 336738
rect 377416 335430 377720 335458
rect 376852 323604 376904 323610
rect 376852 323546 376904 323552
rect 377128 323604 377180 323610
rect 377128 323546 377180 323552
rect 376864 318889 376892 323546
rect 376850 318880 376906 318889
rect 376850 318815 376906 318824
rect 377126 318880 377182 318889
rect 377126 318815 377182 318824
rect 377140 317422 377168 318815
rect 377128 317416 377180 317422
rect 377128 317358 377180 317364
rect 377312 317416 377364 317422
rect 377312 317358 377364 317364
rect 377324 302122 377352 317358
rect 377128 302116 377180 302122
rect 377128 302058 377180 302064
rect 377312 302116 377364 302122
rect 377312 302058 377364 302064
rect 377140 292670 377168 302058
rect 377128 292664 377180 292670
rect 377128 292606 377180 292612
rect 377128 292460 377180 292466
rect 377128 292402 377180 292408
rect 377140 280158 377168 292402
rect 377128 280152 377180 280158
rect 377128 280094 377180 280100
rect 377128 270564 377180 270570
rect 377128 270506 377180 270512
rect 377140 260846 377168 270506
rect 377128 260840 377180 260846
rect 377128 260782 377180 260788
rect 377128 251252 377180 251258
rect 377128 251194 377180 251200
rect 377140 241505 377168 251194
rect 376942 241496 376998 241505
rect 376942 241431 376998 241440
rect 377126 241496 377182 241505
rect 377126 241431 377182 241440
rect 376956 231878 376984 241431
rect 376944 231872 376996 231878
rect 376944 231814 376996 231820
rect 377128 231872 377180 231878
rect 377128 231814 377180 231820
rect 377140 222193 377168 231814
rect 376942 222184 376998 222193
rect 376942 222119 376998 222128
rect 377126 222184 377182 222193
rect 377126 222119 377182 222128
rect 376956 212566 376984 222119
rect 376944 212560 376996 212566
rect 376944 212502 376996 212508
rect 377128 212560 377180 212566
rect 377128 212502 377180 212508
rect 377140 202881 377168 212502
rect 376942 202872 376998 202881
rect 376942 202807 376998 202816
rect 377126 202872 377182 202881
rect 377126 202807 377182 202816
rect 376956 193254 376984 202807
rect 376944 193248 376996 193254
rect 376944 193190 376996 193196
rect 377128 193248 377180 193254
rect 377128 193190 377180 193196
rect 377140 183569 377168 193190
rect 376942 183560 376998 183569
rect 376942 183495 376998 183504
rect 377126 183560 377182 183569
rect 377126 183495 377182 183504
rect 376956 173942 376984 183495
rect 376944 173936 376996 173942
rect 376944 173878 376996 173884
rect 377128 173936 377180 173942
rect 377128 173878 377180 173884
rect 377140 164218 377168 173878
rect 376944 164212 376996 164218
rect 376944 164154 376996 164160
rect 377128 164212 377180 164218
rect 377128 164154 377180 164160
rect 376956 154601 376984 164154
rect 376942 154592 376998 154601
rect 376942 154527 376998 154536
rect 377126 154592 377182 154601
rect 377126 154527 377182 154536
rect 377140 144906 377168 154527
rect 376944 144900 376996 144906
rect 376944 144842 376996 144848
rect 377128 144900 377180 144906
rect 377128 144842 377180 144848
rect 376956 135289 376984 144842
rect 376942 135280 376998 135289
rect 376942 135215 376998 135224
rect 377126 135280 377182 135289
rect 377126 135215 377182 135224
rect 377140 118726 377168 135215
rect 377128 118720 377180 118726
rect 377128 118662 377180 118668
rect 377128 118584 377180 118590
rect 377128 118526 377180 118532
rect 377140 115938 377168 118526
rect 377128 115932 377180 115938
rect 377128 115874 377180 115880
rect 377036 106344 377088 106350
rect 377088 106292 377168 106298
rect 377036 106286 377168 106292
rect 377048 106282 377168 106286
rect 377048 106276 377180 106282
rect 377048 106270 377128 106276
rect 377128 106218 377180 106224
rect 377128 99340 377180 99346
rect 377128 99282 377180 99288
rect 376758 87136 376814 87145
rect 376758 87071 376760 87080
rect 376812 87071 376814 87080
rect 376760 87042 376812 87048
rect 377140 60738 377168 99282
rect 377048 60710 377168 60738
rect 377048 60602 377076 60710
rect 377048 60574 377168 60602
rect 377140 41342 377168 60574
rect 377128 41336 377180 41342
rect 377128 41278 377180 41284
rect 377036 38752 377088 38758
rect 377088 38700 377168 38706
rect 377036 38694 377168 38700
rect 377048 38678 377168 38694
rect 377140 38622 377168 38678
rect 377128 38616 377180 38622
rect 377128 38558 377180 38564
rect 377312 38616 377364 38622
rect 377312 38558 377364 38564
rect 376666 29336 376722 29345
rect 376666 29271 376722 29280
rect 376680 29102 376708 29271
rect 376668 29096 376720 29102
rect 377324 29073 377352 38558
rect 376668 29038 376720 29044
rect 377126 29064 377182 29073
rect 377126 28999 377182 29008
rect 377310 29064 377366 29073
rect 377310 28999 377366 29008
rect 377140 28966 377168 28999
rect 377128 28960 377180 28966
rect 377128 28902 377180 28908
rect 377128 22092 377180 22098
rect 377128 22034 377180 22040
rect 377140 4010 377168 22034
rect 377416 4078 377444 335430
rect 378060 4146 378088 336942
rect 378428 336802 378456 340068
rect 378888 337822 378916 340068
rect 379348 338065 379376 340068
rect 379716 340054 379914 340082
rect 379334 338056 379390 338065
rect 379334 337991 379390 338000
rect 378876 337816 378928 337822
rect 378876 337758 378928 337764
rect 378416 336796 378468 336802
rect 378416 336738 378468 336744
rect 377588 4140 377640 4146
rect 377588 4082 377640 4088
rect 378048 4140 378100 4146
rect 378048 4082 378100 4088
rect 378784 4140 378836 4146
rect 378784 4082 378836 4088
rect 377404 4072 377456 4078
rect 377404 4014 377456 4020
rect 377128 4004 377180 4010
rect 377128 3946 377180 3952
rect 376392 3800 376444 3806
rect 376392 3742 376444 3748
rect 376024 3256 376076 3262
rect 376024 3198 376076 3204
rect 375840 2848 375892 2854
rect 375840 2790 375892 2796
rect 376404 480 376432 3742
rect 377600 480 377628 4082
rect 378796 480 378824 4082
rect 379716 3738 379744 340054
rect 380360 338094 380388 340068
rect 380348 338088 380400 338094
rect 380348 338030 380400 338036
rect 380164 337748 380216 337754
rect 380164 337690 380216 337696
rect 380176 4418 380204 337690
rect 380820 337346 380848 340068
rect 381372 337754 381400 340068
rect 381360 337748 381412 337754
rect 381360 337690 381412 337696
rect 381544 337748 381596 337754
rect 381544 337690 381596 337696
rect 380808 337340 380860 337346
rect 380808 337282 380860 337288
rect 380808 336932 380860 336938
rect 380808 336874 380860 336880
rect 380164 4412 380216 4418
rect 380164 4354 380216 4360
rect 380820 4078 380848 336874
rect 379980 4072 380032 4078
rect 379980 4014 380032 4020
rect 380808 4072 380860 4078
rect 380808 4014 380860 4020
rect 381176 4072 381228 4078
rect 381176 4014 381228 4020
rect 379704 3732 379756 3738
rect 379704 3674 379756 3680
rect 379992 480 380020 4014
rect 381188 480 381216 4014
rect 381556 3602 381584 337690
rect 381832 337482 381860 340068
rect 382292 338026 382320 340068
rect 382280 338020 382332 338026
rect 382280 337962 382332 337968
rect 382844 337754 382872 340068
rect 382832 337748 382884 337754
rect 382832 337690 382884 337696
rect 383304 337618 383332 340068
rect 383292 337612 383344 337618
rect 383292 337554 383344 337560
rect 383764 337550 383792 340068
rect 383856 340054 384330 340082
rect 383752 337544 383804 337550
rect 383752 337486 383804 337492
rect 381820 337476 381872 337482
rect 381820 337418 381872 337424
rect 382188 337408 382240 337414
rect 382188 337350 382240 337356
rect 381636 336864 381688 336870
rect 381636 336806 381688 336812
rect 381648 3806 381676 336806
rect 382200 4078 382228 337350
rect 382188 4072 382240 4078
rect 382188 4014 382240 4020
rect 383568 4072 383620 4078
rect 383568 4014 383620 4020
rect 381636 3800 381688 3806
rect 381636 3742 381688 3748
rect 381544 3596 381596 3602
rect 381544 3538 381596 3544
rect 382372 3460 382424 3466
rect 382372 3402 382424 3408
rect 382384 480 382412 3402
rect 383580 480 383608 4014
rect 383856 3670 383884 340054
rect 384304 337680 384356 337686
rect 384304 337622 384356 337628
rect 384316 4078 384344 337622
rect 384776 336870 384804 340068
rect 384948 337748 385000 337754
rect 384948 337690 385000 337696
rect 384764 336864 384816 336870
rect 384764 336806 384816 336812
rect 384304 4072 384356 4078
rect 384304 4014 384356 4020
rect 383844 3664 383896 3670
rect 383844 3606 383896 3612
rect 384960 610 384988 337690
rect 385236 337006 385264 340068
rect 385328 340054 385802 340082
rect 385224 337000 385276 337006
rect 385224 336942 385276 336948
rect 385328 4146 385356 340054
rect 386248 336938 386276 340068
rect 386708 337414 386736 340068
rect 386696 337408 386748 337414
rect 386696 337350 386748 337356
rect 386800 337226 386828 340190
rect 387720 337686 387748 340068
rect 388180 337754 388208 340068
rect 388444 337816 388496 337822
rect 388444 337758 388496 337764
rect 388168 337748 388220 337754
rect 388168 337690 388220 337696
rect 387708 337680 387760 337686
rect 387708 337622 387760 337628
rect 387064 337476 387116 337482
rect 387064 337418 387116 337424
rect 386616 337198 386828 337226
rect 386236 336932 386288 336938
rect 386236 336874 386288 336880
rect 386236 87100 386288 87106
rect 386236 87042 386288 87048
rect 386420 87100 386472 87106
rect 386420 87042 386472 87048
rect 386248 87009 386276 87042
rect 386432 87009 386460 87042
rect 386234 87000 386290 87009
rect 386234 86935 386290 86944
rect 386418 87000 386474 87009
rect 386418 86935 386474 86944
rect 385316 4140 385368 4146
rect 385316 4082 385368 4088
rect 386616 3466 386644 337198
rect 386604 3460 386656 3466
rect 386604 3402 386656 3408
rect 387076 2922 387104 337418
rect 388260 3528 388312 3534
rect 388260 3470 388312 3476
rect 385868 2916 385920 2922
rect 385868 2858 385920 2864
rect 387064 2916 387116 2922
rect 387064 2858 387116 2864
rect 384672 604 384724 610
rect 384672 546 384724 552
rect 384948 604 385000 610
rect 384948 546 385000 552
rect 384684 480 384712 546
rect 385880 480 385908 2858
rect 387064 2780 387116 2786
rect 387064 2722 387116 2728
rect 387076 480 387104 2722
rect 388272 480 388300 3470
rect 388456 2854 388484 337758
rect 388732 337482 388760 340068
rect 389192 337822 389220 340068
rect 389284 340054 389666 340082
rect 389744 340054 390218 340082
rect 390572 340054 390678 340082
rect 390848 340054 391138 340082
rect 391690 340054 391888 340082
rect 389180 337816 389232 337822
rect 389180 337758 389232 337764
rect 389284 337668 389312 340054
rect 389100 337640 389312 337668
rect 388720 337476 388772 337482
rect 388720 337418 388772 337424
rect 388994 251152 389050 251161
rect 388994 251087 389050 251096
rect 389008 241602 389036 251087
rect 388996 241596 389048 241602
rect 388996 241538 389048 241544
rect 389100 3534 389128 337640
rect 389744 331294 389772 340054
rect 389732 331288 389784 331294
rect 389732 331230 389784 331236
rect 389640 331220 389692 331226
rect 389640 331162 389692 331168
rect 389652 328438 389680 331162
rect 389640 328432 389692 328438
rect 389640 328374 389692 328380
rect 389548 318844 389600 318850
rect 389548 318786 389600 318792
rect 389560 309194 389588 318786
rect 389364 309188 389416 309194
rect 389364 309130 389416 309136
rect 389548 309188 389600 309194
rect 389548 309130 389600 309136
rect 389376 309058 389404 309130
rect 389364 309052 389416 309058
rect 389364 308994 389416 309000
rect 389272 299532 389324 299538
rect 389272 299474 389324 299480
rect 389284 292618 389312 299474
rect 389284 292590 389496 292618
rect 389468 289814 389496 292590
rect 389456 289808 389508 289814
rect 389456 289750 389508 289756
rect 389364 280220 389416 280226
rect 389364 280162 389416 280168
rect 389376 273306 389404 280162
rect 389376 273278 389496 273306
rect 389468 270502 389496 273278
rect 389456 270496 389508 270502
rect 389456 270438 389508 270444
rect 389364 260908 389416 260914
rect 389364 260850 389416 260856
rect 389376 251258 389404 260850
rect 389180 251252 389232 251258
rect 389180 251194 389232 251200
rect 389364 251252 389416 251258
rect 389364 251194 389416 251200
rect 389192 251161 389220 251194
rect 389178 251152 389234 251161
rect 389178 251087 389234 251096
rect 389272 241596 389324 241602
rect 389272 241538 389324 241544
rect 389284 241466 389312 241538
rect 389272 241460 389324 241466
rect 389272 241402 389324 241408
rect 389456 234660 389508 234666
rect 389456 234602 389508 234608
rect 389468 231849 389496 234602
rect 389270 231840 389326 231849
rect 389270 231775 389326 231784
rect 389454 231840 389510 231849
rect 389454 231775 389510 231784
rect 389284 222222 389312 231775
rect 389272 222216 389324 222222
rect 389272 222158 389324 222164
rect 389548 222216 389600 222222
rect 389548 222158 389600 222164
rect 389560 215422 389588 222158
rect 389548 215416 389600 215422
rect 389548 215358 389600 215364
rect 389456 215280 389508 215286
rect 389456 215222 389508 215228
rect 389468 212537 389496 215222
rect 389270 212528 389326 212537
rect 389270 212463 389326 212472
rect 389454 212528 389510 212537
rect 389454 212463 389510 212472
rect 389284 202910 389312 212463
rect 389272 202904 389324 202910
rect 389272 202846 389324 202852
rect 389548 202904 389600 202910
rect 389548 202846 389600 202852
rect 389560 196110 389588 202846
rect 389548 196104 389600 196110
rect 389548 196046 389600 196052
rect 389456 195968 389508 195974
rect 389456 195910 389508 195916
rect 389468 193225 389496 195910
rect 389270 193216 389326 193225
rect 389270 193151 389326 193160
rect 389454 193216 389510 193225
rect 389454 193151 389510 193160
rect 389284 183598 389312 193151
rect 389272 183592 389324 183598
rect 389272 183534 389324 183540
rect 389548 183592 389600 183598
rect 389548 183534 389600 183540
rect 389560 176798 389588 183534
rect 389548 176792 389600 176798
rect 389548 176734 389600 176740
rect 389456 176656 389508 176662
rect 389456 176598 389508 176604
rect 389468 154562 389496 176598
rect 389456 154556 389508 154562
rect 389456 154498 389508 154504
rect 389640 154556 389692 154562
rect 389640 154498 389692 154504
rect 389652 144945 389680 154498
rect 389362 144936 389418 144945
rect 389362 144871 389418 144880
rect 389638 144936 389694 144945
rect 389638 144871 389694 144880
rect 389376 138038 389404 144871
rect 389364 138032 389416 138038
rect 389364 137974 389416 137980
rect 389456 137964 389508 137970
rect 389456 137906 389508 137912
rect 389468 133890 389496 137906
rect 389456 133884 389508 133890
rect 389456 133826 389508 133832
rect 389180 122868 389232 122874
rect 389180 122810 389232 122816
rect 389192 122754 389220 122810
rect 389192 122726 389312 122754
rect 389284 118833 389312 122726
rect 389270 118824 389326 118833
rect 389270 118759 389326 118768
rect 389454 108896 389510 108905
rect 389454 108831 389510 108840
rect 389468 99210 389496 108831
rect 389456 99204 389508 99210
rect 389456 99146 389508 99152
rect 389364 87916 389416 87922
rect 389364 87858 389416 87864
rect 389376 80102 389404 87858
rect 389364 80096 389416 80102
rect 389364 80038 389416 80044
rect 389456 79960 389508 79966
rect 389456 79902 389508 79908
rect 389468 77246 389496 79902
rect 389456 77240 389508 77246
rect 389456 77182 389508 77188
rect 389364 67652 389416 67658
rect 389364 67594 389416 67600
rect 389376 60738 389404 67594
rect 389192 60710 389404 60738
rect 389192 57934 389220 60710
rect 389180 57928 389232 57934
rect 389180 57870 389232 57876
rect 389272 48340 389324 48346
rect 389272 48282 389324 48288
rect 389284 41426 389312 48282
rect 389284 41398 389404 41426
rect 389376 31822 389404 41398
rect 389364 31816 389416 31822
rect 389364 31758 389416 31764
rect 389456 31680 389508 31686
rect 389456 31622 389508 31628
rect 389468 22273 389496 31622
rect 389454 22264 389510 22273
rect 389454 22199 389510 22208
rect 389362 18048 389418 18057
rect 389362 17983 389418 17992
rect 389376 17950 389404 17983
rect 389364 17944 389416 17950
rect 389364 17886 389416 17892
rect 389456 8356 389508 8362
rect 389456 8298 389508 8304
rect 389088 3528 389140 3534
rect 389088 3470 389140 3476
rect 388444 2848 388496 2854
rect 388444 2790 388496 2796
rect 389468 480 389496 8298
rect 390572 1442 390600 340054
rect 390848 4146 390876 340054
rect 391860 336818 391888 340054
rect 392136 336938 392164 340068
rect 392124 336932 392176 336938
rect 392124 336874 392176 336880
rect 391860 336790 392164 336818
rect 390836 4140 390888 4146
rect 390836 4082 390888 4088
rect 391848 4140 391900 4146
rect 391848 4082 391900 4088
rect 390572 1414 390692 1442
rect 390664 480 390692 1414
rect 391860 480 391888 4082
rect 392136 1442 392164 336790
rect 393056 331242 393084 340190
rect 393162 340054 393268 340082
rect 393622 340054 393912 340082
rect 393056 331214 393176 331242
rect 393148 4146 393176 331214
rect 393136 4140 393188 4146
rect 393136 4082 393188 4088
rect 393240 4078 393268 340054
rect 393884 336938 393912 340054
rect 393596 336932 393648 336938
rect 393596 336874 393648 336880
rect 393872 336932 393924 336938
rect 393872 336874 393924 336880
rect 393228 4072 393280 4078
rect 393228 4014 393280 4020
rect 393608 1442 393636 336874
rect 394068 336802 394096 340068
rect 394528 340054 394634 340082
rect 394056 336796 394108 336802
rect 394056 336738 394108 336744
rect 394528 3330 394556 340054
rect 395080 336802 395108 340068
rect 395554 340054 396028 340082
rect 394608 336796 394660 336802
rect 394608 336738 394660 336744
rect 395068 336796 395120 336802
rect 395068 336738 395120 336744
rect 395896 336796 395948 336802
rect 395896 336738 395948 336744
rect 394620 3534 394648 336738
rect 395908 87242 395936 336738
rect 396000 87242 396028 340054
rect 396092 336870 396120 340068
rect 396080 336864 396132 336870
rect 396080 336806 396132 336812
rect 396552 336802 396580 340068
rect 397012 337482 397040 340068
rect 397000 337476 397052 337482
rect 397000 337418 397052 337424
rect 397472 337074 397500 340068
rect 398024 337686 398052 340068
rect 398484 337890 398512 340068
rect 398472 337884 398524 337890
rect 398472 337826 398524 337832
rect 398944 337754 398972 340068
rect 399864 337770 399892 340190
rect 399970 340054 400168 340082
rect 398932 337748 398984 337754
rect 399864 337742 400076 337770
rect 398932 337690 398984 337696
rect 398012 337680 398064 337686
rect 398012 337622 398064 337628
rect 399484 337680 399536 337686
rect 399484 337622 399536 337628
rect 397460 337068 397512 337074
rect 397460 337010 397512 337016
rect 397460 336932 397512 336938
rect 397460 336874 397512 336880
rect 396540 336796 396592 336802
rect 396540 336738 396592 336744
rect 395896 87236 395948 87242
rect 395896 87178 395948 87184
rect 395988 87236 396040 87242
rect 395988 87178 396040 87184
rect 395986 87136 396042 87145
rect 395816 87106 395986 87122
rect 395804 87100 395986 87106
rect 395856 87094 395986 87100
rect 395986 87071 396042 87080
rect 395804 87042 395856 87048
rect 395896 87032 395948 87038
rect 395896 86974 395948 86980
rect 395988 87032 396040 87038
rect 395988 86974 396040 86980
rect 395436 4140 395488 4146
rect 395436 4082 395488 4088
rect 394608 3528 394660 3534
rect 394608 3470 394660 3476
rect 394516 3324 394568 3330
rect 394516 3266 394568 3272
rect 392136 1414 393084 1442
rect 393608 1414 394280 1442
rect 393056 480 393084 1414
rect 394252 480 394280 1414
rect 395448 480 395476 4082
rect 395908 3058 395936 86974
rect 395896 3052 395948 3058
rect 395896 2994 395948 3000
rect 396000 2990 396028 86974
rect 396632 4072 396684 4078
rect 396632 4014 396684 4020
rect 395988 2984 396040 2990
rect 395988 2926 396040 2932
rect 396644 480 396672 4014
rect 397472 1442 397500 336874
rect 398196 336864 398248 336870
rect 398196 336806 398248 336812
rect 398104 336796 398156 336802
rect 398104 336738 398156 336744
rect 398116 4146 398144 336738
rect 398104 4140 398156 4146
rect 398104 4082 398156 4088
rect 398208 2922 398236 336806
rect 398654 76120 398710 76129
rect 398838 76120 398894 76129
rect 398710 76078 398838 76106
rect 398654 76055 398710 76064
rect 398838 76055 398894 76064
rect 399496 3806 399524 337622
rect 399484 3800 399536 3806
rect 399484 3742 399536 3748
rect 400048 3738 400076 337742
rect 400036 3732 400088 3738
rect 400036 3674 400088 3680
rect 400140 3670 400168 340054
rect 400416 337958 400444 340068
rect 400404 337952 400456 337958
rect 400404 337894 400456 337900
rect 400968 337414 400996 340068
rect 400956 337408 401008 337414
rect 400956 337350 401008 337356
rect 401428 337006 401456 340068
rect 401888 337210 401916 340068
rect 402454 340054 402836 340082
rect 402244 337408 402296 337414
rect 402244 337350 402296 337356
rect 401876 337204 401928 337210
rect 401876 337146 401928 337152
rect 401416 337000 401468 337006
rect 401416 336942 401468 336948
rect 400128 3664 400180 3670
rect 400128 3606 400180 3612
rect 402256 3534 402284 337350
rect 402808 4010 402836 340054
rect 402796 4004 402848 4010
rect 402796 3946 402848 3952
rect 402900 3602 402928 340068
rect 403360 337754 403388 340068
rect 403926 340054 404308 340082
rect 403348 337748 403400 337754
rect 403348 337690 403400 337696
rect 403624 337068 403676 337074
rect 403624 337010 403676 337016
rect 402888 3596 402940 3602
rect 402888 3538 402940 3544
rect 399024 3528 399076 3534
rect 399024 3470 399076 3476
rect 402244 3528 402296 3534
rect 402244 3470 402296 3476
rect 398196 2916 398248 2922
rect 398196 2858 398248 2864
rect 397472 1414 397868 1442
rect 397840 480 397868 1414
rect 399036 480 399064 3470
rect 403636 3466 403664 337010
rect 403624 3460 403676 3466
rect 403624 3402 403676 3408
rect 404280 3398 404308 340054
rect 404372 338026 404400 340068
rect 404360 338020 404412 338026
rect 404360 337962 404412 337968
rect 404832 337618 404860 340068
rect 405398 340054 405688 340082
rect 404820 337612 404872 337618
rect 404820 337554 404872 337560
rect 405004 337000 405056 337006
rect 405004 336942 405056 336948
rect 404912 4140 404964 4146
rect 404912 4082 404964 4088
rect 404268 3392 404320 3398
rect 404268 3334 404320 3340
rect 400220 3324 400272 3330
rect 400220 3266 400272 3272
rect 400232 480 400260 3266
rect 401324 3052 401376 3058
rect 401324 2994 401376 3000
rect 401336 480 401364 2994
rect 402520 2984 402572 2990
rect 402520 2926 402572 2932
rect 402532 480 402560 2926
rect 403716 2916 403768 2922
rect 403716 2858 403768 2864
rect 403728 480 403756 2858
rect 404924 480 404952 4082
rect 405016 3330 405044 336942
rect 405004 3324 405056 3330
rect 405004 3266 405056 3272
rect 405660 3126 405688 340054
rect 405844 337550 405872 340068
rect 406304 338094 406332 340068
rect 406870 340054 407068 340082
rect 406292 338088 406344 338094
rect 406292 338030 406344 338036
rect 406384 337680 406436 337686
rect 406384 337622 406436 337628
rect 405832 337544 405884 337550
rect 405832 337486 405884 337492
rect 405924 337476 405976 337482
rect 405924 337418 405976 337424
rect 405648 3120 405700 3126
rect 405648 3062 405700 3068
rect 405936 610 405964 337418
rect 406396 3058 406424 337622
rect 407040 3194 407068 340054
rect 407316 337822 407344 340068
rect 407304 337816 407356 337822
rect 407304 337758 407356 337764
rect 407776 337074 407804 340068
rect 408342 340054 408448 340082
rect 408802 340054 409184 340082
rect 407764 337068 407816 337074
rect 407764 337010 407816 337016
rect 408420 5438 408448 340054
rect 408776 337884 408828 337890
rect 408776 337826 408828 337832
rect 408408 5432 408460 5438
rect 408408 5374 408460 5380
rect 408500 3800 408552 3806
rect 408500 3742 408552 3748
rect 407304 3460 407356 3466
rect 407304 3402 407356 3408
rect 407028 3188 407080 3194
rect 407028 3130 407080 3136
rect 406384 3052 406436 3058
rect 406384 2994 406436 3000
rect 405924 604 405976 610
rect 405924 546 405976 552
rect 406108 604 406160 610
rect 406108 546 406160 552
rect 406120 480 406148 546
rect 407316 480 407344 3402
rect 408512 480 408540 3742
rect 408788 2938 408816 337826
rect 409156 337482 409184 340054
rect 409144 337476 409196 337482
rect 409144 337418 409196 337424
rect 409248 337414 409276 340068
rect 409236 337408 409288 337414
rect 409236 337350 409288 337356
rect 409144 337068 409196 337074
rect 409144 337010 409196 337016
rect 409156 3262 409184 337010
rect 409800 3398 409828 340068
rect 410260 337754 410288 340068
rect 410734 340054 411208 340082
rect 410248 337748 410300 337754
rect 410248 337690 410300 337696
rect 411076 337748 411128 337754
rect 411076 337690 411128 337696
rect 411088 4146 411116 337690
rect 411076 4140 411128 4146
rect 411076 4082 411128 4088
rect 411180 4078 411208 340054
rect 411272 337686 411300 340068
rect 411746 340054 412128 340082
rect 412206 340054 412588 340082
rect 412100 337770 412128 340054
rect 412100 337742 412496 337770
rect 411260 337680 411312 337686
rect 411260 337622 411312 337628
rect 412364 337680 412416 337686
rect 412364 337622 412416 337628
rect 412376 5370 412404 337622
rect 412364 5364 412416 5370
rect 412364 5306 412416 5312
rect 411168 4072 411220 4078
rect 411168 4014 411220 4020
rect 412468 3942 412496 337742
rect 412456 3936 412508 3942
rect 412456 3878 412508 3884
rect 412560 3874 412588 340054
rect 412744 337618 412772 340068
rect 413218 340054 413600 340082
rect 413284 337952 413336 337958
rect 413284 337894 413336 337900
rect 412732 337612 412784 337618
rect 412732 337554 412784 337560
rect 412548 3868 412600 3874
rect 412548 3810 412600 3816
rect 412088 3732 412140 3738
rect 412088 3674 412140 3680
rect 409788 3392 409840 3398
rect 409788 3334 409840 3340
rect 409144 3256 409196 3262
rect 409144 3198 409196 3204
rect 410892 3052 410944 3058
rect 410892 2994 410944 3000
rect 408788 2910 409736 2938
rect 409708 480 409736 2910
rect 410904 480 410932 2994
rect 412100 480 412128 3674
rect 413192 3664 413244 3670
rect 413192 3606 413244 3612
rect 413204 3346 413232 3606
rect 413296 3534 413324 337894
rect 413572 337736 413600 340054
rect 413664 337958 413692 340068
rect 413652 337952 413704 337958
rect 413652 337894 413704 337900
rect 414216 337890 414244 340068
rect 414676 338026 414704 340068
rect 414664 338020 414716 338026
rect 414664 337962 414716 337968
rect 414204 337884 414256 337890
rect 414204 337826 414256 337832
rect 413572 337708 413968 337736
rect 413836 337612 413888 337618
rect 413836 337554 413888 337560
rect 413848 5302 413876 337554
rect 413836 5296 413888 5302
rect 413836 5238 413888 5244
rect 413940 3670 413968 337708
rect 415136 337142 415164 340068
rect 415308 337884 415360 337890
rect 415308 337826 415360 337832
rect 415124 337136 415176 337142
rect 415124 337078 415176 337084
rect 415320 5234 415348 337826
rect 415596 337754 415624 340068
rect 416148 337822 416176 340068
rect 416136 337816 416188 337822
rect 416136 337758 416188 337764
rect 415584 337748 415636 337754
rect 415584 337690 415636 337696
rect 416504 337748 416556 337754
rect 416504 337690 416556 337696
rect 415308 5228 415360 5234
rect 415308 5170 415360 5176
rect 416516 5166 416544 337690
rect 416504 5160 416556 5166
rect 416504 5102 416556 5108
rect 413928 3664 413980 3670
rect 413928 3606 413980 3612
rect 415676 3596 415728 3602
rect 415676 3538 415728 3544
rect 413284 3528 413336 3534
rect 413284 3470 413336 3476
rect 414480 3528 414532 3534
rect 414480 3470 414532 3476
rect 413204 3318 413324 3346
rect 413296 480 413324 3318
rect 414492 480 414520 3470
rect 415688 480 415716 3538
rect 416608 3058 416636 340068
rect 416688 337816 416740 337822
rect 416688 337758 416740 337764
rect 416700 3806 416728 337758
rect 417068 337754 417096 340068
rect 417424 338088 417476 338094
rect 417424 338030 417476 338036
rect 417056 337748 417108 337754
rect 417056 337690 417108 337696
rect 416964 337204 417016 337210
rect 416964 337146 417016 337152
rect 416688 3800 416740 3806
rect 416688 3742 416740 3748
rect 416872 3324 416924 3330
rect 416872 3266 416924 3272
rect 416596 3052 416648 3058
rect 416596 2994 416648 3000
rect 416884 480 416912 3266
rect 416976 2666 417004 337146
rect 417436 2990 417464 338030
rect 417620 337890 417648 340068
rect 417608 337884 417660 337890
rect 417608 337826 417660 337832
rect 417976 337748 418028 337754
rect 417976 337690 418028 337696
rect 417882 157584 417938 157593
rect 417882 157519 417884 157528
rect 417936 157519 417938 157528
rect 417884 157490 417936 157496
rect 417882 110664 417938 110673
rect 417882 110599 417884 110608
rect 417936 110599 417938 110608
rect 417884 110570 417936 110576
rect 417882 87136 417938 87145
rect 417882 87071 417884 87080
rect 417936 87071 417938 87080
rect 417884 87042 417936 87048
rect 417884 76152 417936 76158
rect 417882 76120 417884 76129
rect 417936 76120 417938 76129
rect 417882 76055 417938 76064
rect 417882 63744 417938 63753
rect 417882 63679 417884 63688
rect 417936 63679 417938 63688
rect 417884 63650 417936 63656
rect 417884 40248 417936 40254
rect 417882 40216 417884 40225
rect 417936 40216 417938 40225
rect 417882 40151 417938 40160
rect 417884 29232 417936 29238
rect 417882 29200 417884 29209
rect 417936 29200 417938 29209
rect 417882 29135 417938 29144
rect 417882 16824 417938 16833
rect 417882 16759 417884 16768
rect 417936 16759 417938 16768
rect 417884 16730 417936 16736
rect 417988 5098 418016 337690
rect 417976 5092 418028 5098
rect 417976 5034 418028 5040
rect 418080 3534 418108 340068
rect 418540 337754 418568 340068
rect 419092 338094 419120 340068
rect 419080 338088 419132 338094
rect 419080 338030 419132 338036
rect 419552 337754 419580 340068
rect 418528 337748 418580 337754
rect 418528 337690 418580 337696
rect 419448 337748 419500 337754
rect 419448 337690 419500 337696
rect 419540 337748 419592 337754
rect 419540 337690 419592 337696
rect 418158 157584 418214 157593
rect 418158 157519 418160 157528
rect 418212 157519 418214 157528
rect 418160 157490 418212 157496
rect 418158 110664 418214 110673
rect 418158 110599 418160 110608
rect 418212 110599 418214 110608
rect 418160 110570 418212 110576
rect 418158 87136 418214 87145
rect 418158 87071 418160 87080
rect 418212 87071 418214 87080
rect 418160 87042 418212 87048
rect 418158 63744 418214 63753
rect 418158 63679 418160 63688
rect 418212 63679 418214 63688
rect 418160 63650 418212 63656
rect 418804 29232 418856 29238
rect 418802 29200 418804 29209
rect 418856 29200 418858 29209
rect 418802 29135 418858 29144
rect 418158 16824 418214 16833
rect 418158 16759 418160 16768
rect 418212 16759 418214 16768
rect 418160 16730 418212 16736
rect 419460 5030 419488 337690
rect 420012 337346 420040 340068
rect 420564 337958 420592 340068
rect 420184 337952 420236 337958
rect 420184 337894 420236 337900
rect 420552 337952 420604 337958
rect 420552 337894 420604 337900
rect 420000 337340 420052 337346
rect 420000 337282 420052 337288
rect 419448 5024 419500 5030
rect 419448 4966 419500 4972
rect 419172 4004 419224 4010
rect 419172 3946 419224 3952
rect 418068 3528 418120 3534
rect 418068 3470 418120 3476
rect 417424 2984 417476 2990
rect 417424 2926 417476 2932
rect 416976 2638 418016 2666
rect 417988 480 418016 2638
rect 419184 480 419212 3946
rect 420196 3330 420224 337894
rect 420276 337816 420328 337822
rect 420276 337758 420328 337764
rect 420288 3670 420316 337758
rect 420828 337748 420880 337754
rect 420828 337690 420880 337696
rect 420736 337340 420788 337346
rect 420736 337282 420788 337288
rect 420368 76152 420420 76158
rect 420366 76120 420368 76129
rect 420420 76120 420422 76129
rect 420366 76055 420422 76064
rect 420368 40248 420420 40254
rect 420366 40216 420368 40225
rect 420420 40216 420422 40225
rect 420366 40151 420422 40160
rect 420748 4962 420776 337282
rect 420736 4956 420788 4962
rect 420736 4898 420788 4904
rect 420368 3732 420420 3738
rect 420368 3674 420420 3680
rect 420276 3664 420328 3670
rect 420276 3606 420328 3612
rect 420184 3324 420236 3330
rect 420184 3266 420236 3272
rect 420380 480 420408 3674
rect 420840 3602 420868 337690
rect 421024 337346 421052 340068
rect 421484 337754 421512 340068
rect 422036 337822 422064 340068
rect 422024 337816 422076 337822
rect 422024 337758 422076 337764
rect 422496 337754 422524 340068
rect 421472 337748 421524 337754
rect 421472 337690 421524 337696
rect 422208 337748 422260 337754
rect 422208 337690 422260 337696
rect 422484 337748 422536 337754
rect 422484 337690 422536 337696
rect 421196 337612 421248 337618
rect 421196 337554 421248 337560
rect 421012 337340 421064 337346
rect 421012 337282 421064 337288
rect 420828 3596 420880 3602
rect 420828 3538 420880 3544
rect 421208 3346 421236 337554
rect 421564 337136 421616 337142
rect 421564 337078 421616 337084
rect 421576 4010 421604 337078
rect 422220 4894 422248 337690
rect 423416 337090 423444 340190
rect 423508 337278 423536 340068
rect 423496 337272 423548 337278
rect 423496 337214 423548 337220
rect 423416 337062 423628 337090
rect 422208 4888 422260 4894
rect 422208 4830 422260 4836
rect 423600 4826 423628 337062
rect 423968 336938 423996 340068
rect 424442 340054 424640 340082
rect 424416 337748 424468 337754
rect 424416 337690 424468 337696
rect 424324 337204 424376 337210
rect 424324 337146 424376 337152
rect 423956 336932 424008 336938
rect 423956 336874 424008 336880
rect 423588 4820 423640 4826
rect 423588 4762 423640 4768
rect 421564 4004 421616 4010
rect 421564 3946 421616 3952
rect 423956 3664 424008 3670
rect 423956 3606 424008 3612
rect 422760 3460 422812 3466
rect 422760 3402 422812 3408
rect 421208 3318 421604 3346
rect 421576 480 421604 3318
rect 422772 480 422800 3402
rect 423968 480 423996 3606
rect 424336 3466 424364 337146
rect 424428 3670 424456 337690
rect 424612 336802 424640 340054
rect 424980 336870 425008 340068
rect 425440 337754 425468 340068
rect 425914 340054 426388 340082
rect 426466 340054 426848 340082
rect 425428 337748 425480 337754
rect 425428 337690 425480 337696
rect 424968 336864 425020 336870
rect 424968 336806 425020 336812
rect 424600 336796 424652 336802
rect 424600 336738 424652 336744
rect 424968 336728 425020 336734
rect 424968 336670 425020 336676
rect 424980 4214 425008 336670
rect 426360 5778 426388 340054
rect 426820 337618 426848 340054
rect 426808 337612 426860 337618
rect 426808 337554 426860 337560
rect 426440 337544 426492 337550
rect 426440 337486 426492 337492
rect 426348 5772 426400 5778
rect 426348 5714 426400 5720
rect 424968 4208 425020 4214
rect 424968 4150 425020 4156
rect 424416 3664 424468 3670
rect 424416 3606 424468 3612
rect 424324 3460 424376 3466
rect 424324 3402 424376 3408
rect 425152 3460 425204 3466
rect 425152 3402 425204 3408
rect 425164 480 425192 3402
rect 426452 3346 426480 337486
rect 426912 337074 426940 340068
rect 427386 340054 427768 340082
rect 427084 337680 427136 337686
rect 427084 337622 427136 337628
rect 426900 337068 426952 337074
rect 426900 337010 426952 337016
rect 427096 3670 427124 337622
rect 427740 5846 427768 340054
rect 427924 337210 427952 340068
rect 428384 337618 428412 340068
rect 428858 340054 429148 340082
rect 428464 337748 428516 337754
rect 428464 337690 428516 337696
rect 428372 337612 428424 337618
rect 428372 337554 428424 337560
rect 427912 337204 427964 337210
rect 427912 337146 427964 337152
rect 427728 5840 427780 5846
rect 427728 5782 427780 5788
rect 427084 3664 427136 3670
rect 427084 3606 427136 3612
rect 426452 3318 427584 3346
rect 426348 3120 426400 3126
rect 426348 3062 426400 3068
rect 426360 480 426388 3062
rect 427556 480 427584 3318
rect 428476 3126 428504 337690
rect 429120 5914 429148 340054
rect 429396 337754 429424 340068
rect 429752 338020 429804 338026
rect 429752 337962 429804 337968
rect 429384 337748 429436 337754
rect 429384 337690 429436 337696
rect 429764 336988 429792 337962
rect 429856 337142 429884 340068
rect 430330 340054 430436 340082
rect 429844 337136 429896 337142
rect 429844 337078 429896 337084
rect 429764 336960 429884 336988
rect 429108 5908 429160 5914
rect 429108 5850 429160 5856
rect 428464 3120 428516 3126
rect 428464 3062 428516 3068
rect 429856 2990 429884 336960
rect 430408 6118 430436 340054
rect 430488 337748 430540 337754
rect 430488 337690 430540 337696
rect 430396 6112 430448 6118
rect 430396 6054 430448 6060
rect 430500 5982 430528 337690
rect 430868 337686 430896 340068
rect 430856 337680 430908 337686
rect 430856 337622 430908 337628
rect 431328 337618 431356 340068
rect 431408 338088 431460 338094
rect 431408 338030 431460 338036
rect 431224 337612 431276 337618
rect 431224 337554 431276 337560
rect 431316 337612 431368 337618
rect 431316 337554 431368 337560
rect 430488 5976 430540 5982
rect 430488 5918 430540 5924
rect 431132 3664 431184 3670
rect 431132 3606 431184 3612
rect 429936 3188 429988 3194
rect 429936 3130 429988 3136
rect 428740 2984 428792 2990
rect 428740 2926 428792 2932
rect 429844 2984 429896 2990
rect 429844 2926 429896 2932
rect 428752 480 428780 2926
rect 429948 480 429976 3130
rect 431144 480 431172 3606
rect 431236 3194 431264 337554
rect 431420 337498 431448 338030
rect 431328 337470 431448 337498
rect 431224 3188 431276 3194
rect 431224 3130 431276 3136
rect 431328 3058 431356 337470
rect 431788 6866 431816 340068
rect 432340 337754 432368 340068
rect 432328 337748 432380 337754
rect 432328 337690 432380 337696
rect 431868 337680 431920 337686
rect 431868 337622 431920 337628
rect 431776 6860 431828 6866
rect 431776 6802 431828 6808
rect 431880 6050 431908 337622
rect 432800 337210 432828 340068
rect 433156 337748 433208 337754
rect 433156 337690 433208 337696
rect 432788 337204 432840 337210
rect 432788 337146 432840 337152
rect 433168 6798 433196 337690
rect 433156 6792 433208 6798
rect 433156 6734 433208 6740
rect 433260 6662 433288 340068
rect 433720 337754 433748 340068
rect 433708 337748 433760 337754
rect 433708 337690 433760 337696
rect 433524 337476 433576 337482
rect 433524 337418 433576 337424
rect 433248 6656 433300 6662
rect 433248 6598 433300 6604
rect 431868 6044 431920 6050
rect 431868 5986 431920 5992
rect 433536 5522 433564 337418
rect 434272 337414 434300 340068
rect 434628 337748 434680 337754
rect 434628 337690 434680 337696
rect 433984 337408 434036 337414
rect 433984 337350 434036 337356
rect 434260 337408 434312 337414
rect 434260 337350 434312 337356
rect 433536 5494 433840 5522
rect 433524 5432 433576 5438
rect 433524 5374 433576 5380
rect 432328 3256 432380 3262
rect 432328 3198 432380 3204
rect 431316 3052 431368 3058
rect 431316 2994 431368 3000
rect 432340 480 432368 3198
rect 433536 480 433564 5374
rect 433812 3074 433840 5494
rect 433996 3398 434024 337350
rect 434640 6730 434668 337690
rect 434732 337686 434760 340068
rect 435192 337754 435220 340068
rect 435744 338094 435772 340068
rect 435732 338088 435784 338094
rect 435732 338030 435784 338036
rect 436204 337754 436232 340068
rect 435180 337748 435232 337754
rect 435180 337690 435232 337696
rect 436008 337748 436060 337754
rect 436008 337690 436060 337696
rect 436192 337748 436244 337754
rect 436192 337690 436244 337696
rect 434720 337680 434772 337686
rect 434720 337622 434772 337628
rect 435916 337680 435968 337686
rect 435916 337622 435968 337628
rect 434628 6724 434680 6730
rect 434628 6666 434680 6672
rect 435928 6594 435956 337622
rect 435916 6588 435968 6594
rect 435916 6530 435968 6536
rect 436020 6526 436048 337690
rect 436664 337686 436692 340068
rect 437216 338026 437244 340068
rect 437204 338020 437256 338026
rect 437204 337962 437256 337968
rect 437388 337748 437440 337754
rect 437388 337690 437440 337696
rect 436652 337680 436704 337686
rect 436652 337622 436704 337628
rect 437296 337680 437348 337686
rect 437296 337622 437348 337628
rect 437202 157584 437258 157593
rect 437202 157519 437204 157528
rect 437256 157519 437258 157528
rect 437204 157490 437256 157496
rect 437202 110664 437258 110673
rect 437202 110599 437204 110608
rect 437256 110599 437258 110608
rect 437204 110570 437256 110576
rect 437204 87168 437256 87174
rect 437202 87136 437204 87145
rect 437256 87136 437258 87145
rect 437202 87071 437258 87080
rect 437202 76120 437258 76129
rect 437202 76055 437204 76064
rect 437256 76055 437258 76064
rect 437204 76026 437256 76032
rect 437202 63744 437258 63753
rect 437202 63679 437204 63688
rect 437256 63679 437258 63688
rect 437204 63650 437256 63656
rect 437204 40248 437256 40254
rect 437202 40216 437204 40225
rect 437256 40216 437258 40225
rect 437202 40151 437258 40160
rect 437202 29200 437258 29209
rect 437202 29135 437204 29144
rect 437256 29135 437258 29144
rect 437204 29106 437256 29112
rect 437202 16824 437258 16833
rect 437202 16759 437204 16768
rect 437256 16759 437258 16768
rect 437204 16730 437256 16736
rect 436008 6520 436060 6526
rect 436008 6462 436060 6468
rect 437308 6322 437336 337622
rect 437400 6458 437428 337690
rect 437676 337482 437704 340068
rect 438150 340054 438624 340082
rect 438124 337816 438176 337822
rect 438124 337758 438176 337764
rect 437664 337476 437716 337482
rect 437664 337418 437716 337424
rect 437478 157584 437534 157593
rect 437478 157519 437480 157528
rect 437532 157519 437534 157528
rect 437480 157490 437532 157496
rect 437478 110664 437534 110673
rect 437478 110599 437480 110608
rect 437532 110599 437534 110608
rect 437480 110570 437532 110576
rect 437480 87168 437532 87174
rect 437478 87136 437480 87145
rect 437532 87136 437534 87145
rect 437478 87071 437534 87080
rect 437478 76120 437534 76129
rect 437478 76055 437480 76064
rect 437532 76055 437534 76064
rect 437480 76026 437532 76032
rect 437478 63744 437534 63753
rect 437478 63679 437480 63688
rect 437532 63679 437534 63688
rect 437480 63650 437532 63656
rect 437480 40248 437532 40254
rect 437478 40216 437480 40225
rect 437532 40216 437534 40225
rect 437478 40151 437534 40160
rect 437478 29200 437534 29209
rect 437478 29135 437480 29144
rect 437532 29135 437534 29144
rect 437480 29106 437532 29112
rect 437478 16824 437534 16833
rect 437478 16759 437480 16768
rect 437532 16759 437534 16768
rect 437480 16730 437532 16736
rect 437388 6452 437440 6458
rect 437388 6394 437440 6400
rect 437296 6316 437348 6322
rect 437296 6258 437348 6264
rect 438136 3398 438164 337758
rect 438596 337668 438624 340054
rect 438688 337822 438716 340068
rect 438676 337816 438728 337822
rect 438676 337758 438728 337764
rect 439148 337754 439176 340068
rect 439622 340054 440096 340082
rect 439136 337748 439188 337754
rect 439136 337690 439188 337696
rect 438596 337640 438808 337668
rect 438676 337476 438728 337482
rect 438676 337418 438728 337424
rect 438688 6390 438716 337418
rect 438676 6384 438728 6390
rect 438676 6326 438728 6332
rect 438780 6254 438808 337640
rect 439504 337408 439556 337414
rect 439504 337350 439556 337356
rect 438768 6248 438820 6254
rect 438768 6190 438820 6196
rect 438216 4140 438268 4146
rect 438216 4082 438268 4088
rect 433984 3392 434036 3398
rect 433984 3334 434036 3340
rect 435824 3392 435876 3398
rect 435824 3334 435876 3340
rect 438124 3392 438176 3398
rect 438124 3334 438176 3340
rect 433812 3046 434668 3074
rect 434640 480 434668 3046
rect 435836 480 435864 3334
rect 437020 3256 437072 3262
rect 437020 3198 437072 3204
rect 437032 480 437060 3198
rect 438228 480 438256 4082
rect 439516 4078 439544 337350
rect 439596 336864 439648 336870
rect 439596 336806 439648 336812
rect 439412 4072 439464 4078
rect 439412 4014 439464 4020
rect 439504 4072 439556 4078
rect 439504 4014 439556 4020
rect 439424 480 439452 4014
rect 439608 2854 439636 336806
rect 440068 7342 440096 340054
rect 440160 337906 440188 340068
rect 440160 337878 440280 337906
rect 440148 337748 440200 337754
rect 440148 337690 440200 337696
rect 440056 7336 440108 7342
rect 440056 7278 440108 7284
rect 440160 6186 440188 337690
rect 440252 337686 440280 337878
rect 440620 337822 440648 340068
rect 441094 340054 441476 340082
rect 440608 337816 440660 337822
rect 440608 337758 440660 337764
rect 440240 337680 440292 337686
rect 440240 337622 440292 337628
rect 441448 7410 441476 340054
rect 441528 337816 441580 337822
rect 441528 337758 441580 337764
rect 441436 7404 441488 7410
rect 441436 7346 441488 7352
rect 440148 6180 440200 6186
rect 440148 6122 440200 6128
rect 440608 5364 440660 5370
rect 440608 5306 440660 5312
rect 439596 2848 439648 2854
rect 439596 2790 439648 2796
rect 440620 480 440648 5306
rect 441540 4282 441568 337758
rect 441632 336870 441660 340068
rect 442092 337822 442120 340068
rect 442566 340054 442856 340082
rect 442356 338020 442408 338026
rect 442356 337962 442408 337968
rect 442080 337816 442132 337822
rect 442080 337758 442132 337764
rect 442264 337544 442316 337550
rect 442264 337486 442316 337492
rect 441620 336864 441672 336870
rect 441620 336806 441672 336812
rect 441528 4276 441580 4282
rect 441528 4218 441580 4224
rect 442276 4146 442304 337486
rect 442264 4140 442316 4146
rect 442264 4082 442316 4088
rect 442368 3942 442396 337962
rect 442828 7478 442856 340054
rect 442908 337816 442960 337822
rect 442908 337758 442960 337764
rect 442816 7472 442868 7478
rect 442816 7414 442868 7420
rect 442920 4350 442948 337758
rect 443104 337482 443132 340068
rect 443564 337686 443592 340068
rect 444038 340054 444236 340082
rect 443552 337680 443604 337686
rect 443552 337622 443604 337628
rect 443092 337476 443144 337482
rect 443092 337418 443144 337424
rect 443644 336864 443696 336870
rect 443644 336806 443696 336812
rect 442908 4344 442960 4350
rect 442908 4286 442960 4292
rect 441804 3936 441856 3942
rect 441804 3878 441856 3884
rect 442356 3936 442408 3942
rect 442356 3878 442408 3884
rect 441816 480 441844 3878
rect 443656 3874 443684 336806
rect 444208 7546 444236 340054
rect 444576 337822 444604 340068
rect 444564 337816 444616 337822
rect 444564 337758 444616 337764
rect 445036 337686 445064 340068
rect 444288 337680 444340 337686
rect 444288 337622 444340 337628
rect 445024 337680 445076 337686
rect 445024 337622 445076 337628
rect 444196 7540 444248 7546
rect 444196 7482 444248 7488
rect 444196 5296 444248 5302
rect 444196 5238 444248 5244
rect 443000 3868 443052 3874
rect 443000 3810 443052 3816
rect 443644 3868 443696 3874
rect 443644 3810 443696 3816
rect 443012 480 443040 3810
rect 444208 480 444236 5238
rect 444300 4418 444328 337622
rect 445496 8294 445524 340068
rect 446048 338026 446076 340068
rect 446036 338020 446088 338026
rect 446036 337962 446088 337968
rect 445668 337816 445720 337822
rect 445668 337758 445720 337764
rect 445576 337680 445628 337686
rect 445576 337622 445628 337628
rect 445484 8288 445536 8294
rect 445484 8230 445536 8236
rect 445588 4486 445616 337622
rect 445576 4480 445628 4486
rect 445576 4422 445628 4428
rect 444288 4412 444340 4418
rect 444288 4354 444340 4360
rect 445680 4146 445708 337758
rect 446508 337686 446536 340068
rect 446496 337680 446548 337686
rect 446496 337622 446548 337628
rect 446968 8226 446996 340068
rect 447048 337680 447100 337686
rect 447048 337622 447100 337628
rect 446956 8220 447008 8226
rect 446956 8162 447008 8168
rect 447060 4554 447088 337622
rect 447520 337550 447548 340068
rect 447994 340054 448376 340082
rect 448244 337680 448296 337686
rect 448244 337622 448296 337628
rect 447508 337544 447560 337550
rect 447508 337486 447560 337492
rect 448256 8158 448284 337622
rect 448244 8152 448296 8158
rect 448244 8094 448296 8100
rect 447784 5228 447836 5234
rect 447784 5170 447836 5176
rect 447048 4548 447100 4554
rect 447048 4490 447100 4496
rect 445668 4140 445720 4146
rect 445668 4082 445720 4088
rect 446312 3936 446364 3942
rect 446364 3884 446536 3890
rect 446312 3878 446536 3884
rect 446324 3862 446536 3878
rect 445392 3800 445444 3806
rect 445392 3742 445444 3748
rect 445404 480 445432 3742
rect 446508 3670 446536 3862
rect 446588 3868 446640 3874
rect 446588 3810 446640 3816
rect 446496 3664 446548 3670
rect 446496 3606 446548 3612
rect 446600 3482 446628 3810
rect 446232 3454 446628 3482
rect 446232 3262 446260 3454
rect 446588 3324 446640 3330
rect 446588 3266 446640 3272
rect 446220 3256 446272 3262
rect 446220 3198 446272 3204
rect 446600 480 446628 3266
rect 447796 480 447824 5170
rect 448348 4622 448376 340054
rect 448440 337686 448468 340068
rect 448992 337822 449020 340068
rect 449466 340054 449848 340082
rect 448980 337816 449032 337822
rect 448980 337758 449032 337764
rect 448428 337680 448480 337686
rect 448428 337622 448480 337628
rect 449164 337612 449216 337618
rect 449164 337554 449216 337560
rect 448428 337544 448480 337550
rect 448428 337486 448480 337492
rect 448336 4616 448388 4622
rect 448336 4558 448388 4564
rect 448440 4078 448468 337486
rect 448428 4072 448480 4078
rect 448428 4014 448480 4020
rect 449176 3738 449204 337554
rect 449820 4690 449848 340054
rect 449912 337686 449940 340068
rect 449900 337680 449952 337686
rect 449900 337622 449952 337628
rect 450464 337618 450492 340068
rect 450938 340054 451136 340082
rect 451004 337680 451056 337686
rect 451004 337622 451056 337628
rect 450452 337612 450504 337618
rect 450452 337554 450504 337560
rect 451016 8090 451044 337622
rect 451004 8084 451056 8090
rect 451004 8026 451056 8032
rect 451108 4758 451136 340054
rect 451384 337822 451412 340068
rect 451844 338026 451872 340068
rect 452410 340054 452608 340082
rect 451832 338020 451884 338026
rect 451832 337962 451884 337968
rect 451372 337816 451424 337822
rect 451372 337758 451424 337764
rect 452476 337816 452528 337822
rect 452476 337758 452528 337764
rect 451188 337612 451240 337618
rect 451188 337554 451240 337560
rect 451096 4752 451148 4758
rect 451096 4694 451148 4700
rect 449808 4684 449860 4690
rect 449808 4626 449860 4632
rect 451200 4010 451228 337554
rect 452488 8022 452516 337758
rect 452476 8016 452528 8022
rect 452476 7958 452528 7964
rect 452580 5506 452608 340054
rect 452856 337822 452884 340068
rect 452844 337816 452896 337822
rect 452844 337758 452896 337764
rect 453316 337618 453344 340068
rect 453764 337816 453816 337822
rect 453764 337758 453816 337764
rect 453304 337612 453356 337618
rect 453304 337554 453356 337560
rect 453776 7954 453804 337758
rect 453764 7948 453816 7954
rect 453764 7890 453816 7896
rect 452568 5500 452620 5506
rect 452568 5442 452620 5448
rect 453868 5438 453896 340068
rect 454328 337822 454356 340068
rect 454788 337958 454816 340068
rect 454776 337952 454828 337958
rect 454776 337894 454828 337900
rect 454316 337816 454368 337822
rect 454316 337758 454368 337764
rect 455236 337816 455288 337822
rect 455236 337758 455288 337764
rect 453948 337612 454000 337618
rect 453948 337554 454000 337560
rect 453856 5432 453908 5438
rect 453856 5374 453908 5380
rect 451280 5160 451332 5166
rect 451280 5102 451332 5108
rect 450176 4004 450228 4010
rect 450176 3946 450228 3952
rect 451188 4004 451240 4010
rect 451188 3946 451240 3952
rect 449164 3732 449216 3738
rect 449164 3674 449216 3680
rect 448980 2984 449032 2990
rect 448980 2926 449032 2932
rect 448992 480 449020 2926
rect 450188 480 450216 3946
rect 451292 480 451320 5102
rect 453960 3942 453988 337554
rect 455248 7886 455276 337758
rect 455236 7880 455288 7886
rect 455236 7822 455288 7828
rect 455340 5370 455368 340068
rect 455604 337884 455656 337890
rect 455604 337826 455656 337832
rect 455328 5364 455380 5370
rect 455328 5306 455380 5312
rect 454868 5092 454920 5098
rect 454868 5034 454920 5040
rect 453672 3936 453724 3942
rect 453672 3878 453724 3884
rect 453948 3936 454000 3942
rect 453948 3878 454000 3884
rect 452476 3868 452528 3874
rect 452476 3810 452528 3816
rect 452488 480 452516 3810
rect 453684 480 453712 3878
rect 454880 480 454908 5034
rect 455616 626 455644 337826
rect 455800 337822 455828 340068
rect 456274 340054 456748 340082
rect 455788 337816 455840 337822
rect 455788 337758 455840 337764
rect 456616 337816 456668 337822
rect 456616 337758 456668 337764
rect 456522 157584 456578 157593
rect 456522 157519 456524 157528
rect 456576 157519 456578 157528
rect 456524 157490 456576 157496
rect 456524 110696 456576 110702
rect 456522 110664 456524 110673
rect 456576 110664 456578 110673
rect 456522 110599 456578 110608
rect 456524 87168 456576 87174
rect 456522 87136 456524 87145
rect 456576 87136 456578 87145
rect 456522 87071 456578 87080
rect 456522 76120 456578 76129
rect 456522 76055 456524 76064
rect 456576 76055 456578 76064
rect 456524 76026 456576 76032
rect 456522 63744 456578 63753
rect 456522 63679 456524 63688
rect 456576 63679 456578 63688
rect 456524 63650 456576 63656
rect 456522 40216 456578 40225
rect 456522 40151 456524 40160
rect 456576 40151 456578 40160
rect 456524 40122 456576 40128
rect 456524 29232 456576 29238
rect 456522 29200 456524 29209
rect 456576 29200 456578 29209
rect 456522 29135 456578 29144
rect 456524 16856 456576 16862
rect 456522 16824 456524 16833
rect 456576 16824 456578 16833
rect 456522 16759 456578 16768
rect 456628 7818 456656 337758
rect 456616 7812 456668 7818
rect 456616 7754 456668 7760
rect 456720 3806 456748 340054
rect 456812 336870 456840 340068
rect 456800 336864 456852 336870
rect 456800 336806 456852 336812
rect 457272 336802 457300 340068
rect 457732 337890 457760 340068
rect 457720 337884 457772 337890
rect 457720 337826 457772 337832
rect 458088 336864 458140 336870
rect 458088 336806 458140 336812
rect 457260 336796 457312 336802
rect 457260 336738 457312 336744
rect 457996 336796 458048 336802
rect 457996 336738 458048 336744
rect 456890 157584 456946 157593
rect 456890 157519 456892 157528
rect 456944 157519 456946 157528
rect 456892 157490 456944 157496
rect 456984 87168 457036 87174
rect 456982 87136 456984 87145
rect 457036 87136 457038 87145
rect 456982 87071 457038 87080
rect 456798 76120 456854 76129
rect 456798 76055 456800 76064
rect 456852 76055 456854 76064
rect 456800 76026 456852 76032
rect 456890 63744 456946 63753
rect 456890 63679 456892 63688
rect 456944 63679 456946 63688
rect 456892 63650 456944 63656
rect 456890 40216 456946 40225
rect 456890 40151 456892 40160
rect 456944 40151 456946 40160
rect 456892 40122 456944 40128
rect 456984 29232 457036 29238
rect 456982 29200 456984 29209
rect 457036 29200 457038 29209
rect 456982 29135 457038 29144
rect 458008 7750 458036 336738
rect 457996 7744 458048 7750
rect 457996 7686 458048 7692
rect 458100 4962 458128 336806
rect 458284 336802 458312 340068
rect 458758 340054 458956 340082
rect 458272 336796 458324 336802
rect 458272 336738 458324 336744
rect 458928 335646 458956 340054
rect 459204 336870 459232 340068
rect 459192 336864 459244 336870
rect 459192 336806 459244 336812
rect 459756 336802 459784 340068
rect 460216 337822 460244 340068
rect 460676 337958 460704 340068
rect 460664 337952 460716 337958
rect 460664 337894 460716 337900
rect 460204 337816 460256 337822
rect 460204 337758 460256 337764
rect 460756 337816 460808 337822
rect 460756 337758 460808 337764
rect 460296 337272 460348 337278
rect 460296 337214 460348 337220
rect 460204 336864 460256 336870
rect 460204 336806 460256 336812
rect 459468 336796 459520 336802
rect 459468 336738 459520 336744
rect 459744 336796 459796 336802
rect 459744 336738 459796 336744
rect 458916 335640 458968 335646
rect 458916 335582 458968 335588
rect 459376 335640 459428 335646
rect 459376 335582 459428 335588
rect 458824 110696 458876 110702
rect 458822 110664 458824 110673
rect 458876 110664 458878 110673
rect 458822 110599 458878 110608
rect 458824 16856 458876 16862
rect 458822 16824 458824 16833
rect 458876 16824 458878 16833
rect 458822 16759 458878 16768
rect 459388 7682 459416 335582
rect 459376 7676 459428 7682
rect 459376 7618 459428 7624
rect 459480 5302 459508 336738
rect 459468 5296 459520 5302
rect 459468 5238 459520 5244
rect 458456 5024 458508 5030
rect 458456 4966 458508 4972
rect 458088 4956 458140 4962
rect 458088 4898 458140 4904
rect 456708 3800 456760 3806
rect 456708 3742 456760 3748
rect 457260 3528 457312 3534
rect 457260 3470 457312 3476
rect 455616 598 456104 626
rect 456076 480 456104 598
rect 457272 480 457300 3470
rect 458468 480 458496 4966
rect 460216 3738 460244 336806
rect 460308 3806 460336 337214
rect 460768 7614 460796 337758
rect 461228 336802 461256 340068
rect 461688 338026 461716 340068
rect 462162 340054 462268 340082
rect 461676 338020 461728 338026
rect 461676 337962 461728 337968
rect 460848 336796 460900 336802
rect 460848 336738 460900 336744
rect 461216 336796 461268 336802
rect 461216 336738 461268 336744
rect 462136 336796 462188 336802
rect 462136 336738 462188 336744
rect 460756 7608 460808 7614
rect 460756 7550 460808 7556
rect 460860 5234 460888 336738
rect 460848 5228 460900 5234
rect 460848 5170 460900 5176
rect 462148 4826 462176 336738
rect 462136 4820 462188 4826
rect 462136 4762 462188 4768
rect 460296 3800 460348 3806
rect 460296 3742 460348 3748
rect 460204 3732 460256 3738
rect 460204 3674 460256 3680
rect 462240 3602 462268 340054
rect 462700 336802 462728 340068
rect 463174 340054 463464 340082
rect 463436 336920 463464 340054
rect 463620 337278 463648 340068
rect 463884 337340 463936 337346
rect 463884 337282 463936 337288
rect 463608 337272 463660 337278
rect 463608 337214 463660 337220
rect 463436 336892 463648 336920
rect 462688 336796 462740 336802
rect 462688 336738 462740 336744
rect 463516 336796 463568 336802
rect 463516 336738 463568 336744
rect 463528 5166 463556 336738
rect 463516 5160 463568 5166
rect 463516 5102 463568 5108
rect 463240 3800 463292 3806
rect 463240 3742 463292 3748
rect 460848 3596 460900 3602
rect 460848 3538 460900 3544
rect 462228 3596 462280 3602
rect 462228 3538 462280 3544
rect 459652 3052 459704 3058
rect 459652 2994 459704 3000
rect 459664 480 459692 2994
rect 460860 480 460888 3538
rect 462044 2780 462096 2786
rect 462044 2722 462096 2728
rect 462056 480 462084 2722
rect 463252 480 463280 3742
rect 463620 3670 463648 336892
rect 463896 325718 463924 337282
rect 464172 336802 464200 340068
rect 464646 340054 464936 340082
rect 464908 336920 464936 340054
rect 465092 337346 465120 340068
rect 465658 340054 465948 340082
rect 466118 340054 466316 340082
rect 465080 337340 465132 337346
rect 465080 337282 465132 337288
rect 464908 336892 465120 336920
rect 465092 336802 465120 336892
rect 464160 336796 464212 336802
rect 464160 336738 464212 336744
rect 464988 336796 465040 336802
rect 464988 336738 465040 336744
rect 465080 336796 465132 336802
rect 465080 336738 465132 336744
rect 463700 325712 463752 325718
rect 463700 325654 463752 325660
rect 463884 325712 463936 325718
rect 463884 325654 463936 325660
rect 463712 316010 463740 325654
rect 463712 315982 463924 316010
rect 463896 306406 463924 315982
rect 463700 306400 463752 306406
rect 463700 306342 463752 306348
rect 463884 306400 463936 306406
rect 463884 306342 463936 306348
rect 463712 296698 463740 306342
rect 463712 296670 463924 296698
rect 463896 287094 463924 296670
rect 463700 287088 463752 287094
rect 463700 287030 463752 287036
rect 463884 287088 463936 287094
rect 463884 287030 463936 287036
rect 463712 277386 463740 287030
rect 463712 277358 463924 277386
rect 463896 267782 463924 277358
rect 463700 267776 463752 267782
rect 463884 267776 463936 267782
rect 463752 267724 463832 267730
rect 463700 267718 463832 267724
rect 463884 267718 463936 267724
rect 463712 267702 463832 267718
rect 463804 267594 463832 267702
rect 463804 267566 463924 267594
rect 463896 263514 463924 267566
rect 463804 263486 463924 263514
rect 463804 260846 463832 263486
rect 463792 260840 463844 260846
rect 463792 260782 463844 260788
rect 463700 251252 463752 251258
rect 463700 251194 463752 251200
rect 463712 244202 463740 251194
rect 463712 244174 463832 244202
rect 463804 234682 463832 244174
rect 463804 234654 464016 234682
rect 463988 231849 464016 234654
rect 463790 231840 463846 231849
rect 463790 231775 463846 231784
rect 463974 231840 464030 231849
rect 463974 231775 464030 231784
rect 463804 222222 463832 231775
rect 463792 222216 463844 222222
rect 463792 222158 463844 222164
rect 464068 222216 464120 222222
rect 464068 222158 464120 222164
rect 464080 215422 464108 222158
rect 464068 215416 464120 215422
rect 464068 215358 464120 215364
rect 463976 215280 464028 215286
rect 463976 215222 464028 215228
rect 463988 212537 464016 215222
rect 463790 212528 463846 212537
rect 463790 212463 463846 212472
rect 463974 212528 464030 212537
rect 463974 212463 464030 212472
rect 463804 202910 463832 212463
rect 463792 202904 463844 202910
rect 463792 202846 463844 202852
rect 464068 202904 464120 202910
rect 464068 202846 464120 202852
rect 464080 196110 464108 202846
rect 464068 196104 464120 196110
rect 464068 196046 464120 196052
rect 463976 195968 464028 195974
rect 463976 195910 464028 195916
rect 463988 193225 464016 195910
rect 463790 193216 463846 193225
rect 463790 193151 463846 193160
rect 463974 193216 464030 193225
rect 463974 193151 464030 193160
rect 463804 183598 463832 193151
rect 463792 183592 463844 183598
rect 463792 183534 463844 183540
rect 464068 183592 464120 183598
rect 464068 183534 464120 183540
rect 464080 176730 464108 183534
rect 463884 176724 463936 176730
rect 463884 176666 463936 176672
rect 464068 176724 464120 176730
rect 464068 176666 464120 176672
rect 463896 166954 463924 176666
rect 463804 166926 463924 166954
rect 463804 164218 463832 166926
rect 463792 164212 463844 164218
rect 463792 164154 463844 164160
rect 464068 164212 464120 164218
rect 464068 164154 464120 164160
rect 464080 154601 464108 164154
rect 463882 154592 463938 154601
rect 463882 154527 463938 154536
rect 464066 154592 464122 154601
rect 464066 154527 464122 154536
rect 463896 130422 463924 154527
rect 463884 130416 463936 130422
rect 463884 130358 463936 130364
rect 464068 130416 464120 130422
rect 464068 130358 464120 130364
rect 464080 125633 464108 130358
rect 463882 125624 463938 125633
rect 463882 125559 463938 125568
rect 464066 125624 464122 125633
rect 464066 125559 464122 125568
rect 463896 118726 463924 125559
rect 463884 118720 463936 118726
rect 463884 118662 463936 118668
rect 463976 118652 464028 118658
rect 463976 118594 464028 118600
rect 463988 109070 464016 118594
rect 463792 109064 463844 109070
rect 463792 109006 463844 109012
rect 463976 109064 464028 109070
rect 463976 109006 464028 109012
rect 463804 103578 463832 109006
rect 463804 103550 463924 103578
rect 463896 93906 463924 103550
rect 463700 93900 463752 93906
rect 463700 93842 463752 93848
rect 463884 93900 463936 93906
rect 463884 93842 463936 93848
rect 463712 93786 463740 93842
rect 463712 93758 463832 93786
rect 463804 80102 463832 93758
rect 463792 80096 463844 80102
rect 463792 80038 463844 80044
rect 463792 79960 463844 79966
rect 463792 79902 463844 79908
rect 463804 70394 463832 79902
rect 463712 70366 463832 70394
rect 463608 3664 463660 3670
rect 463608 3606 463660 3612
rect 463712 610 463740 70366
rect 465000 5098 465028 336738
rect 465920 331242 465948 340054
rect 465920 331214 466224 331242
rect 464988 5092 465040 5098
rect 464988 5034 465040 5040
rect 465632 5024 465684 5030
rect 465632 4966 465684 4972
rect 463700 604 463752 610
rect 463700 546 463752 552
rect 464436 604 464488 610
rect 464436 546 464488 552
rect 464448 480 464476 546
rect 465644 480 465672 4966
rect 466196 4962 466224 331214
rect 466184 4956 466236 4962
rect 466184 4898 466236 4904
rect 466288 3534 466316 340054
rect 466368 337340 466420 337346
rect 466368 337282 466420 337288
rect 466380 3602 466408 337282
rect 466564 336938 466592 340068
rect 467116 337958 467144 340068
rect 467104 337952 467156 337958
rect 467104 337894 467156 337900
rect 467576 337385 467604 340068
rect 468036 337958 468064 340068
rect 468602 340054 468984 340082
rect 467748 337952 467800 337958
rect 467748 337894 467800 337900
rect 468024 337952 468076 337958
rect 468024 337894 468076 337900
rect 467562 337376 467618 337385
rect 467562 337311 467618 337320
rect 466552 336932 466604 336938
rect 466552 336874 466604 336880
rect 467760 4865 467788 337894
rect 468760 8356 468812 8362
rect 468760 8298 468812 8304
rect 467746 4856 467802 4865
rect 467746 4791 467802 4800
rect 466368 3596 466420 3602
rect 466368 3538 466420 3544
rect 466276 3528 466328 3534
rect 466276 3470 466328 3476
rect 467932 3460 467984 3466
rect 467932 3402 467984 3408
rect 466828 2848 466880 2854
rect 466828 2790 466880 2796
rect 466840 480 466868 2790
rect 467944 480 467972 3402
rect 468772 3369 468800 8298
rect 468956 5574 468984 340054
rect 469048 8362 469076 340068
rect 469128 337952 469180 337958
rect 469128 337894 469180 337900
rect 469036 8356 469088 8362
rect 469036 8298 469088 8304
rect 469140 7970 469168 337894
rect 469508 337278 469536 340068
rect 469496 337272 469548 337278
rect 469496 337214 469548 337220
rect 469220 336864 469272 336870
rect 469220 336806 469272 336812
rect 469048 7942 469168 7970
rect 468944 5568 468996 5574
rect 468944 5510 468996 5516
rect 469048 3466 469076 7942
rect 469128 4888 469180 4894
rect 469128 4830 469180 4836
rect 469036 3460 469088 3466
rect 469036 3402 469088 3408
rect 468758 3360 468814 3369
rect 468758 3295 468814 3304
rect 469140 480 469168 4830
rect 469232 610 469260 336806
rect 469876 252550 469904 580246
rect 469968 299470 469996 581198
rect 470048 577924 470100 577930
rect 470048 577866 470100 577872
rect 470060 322930 470088 577866
rect 470152 346390 470180 581266
rect 470244 393310 470272 581334
rect 470336 416770 470364 581402
rect 470428 440230 470456 581470
rect 470520 463690 470548 581538
rect 471256 499526 471284 583646
rect 580540 583636 580592 583642
rect 580540 583578 580592 583584
rect 580264 583568 580316 583574
rect 580264 583510 580316 583516
rect 552664 581188 552716 581194
rect 552664 581130 552716 581136
rect 552676 546446 552704 581130
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 580242 580212 580751
rect 580172 580236 580224 580242
rect 580172 580178 580224 580184
rect 579804 579216 579856 579222
rect 579804 579158 579856 579164
rect 579712 567180 579764 567186
rect 579712 567122 579764 567128
rect 579724 557666 579752 567122
rect 579712 557660 579764 557666
rect 579712 557602 579764 557608
rect 579712 557524 579764 557530
rect 579712 557466 579764 557472
rect 579724 557297 579752 557466
rect 579710 557288 579766 557297
rect 579710 557223 579766 557232
rect 579620 547868 579672 547874
rect 579620 547810 579672 547816
rect 552664 546440 552716 546446
rect 552664 546382 552716 546388
rect 579632 538286 579660 547810
rect 579712 546440 579764 546446
rect 579712 546382 579764 546388
rect 579724 545601 579752 546382
rect 579710 545592 579766 545601
rect 579710 545527 579766 545536
rect 579620 538280 579672 538286
rect 579620 538222 579672 538228
rect 579712 534064 579764 534070
rect 579712 534006 579764 534012
rect 579724 533905 579752 534006
rect 579710 533896 579766 533905
rect 579710 533831 579766 533840
rect 579712 528556 579764 528562
rect 579712 528498 579764 528504
rect 579724 518974 579752 528498
rect 579712 518968 579764 518974
rect 579712 518910 579764 518916
rect 579712 510604 579764 510610
rect 579712 510546 579764 510552
rect 579724 510377 579752 510546
rect 579710 510368 579766 510377
rect 579710 510303 579766 510312
rect 579712 509244 579764 509250
rect 579712 509186 579764 509192
rect 579724 499662 579752 509186
rect 579712 499656 579764 499662
rect 579712 499598 579764 499604
rect 471244 499520 471296 499526
rect 471244 499462 471296 499468
rect 579712 499520 579764 499526
rect 579712 499462 579764 499468
rect 579724 498681 579752 499462
rect 579710 498672 579766 498681
rect 579710 498607 579766 498616
rect 579712 489864 579764 489870
rect 579712 489806 579764 489812
rect 579724 480282 579752 489806
rect 579712 480276 579764 480282
rect 579712 480218 579764 480224
rect 579620 470552 579672 470558
rect 579620 470494 579672 470500
rect 470508 463684 470560 463690
rect 470508 463626 470560 463632
rect 579632 460970 579660 470494
rect 579712 463684 579764 463690
rect 579712 463626 579764 463632
rect 579724 463457 579752 463626
rect 579710 463448 579766 463457
rect 579710 463383 579766 463392
rect 579620 460964 579672 460970
rect 579620 460906 579672 460912
rect 579816 451761 579844 579158
rect 579896 579148 579948 579154
rect 579896 579090 579948 579096
rect 579802 451752 579858 451761
rect 579802 451687 579858 451696
rect 579804 451240 579856 451246
rect 579804 451182 579856 451188
rect 579816 441658 579844 451182
rect 579804 441652 579856 441658
rect 579804 441594 579856 441600
rect 470416 440224 470468 440230
rect 470416 440166 470468 440172
rect 579804 440224 579856 440230
rect 579804 440166 579856 440172
rect 579816 439929 579844 440166
rect 579802 439920 579858 439929
rect 579802 439855 579858 439864
rect 579804 431928 579856 431934
rect 579804 431870 579856 431876
rect 579816 422346 579844 431870
rect 579804 422340 579856 422346
rect 579804 422282 579856 422288
rect 470324 416764 470376 416770
rect 470324 416706 470376 416712
rect 579804 416764 579856 416770
rect 579804 416706 579856 416712
rect 579816 416537 579844 416706
rect 579802 416528 579858 416537
rect 579802 416463 579858 416472
rect 579804 412616 579856 412622
rect 579804 412558 579856 412564
rect 579816 403034 579844 412558
rect 579908 404841 579936 579090
rect 580080 579080 580132 579086
rect 580080 579022 580132 579028
rect 579988 579012 580040 579018
rect 579988 578954 580040 578960
rect 579894 404832 579950 404841
rect 579894 404767 579950 404776
rect 579804 403028 579856 403034
rect 579804 402970 579856 402976
rect 470232 393304 470284 393310
rect 470232 393246 470284 393252
rect 579896 393304 579948 393310
rect 579896 393246 579948 393252
rect 579804 393236 579856 393242
rect 579804 393178 579856 393184
rect 579816 384334 579844 393178
rect 579908 393009 579936 393246
rect 579894 393000 579950 393009
rect 579894 392935 579950 392944
rect 579804 384328 579856 384334
rect 579804 384270 579856 384276
rect 580000 369617 580028 578954
rect 579986 369608 580042 369617
rect 579986 369543 580042 369552
rect 579988 361276 580040 361282
rect 579988 361218 580040 361224
rect 580000 360194 580028 361218
rect 579804 360188 579856 360194
rect 579804 360130 579856 360136
rect 579988 360188 580040 360194
rect 579988 360130 580040 360136
rect 579816 357626 579844 360130
rect 580092 357921 580120 579022
rect 580172 578944 580224 578950
rect 580172 578886 580224 578892
rect 580078 357912 580134 357921
rect 580078 357847 580134 357856
rect 579816 357598 580120 357626
rect 470140 346384 470192 346390
rect 470140 346326 470192 346332
rect 579804 346384 579856 346390
rect 579804 346326 579856 346332
rect 579816 346089 579844 346326
rect 579802 346080 579858 346089
rect 579802 346015 579858 346024
rect 580092 345098 580120 357598
rect 580080 345092 580132 345098
rect 580080 345034 580132 345040
rect 580080 344956 580132 344962
rect 580080 344898 580132 344904
rect 499580 338088 499632 338094
rect 499580 338030 499632 338036
rect 470600 337340 470652 337346
rect 470600 337282 470652 337288
rect 470692 337340 470744 337346
rect 470692 337282 470744 337288
rect 470506 337240 470562 337249
rect 470506 337175 470562 337184
rect 470520 336938 470548 337175
rect 470508 336932 470560 336938
rect 470508 336874 470560 336880
rect 470612 328438 470640 337282
rect 470704 337249 470732 337282
rect 470690 337240 470746 337249
rect 470690 337175 470746 337184
rect 492680 337204 492732 337210
rect 492680 337146 492732 337152
rect 485780 337136 485832 337142
rect 485780 337078 485832 337084
rect 477592 337068 477644 337074
rect 477592 337010 477644 337016
rect 475384 337000 475436 337006
rect 475384 336942 475436 336948
rect 470600 328432 470652 328438
rect 470600 328374 470652 328380
rect 470048 322924 470100 322930
rect 470048 322866 470100 322872
rect 470600 318844 470652 318850
rect 470600 318786 470652 318792
rect 470612 309126 470640 318786
rect 470600 309120 470652 309126
rect 470600 309062 470652 309068
rect 470600 299532 470652 299538
rect 470600 299474 470652 299480
rect 469956 299464 470008 299470
rect 469956 299406 470008 299412
rect 470612 289814 470640 299474
rect 470600 289808 470652 289814
rect 470600 289750 470652 289756
rect 470600 280220 470652 280226
rect 470600 280162 470652 280168
rect 470612 270502 470640 280162
rect 470600 270496 470652 270502
rect 470600 270438 470652 270444
rect 470600 260908 470652 260914
rect 470600 260850 470652 260856
rect 469864 252544 469916 252550
rect 469864 252486 469916 252492
rect 470612 251190 470640 260850
rect 470600 251184 470652 251190
rect 470600 251126 470652 251132
rect 470600 241528 470652 241534
rect 470600 241470 470652 241476
rect 470612 231849 470640 241470
rect 470414 231840 470470 231849
rect 470414 231775 470470 231784
rect 470598 231840 470654 231849
rect 470598 231775 470654 231784
rect 470428 222222 470456 231775
rect 470416 222216 470468 222222
rect 470416 222158 470468 222164
rect 470600 222216 470652 222222
rect 470600 222158 470652 222164
rect 470612 212537 470640 222158
rect 470414 212528 470470 212537
rect 470414 212463 470470 212472
rect 470598 212528 470654 212537
rect 470598 212463 470654 212472
rect 470428 202910 470456 212463
rect 470416 202904 470468 202910
rect 470416 202846 470468 202852
rect 470600 202904 470652 202910
rect 470600 202846 470652 202852
rect 470612 193225 470640 202846
rect 470414 193216 470470 193225
rect 470414 193151 470470 193160
rect 470598 193216 470654 193225
rect 470598 193151 470654 193160
rect 470428 183598 470456 193151
rect 470416 183592 470468 183598
rect 470416 183534 470468 183540
rect 470600 183592 470652 183598
rect 470600 183534 470652 183540
rect 470612 173913 470640 183534
rect 470414 173904 470470 173913
rect 470414 173839 470470 173848
rect 470598 173904 470654 173913
rect 470598 173839 470654 173848
rect 470428 164257 470456 173839
rect 470414 164248 470470 164257
rect 470414 164183 470470 164192
rect 470598 164248 470654 164257
rect 470598 164183 470654 164192
rect 470612 154562 470640 164183
rect 470416 154556 470468 154562
rect 470416 154498 470468 154504
rect 470600 154556 470652 154562
rect 470600 154498 470652 154504
rect 470428 144945 470456 154498
rect 470414 144936 470470 144945
rect 470414 144871 470470 144880
rect 470598 144936 470654 144945
rect 470598 144871 470654 144880
rect 470612 135250 470640 144871
rect 470416 135244 470468 135250
rect 470416 135186 470468 135192
rect 470600 135244 470652 135250
rect 470600 135186 470652 135192
rect 470428 125633 470456 135186
rect 470414 125624 470470 125633
rect 470414 125559 470470 125568
rect 470598 125624 470654 125633
rect 470598 125559 470654 125568
rect 470612 57934 470640 125559
rect 470600 57928 470652 57934
rect 470600 57870 470652 57876
rect 470600 48340 470652 48346
rect 470600 48282 470652 48288
rect 470612 5642 470640 48282
rect 470600 5636 470652 5642
rect 470600 5578 470652 5584
rect 472716 4208 472768 4214
rect 472716 4150 472768 4156
rect 469220 604 469272 610
rect 469220 546 469272 552
rect 470324 604 470376 610
rect 470324 546 470376 552
rect 471520 604 471572 610
rect 471520 546 471572 552
rect 470336 480 470364 546
rect 471532 480 471560 546
rect 472728 480 472756 4150
rect 475396 3126 475424 336942
rect 476026 87272 476082 87281
rect 476026 87207 476082 87216
rect 476040 87122 476068 87207
rect 476210 87136 476266 87145
rect 476040 87094 476210 87122
rect 476210 87071 476266 87080
rect 476026 29336 476082 29345
rect 476026 29271 476082 29280
rect 476040 29186 476068 29271
rect 476210 29200 476266 29209
rect 476040 29158 476210 29186
rect 476210 29135 476266 29144
rect 476304 5772 476356 5778
rect 476304 5714 476356 5720
rect 475108 3120 475160 3126
rect 475108 3062 475160 3068
rect 475384 3120 475436 3126
rect 475384 3062 475436 3068
rect 473912 2916 473964 2922
rect 473912 2858 473964 2864
rect 473924 480 473952 2858
rect 475120 480 475148 3062
rect 476316 480 476344 5714
rect 477604 3346 477632 337010
rect 482926 111072 482982 111081
rect 482926 111007 482982 111016
rect 482940 110673 482968 111007
rect 482926 110664 482982 110673
rect 482926 110599 482982 110608
rect 482926 76528 482982 76537
rect 482926 76463 482982 76472
rect 482940 76129 482968 76463
rect 482926 76120 482982 76129
rect 482926 76055 482982 76064
rect 482926 17232 482982 17241
rect 482926 17167 482982 17176
rect 482940 16833 482968 17167
rect 482926 16824 482982 16833
rect 482926 16759 482982 16768
rect 484584 5976 484636 5982
rect 484584 5918 484636 5924
rect 483480 5908 483532 5914
rect 483480 5850 483532 5856
rect 479892 5840 479944 5846
rect 479892 5782 479944 5788
rect 477604 3318 478736 3346
rect 477500 3120 477552 3126
rect 477500 3062 477552 3068
rect 477512 480 477540 3062
rect 478708 480 478736 3318
rect 479904 480 479932 5782
rect 482284 3120 482336 3126
rect 482284 3062 482336 3068
rect 481088 2984 481140 2990
rect 481088 2926 481140 2932
rect 481100 480 481128 2926
rect 482296 480 482324 3062
rect 483492 480 483520 5850
rect 484596 480 484624 5918
rect 485792 480 485820 337078
rect 487802 110936 487858 110945
rect 487802 110871 487858 110880
rect 487816 110537 487844 110871
rect 487802 110528 487858 110537
rect 487802 110463 487858 110472
rect 491206 87408 491262 87417
rect 491206 87343 491262 87352
rect 491220 87009 491248 87343
rect 491206 87000 491262 87009
rect 491206 86935 491262 86944
rect 487802 76392 487858 76401
rect 487802 76327 487858 76336
rect 487816 75993 487844 76327
rect 487802 75984 487858 75993
rect 487802 75919 487858 75928
rect 491206 29472 491262 29481
rect 491206 29407 491262 29416
rect 491220 29073 491248 29407
rect 491206 29064 491262 29073
rect 491206 28999 491262 29008
rect 487802 17096 487858 17105
rect 487802 17031 487858 17040
rect 487816 16697 487844 17031
rect 487802 16688 487858 16697
rect 487802 16623 487858 16632
rect 490564 6860 490616 6866
rect 490564 6802 490616 6808
rect 486976 6112 487028 6118
rect 486976 6054 487028 6060
rect 486988 480 487016 6054
rect 488172 6044 488224 6050
rect 488172 5986 488224 5992
rect 488184 480 488212 5986
rect 489368 3052 489420 3058
rect 489368 2994 489420 3000
rect 489380 480 489408 2994
rect 490576 480 490604 6802
rect 491760 6792 491812 6798
rect 491760 6734 491812 6740
rect 491772 480 491800 6734
rect 492692 3482 492720 337146
rect 494612 87168 494664 87174
rect 494612 87110 494664 87116
rect 494624 87009 494652 87110
rect 494610 87000 494666 87009
rect 494610 86935 494666 86944
rect 492772 29096 492824 29102
rect 492770 29064 492772 29073
rect 492824 29064 492826 29073
rect 492770 28999 492826 29008
rect 495348 6724 495400 6730
rect 495348 6666 495400 6672
rect 494152 6656 494204 6662
rect 494152 6598 494204 6604
rect 492692 3454 492996 3482
rect 492968 480 492996 3454
rect 494164 480 494192 6598
rect 495360 480 495388 6666
rect 497740 6588 497792 6594
rect 497740 6530 497792 6536
rect 496544 3256 496596 3262
rect 496544 3198 496596 3204
rect 496556 480 496584 3198
rect 497752 480 497780 6530
rect 498936 6520 498988 6526
rect 498936 6462 498988 6468
rect 498948 480 498976 6462
rect 499592 3482 499620 338030
rect 525064 338020 525116 338026
rect 525064 337962 525116 337968
rect 523684 337884 523736 337890
rect 523684 337826 523736 337832
rect 520924 337816 520976 337822
rect 520924 337758 520976 337764
rect 506480 337748 506532 337754
rect 506480 337690 506532 337696
rect 505744 336796 505796 336802
rect 505744 336738 505796 336744
rect 502246 87272 502302 87281
rect 502246 87207 502302 87216
rect 502260 87174 502288 87207
rect 502248 87168 502300 87174
rect 502248 87110 502300 87116
rect 502246 29336 502302 29345
rect 502246 29271 502302 29280
rect 502260 29102 502288 29271
rect 502248 29096 502300 29102
rect 502248 29038 502300 29044
rect 501236 6452 501288 6458
rect 501236 6394 501288 6400
rect 499592 3454 500172 3482
rect 500144 480 500172 3454
rect 501248 480 501276 6394
rect 504824 6384 504876 6390
rect 504824 6326 504876 6332
rect 502432 6316 502484 6322
rect 502432 6258 502484 6264
rect 502444 480 502472 6258
rect 503628 3324 503680 3330
rect 503628 3266 503680 3272
rect 503640 480 503668 3266
rect 504836 480 504864 6326
rect 505756 3194 505784 336738
rect 506020 6248 506072 6254
rect 506020 6190 506072 6196
rect 505744 3188 505796 3194
rect 505744 3130 505796 3136
rect 506032 480 506060 6190
rect 506492 3482 506520 337690
rect 518164 337680 518216 337686
rect 518164 337622 518216 337628
rect 516784 337544 516836 337550
rect 516784 337486 516836 337492
rect 514024 337476 514076 337482
rect 514024 337418 514076 337424
rect 510620 337408 510672 337414
rect 510620 337350 510672 337356
rect 512642 337376 512698 337385
rect 509884 336864 509936 336870
rect 509884 336806 509936 336812
rect 509608 7336 509660 7342
rect 509608 7278 509660 7284
rect 508412 6180 508464 6186
rect 508412 6122 508464 6128
rect 506492 3454 507256 3482
rect 507228 480 507256 3454
rect 508424 480 508452 6122
rect 509620 480 509648 7278
rect 509896 3058 509924 336806
rect 510632 3482 510660 337350
rect 512642 337311 512698 337320
rect 512000 4276 512052 4282
rect 512000 4218 512052 4224
rect 510632 3454 510844 3482
rect 509884 3052 509936 3058
rect 509884 2994 509936 3000
rect 510816 480 510844 3454
rect 512012 480 512040 4218
rect 512656 3262 512684 337311
rect 513196 7404 513248 7410
rect 513196 7346 513248 7352
rect 512644 3256 512696 3262
rect 512644 3198 512696 3204
rect 513208 480 513236 7346
rect 514036 3398 514064 337418
rect 516796 11778 516824 337486
rect 516704 11750 516824 11778
rect 516704 6934 516732 11750
rect 516784 7472 516836 7478
rect 516784 7414 516836 7420
rect 516692 6928 516744 6934
rect 516692 6870 516744 6876
rect 515588 4344 515640 4350
rect 515588 4286 515640 4292
rect 514024 3392 514076 3398
rect 514024 3334 514076 3340
rect 514392 3324 514444 3330
rect 514392 3266 514444 3272
rect 514404 480 514432 3266
rect 515600 480 515628 4286
rect 516796 480 516824 7414
rect 516876 6928 516928 6934
rect 516876 6870 516928 6876
rect 516888 3330 516916 6870
rect 517888 3392 517940 3398
rect 517888 3334 517940 3340
rect 516876 3324 516928 3330
rect 516876 3266 516928 3272
rect 517900 480 517928 3334
rect 518176 2854 518204 337622
rect 520280 7540 520332 7546
rect 520280 7482 520332 7488
rect 519084 4412 519136 4418
rect 519084 4354 519136 4360
rect 518164 2848 518216 2854
rect 518164 2790 518216 2796
rect 519096 480 519124 4354
rect 520292 480 520320 7482
rect 520936 2990 520964 337758
rect 521016 337612 521068 337618
rect 521016 337554 521068 337560
rect 520924 2984 520976 2990
rect 520924 2926 520976 2932
rect 521028 2922 521056 337554
rect 522672 4480 522724 4486
rect 522672 4422 522724 4428
rect 521476 4140 521528 4146
rect 521476 4082 521528 4088
rect 521016 2916 521068 2922
rect 521016 2858 521068 2864
rect 521488 480 521516 4082
rect 522684 480 522712 4422
rect 523696 3058 523724 337826
rect 523868 8288 523920 8294
rect 523868 8230 523920 8236
rect 523684 3052 523736 3058
rect 523684 2994 523736 3000
rect 523880 480 523908 8230
rect 525076 6882 525104 337962
rect 527824 337952 527876 337958
rect 527824 337894 527876 337900
rect 527456 8220 527508 8226
rect 527456 8162 527508 8168
rect 524984 6854 525104 6882
rect 524984 3126 525012 6854
rect 526260 4548 526312 4554
rect 526260 4490 526312 4496
rect 525064 3392 525116 3398
rect 525064 3334 525116 3340
rect 524972 3120 525024 3126
rect 524972 3062 525024 3068
rect 525076 480 525104 3334
rect 526272 480 526300 4490
rect 527468 480 527496 8162
rect 527836 3398 527864 337894
rect 529204 337340 529256 337346
rect 529204 337282 529256 337288
rect 529216 4146 529244 337282
rect 530584 337272 530636 337278
rect 530584 337214 530636 337220
rect 529848 4616 529900 4622
rect 529848 4558 529900 4564
rect 529204 4140 529256 4146
rect 529204 4082 529256 4088
rect 528652 4072 528704 4078
rect 528652 4014 528704 4020
rect 527824 3392 527876 3398
rect 527824 3334 527876 3340
rect 528664 480 528692 4014
rect 529860 480 529888 4558
rect 530596 4078 530624 337214
rect 580092 335442 580120 344898
rect 580080 335436 580132 335442
rect 580080 335378 580132 335384
rect 580080 335300 580132 335306
rect 580080 335242 580132 335248
rect 580092 325718 580120 335242
rect 580080 325712 580132 325718
rect 579986 325680 580042 325689
rect 580080 325654 580132 325660
rect 579986 325615 580042 325624
rect 580000 316130 580028 325615
rect 580080 322924 580132 322930
rect 580080 322866 580132 322872
rect 580092 322697 580120 322866
rect 580078 322688 580134 322697
rect 580078 322623 580134 322632
rect 579988 316124 580040 316130
rect 579988 316066 580040 316072
rect 580080 315988 580132 315994
rect 580080 315930 580132 315936
rect 580092 306406 580120 315930
rect 580184 310865 580212 578886
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 580080 306400 580132 306406
rect 580078 306368 580080 306377
rect 580132 306368 580134 306377
rect 580078 306303 580134 306312
rect 580092 296818 580120 306303
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 299169 580212 299406
rect 580170 299160 580226 299169
rect 580170 299095 580226 299104
rect 580080 296812 580132 296818
rect 580080 296754 580132 296760
rect 580172 296676 580224 296682
rect 580172 296618 580224 296624
rect 580184 287094 580212 296618
rect 580172 287088 580224 287094
rect 580172 287030 580224 287036
rect 580172 277364 580224 277370
rect 580172 277306 580224 277312
rect 580184 275777 580212 277306
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 579620 252544 579672 252550
rect 579620 252486 579672 252492
rect 579632 252249 579660 252486
rect 579618 252240 579674 252249
rect 579618 252175 579674 252184
rect 580276 134881 580304 583510
rect 580356 578672 580408 578678
rect 580356 578614 580408 578620
rect 580368 170105 580396 578614
rect 580448 578604 580500 578610
rect 580448 578546 580500 578552
rect 580460 181937 580488 578546
rect 580552 205329 580580 583578
rect 580908 581120 580960 581126
rect 580908 581062 580960 581068
rect 580816 578876 580868 578882
rect 580816 578818 580868 578824
rect 580632 578808 580684 578814
rect 580632 578750 580684 578756
rect 580644 217025 580672 578750
rect 580724 578740 580776 578746
rect 580724 578682 580776 578688
rect 580736 228857 580764 578682
rect 580828 263945 580856 578818
rect 580920 567186 580948 581062
rect 580908 567180 580960 567186
rect 580908 567122 580960 567128
rect 580908 557592 580960 557598
rect 580908 557534 580960 557540
rect 580920 547874 580948 557534
rect 580908 547868 580960 547874
rect 580908 547810 580960 547816
rect 580908 538280 580960 538286
rect 580908 538222 580960 538228
rect 580920 528562 580948 538222
rect 580908 528556 580960 528562
rect 580908 528498 580960 528504
rect 580908 518968 580960 518974
rect 580908 518910 580960 518916
rect 580920 509250 580948 518910
rect 580908 509244 580960 509250
rect 580908 509186 580960 509192
rect 580908 499588 580960 499594
rect 580908 499530 580960 499536
rect 580920 489870 580948 499530
rect 580908 489864 580960 489870
rect 580908 489806 580960 489812
rect 580908 480276 580960 480282
rect 580908 480218 580960 480224
rect 580920 470558 580948 480218
rect 580908 470552 580960 470558
rect 580908 470494 580960 470500
rect 580908 460964 580960 460970
rect 580908 460906 580960 460912
rect 580920 451246 580948 460906
rect 580908 451240 580960 451246
rect 580908 451182 580960 451188
rect 580908 441652 580960 441658
rect 580908 441594 580960 441600
rect 580920 431934 580948 441594
rect 580908 431928 580960 431934
rect 580908 431870 580960 431876
rect 580908 422340 580960 422346
rect 580908 422282 580960 422288
rect 580920 412622 580948 422282
rect 580908 412616 580960 412622
rect 580908 412558 580960 412564
rect 580908 403028 580960 403034
rect 580908 402970 580960 402976
rect 580920 393310 580948 402970
rect 580908 393304 580960 393310
rect 580908 393246 580960 393252
rect 580908 384328 580960 384334
rect 580908 384270 580960 384276
rect 580920 361282 580948 384270
rect 580908 361276 580960 361282
rect 580908 361218 580960 361224
rect 580908 345092 580960 345098
rect 580908 345034 580960 345040
rect 580920 344962 580948 345034
rect 580908 344956 580960 344962
rect 580908 344898 580960 344904
rect 581000 335436 581052 335442
rect 581000 335378 581052 335384
rect 581012 335306 581040 335378
rect 581000 335300 581052 335306
rect 581000 335242 581052 335248
rect 580908 325712 580960 325718
rect 580906 325680 580908 325689
rect 580960 325680 580962 325689
rect 580906 325615 580962 325624
rect 581000 316124 581052 316130
rect 581000 316066 581052 316072
rect 581012 315994 581040 316066
rect 581000 315988 581052 315994
rect 581000 315930 581052 315936
rect 580908 306400 580960 306406
rect 580906 306368 580908 306377
rect 580960 306368 580962 306377
rect 580906 306303 580962 306312
rect 581000 296812 581052 296818
rect 581000 296754 581052 296760
rect 581012 296682 581040 296754
rect 581000 296676 581052 296682
rect 581000 296618 581052 296624
rect 580908 287088 580960 287094
rect 580908 287030 580960 287036
rect 580920 277370 580948 287030
rect 580908 277364 580960 277370
rect 580908 277306 580960 277312
rect 580814 263936 580870 263945
rect 580814 263871 580870 263880
rect 580722 228848 580778 228857
rect 580722 228783 580778 228792
rect 580630 217016 580686 217025
rect 580630 216951 580686 216960
rect 580538 205320 580594 205329
rect 580538 205255 580594 205264
rect 580446 181928 580502 181937
rect 580446 181863 580502 181872
rect 580354 170096 580410 170105
rect 580354 170031 580410 170040
rect 580262 134872 580318 134881
rect 580262 134807 580318 134816
rect 531044 8152 531096 8158
rect 531044 8094 531096 8100
rect 530584 4072 530636 4078
rect 530584 4014 530636 4020
rect 531056 480 531084 8094
rect 534540 8084 534592 8090
rect 534540 8026 534592 8032
rect 533436 4684 533488 4690
rect 533436 4626 533488 4632
rect 532240 2848 532292 2854
rect 532240 2790 532292 2796
rect 532252 480 532280 2790
rect 533448 480 533476 4626
rect 534552 480 534580 8026
rect 538128 8016 538180 8022
rect 538128 7958 538180 7964
rect 536932 4752 536984 4758
rect 536932 4694 536984 4700
rect 535736 4004 535788 4010
rect 535736 3946 535788 3952
rect 535748 480 535776 3946
rect 536944 480 536972 4694
rect 538140 480 538168 7958
rect 541716 7948 541768 7954
rect 541716 7890 541768 7896
rect 540520 5500 540572 5506
rect 540520 5442 540572 5448
rect 539324 2916 539376 2922
rect 539324 2858 539376 2864
rect 539336 480 539364 2858
rect 540532 480 540560 5442
rect 541728 480 541756 7890
rect 545304 7880 545356 7886
rect 545304 7822 545356 7828
rect 544108 5432 544160 5438
rect 544108 5374 544160 5380
rect 542912 3936 542964 3942
rect 542912 3878 542964 3884
rect 542924 480 542952 3878
rect 544120 480 544148 5374
rect 545316 480 545344 7822
rect 548892 7812 548944 7818
rect 548892 7754 548944 7760
rect 547696 5364 547748 5370
rect 547696 5306 547748 5312
rect 546500 2984 546552 2990
rect 546500 2926 546552 2932
rect 546512 480 546540 2926
rect 547708 480 547736 5306
rect 548904 480 548932 7754
rect 552388 7744 552440 7750
rect 552388 7686 552440 7692
rect 551192 5296 551244 5302
rect 551192 5238 551244 5244
rect 550088 3868 550140 3874
rect 550088 3810 550140 3816
rect 550100 480 550128 3810
rect 551204 480 551232 5238
rect 552400 480 552428 7686
rect 555976 7676 556028 7682
rect 555976 7618 556028 7624
rect 554780 5228 554832 5234
rect 554780 5170 554832 5176
rect 553584 3052 553636 3058
rect 553584 2994 553636 3000
rect 553596 480 553624 2994
rect 554792 480 554820 5170
rect 555988 480 556016 7618
rect 559564 7608 559616 7614
rect 559564 7550 559616 7556
rect 558368 5160 558420 5166
rect 558368 5102 558420 5108
rect 557172 3800 557224 3806
rect 557172 3742 557224 3748
rect 557184 480 557212 3742
rect 558380 480 558408 5102
rect 559576 480 559604 7550
rect 561956 5092 562008 5098
rect 561956 5034 562008 5040
rect 560760 3120 560812 3126
rect 560760 3062 560812 3068
rect 560772 480 560800 3062
rect 561968 480 561996 5034
rect 565544 5024 565596 5030
rect 565544 4966 565596 4972
rect 564348 3732 564400 3738
rect 564348 3674 564400 3680
rect 563152 3188 563204 3194
rect 563152 3130 563204 3136
rect 563164 480 563192 3130
rect 564360 480 564388 3674
rect 565556 480 565584 4966
rect 569040 4956 569092 4962
rect 569040 4898 569092 4904
rect 566740 3664 566792 3670
rect 566740 3606 566792 3612
rect 566752 480 566780 3606
rect 567844 3392 567896 3398
rect 567844 3334 567896 3340
rect 567856 480 567884 3334
rect 569052 480 569080 4898
rect 572628 4888 572680 4894
rect 572628 4830 572680 4836
rect 576214 4856 576270 4865
rect 571432 3596 571484 3602
rect 571432 3538 571484 3544
rect 570236 3256 570288 3262
rect 570236 3198 570288 3204
rect 570248 480 570276 3198
rect 571444 480 571472 3538
rect 572640 480 572668 4830
rect 576214 4791 576270 4800
rect 579804 4820 579856 4826
rect 575020 4140 575072 4146
rect 575020 4082 575072 4088
rect 573824 3528 573876 3534
rect 573824 3470 573876 3476
rect 573836 480 573864 3470
rect 575032 480 575060 4082
rect 576228 480 576256 4791
rect 579804 4762 579856 4768
rect 578608 3460 578660 3466
rect 578608 3402 578660 3408
rect 577412 3324 577464 3330
rect 577412 3266 577464 3272
rect 577424 480 577452 3266
rect 578620 480 578648 3402
rect 579816 480 579844 4762
rect 582196 4072 582248 4078
rect 582196 4014 582248 4020
rect 580998 3360 581054 3369
rect 580998 3295 581054 3304
rect 581012 480 581040 3295
rect 582208 480 582236 4014
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 8114 700304 8170 700360
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 3054 567296 3110 567352
rect 3054 553016 3110 553072
rect 3054 538636 3056 538656
rect 3056 538636 3108 538656
rect 3108 538636 3110 538656
rect 3054 538600 3110 538636
rect 3054 509904 3110 509960
rect 2778 495524 2780 495544
rect 2780 495524 2832 495544
rect 2832 495524 2834 495544
rect 2778 495488 2834 495524
rect 2962 481108 2964 481128
rect 2964 481108 3016 481128
rect 3016 481108 3018 481128
rect 2962 481072 3018 481108
rect 3146 452376 3202 452432
rect 3146 437960 3202 438016
rect 3146 423680 3202 423736
rect 3238 394984 3294 395040
rect 3238 380568 3294 380624
rect 3330 366152 3386 366208
rect 3330 323040 3386 323096
rect 2778 308796 2780 308816
rect 2780 308796 2832 308816
rect 2832 308796 2834 308816
rect 2778 308760 2834 308796
rect 2962 295160 3018 295216
rect 2962 294344 3018 294400
rect 2778 251232 2834 251288
rect 3054 236952 3110 237008
rect 2778 165008 2834 165064
rect 3330 150728 3386 150784
rect 2778 136348 2780 136368
rect 2780 136348 2832 136368
rect 2832 136348 2834 136368
rect 2778 136312 2834 136348
rect 2778 122032 2834 122088
rect 4894 583208 4950 583264
rect 4066 280064 4122 280120
rect 3974 265648 4030 265704
rect 3882 222536 3938 222592
rect 3790 208120 3846 208176
rect 3698 193840 3754 193896
rect 3606 179424 3662 179480
rect 3514 107616 3570 107672
rect 3422 93200 3478 93256
rect 2778 78920 2834 78976
rect 3330 64504 3386 64560
rect 2778 50124 2780 50144
rect 2780 50124 2832 50144
rect 2832 50124 2834 50144
rect 2778 50088 2834 50124
rect 3146 35844 3148 35864
rect 3148 35844 3200 35864
rect 3200 35844 3202 35864
rect 3146 35808 3202 35844
rect 10322 337320 10378 337376
rect 2778 7112 2834 7168
rect 6458 3304 6514 3360
rect 24122 582528 24178 582584
rect 247682 582664 247738 582720
rect 293958 583072 294014 583128
rect 378138 700304 378194 700360
rect 580170 697992 580226 698048
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 460294 583208 460350 583264
rect 420274 582936 420330 582992
rect 426622 582800 426678 582856
rect 462410 582528 462466 582584
rect 231122 579264 231178 579320
rect 232962 579264 233018 579320
rect 235262 579264 235318 579320
rect 237194 579264 237250 579320
rect 239402 579264 239458 579320
rect 241426 579264 241482 579320
rect 243266 579264 243322 579320
rect 249522 579264 249578 579320
rect 468574 579264 468630 579320
rect 51630 6160 51686 6216
rect 132498 337220 132500 337240
rect 132500 337220 132552 337240
rect 132552 337220 132554 337240
rect 132498 337184 132554 337220
rect 142066 337220 142068 337240
rect 142068 337220 142120 337240
rect 142120 337220 142122 337240
rect 142066 337184 142122 337220
rect 151818 337220 151820 337240
rect 151820 337220 151872 337240
rect 151872 337220 151874 337240
rect 151818 337184 151874 337220
rect 161386 337220 161388 337240
rect 161388 337220 161440 337240
rect 161440 337220 161442 337240
rect 161386 337184 161442 337220
rect 171138 337220 171140 337240
rect 171140 337220 171192 337240
rect 171192 337220 171194 337240
rect 171138 337184 171194 337220
rect 180706 337220 180708 337240
rect 180708 337220 180760 337240
rect 180760 337220 180762 337240
rect 180706 337184 180762 337220
rect 190458 337220 190460 337240
rect 190460 337220 190512 337240
rect 190512 337220 190514 337240
rect 190458 337184 190514 337220
rect 200026 337220 200028 337240
rect 200028 337220 200080 337240
rect 200080 337220 200082 337240
rect 200026 337184 200082 337220
rect 209778 337220 209780 337240
rect 209780 337220 209832 337240
rect 209832 337220 209834 337240
rect 209778 337184 209834 337220
rect 219346 337220 219348 337240
rect 219348 337220 219400 337240
rect 219400 337220 219402 337240
rect 219346 337184 219402 337220
rect 132590 8880 132646 8936
rect 129002 7520 129058 7576
rect 208674 4800 208730 4856
rect 229190 337220 229192 337240
rect 229192 337220 229244 337240
rect 229244 337220 229246 337240
rect 229190 337184 229246 337220
rect 231950 337320 232006 337376
rect 230754 202816 230810 202872
rect 231030 202816 231086 202872
rect 230754 183504 230810 183560
rect 231030 183504 231086 183560
rect 232226 202816 232282 202872
rect 232318 202680 232374 202736
rect 232226 183504 232282 183560
rect 232318 183368 232374 183424
rect 232042 3304 232098 3360
rect 234618 337220 234620 337240
rect 234620 337220 234672 337240
rect 234672 337220 234674 337240
rect 234618 337184 234674 337220
rect 234894 135224 234950 135280
rect 235170 135224 235226 135280
rect 235998 135224 236054 135280
rect 235078 96600 235134 96656
rect 235262 96600 235318 96656
rect 236274 251096 236330 251152
rect 236458 251096 236514 251152
rect 236274 231784 236330 231840
rect 236458 231784 236514 231840
rect 236274 212472 236330 212528
rect 236458 212472 236514 212528
rect 236274 193160 236330 193216
rect 236458 193160 236514 193216
rect 236274 183540 236276 183560
rect 236276 183540 236328 183560
rect 236328 183540 236330 183560
rect 236274 183504 236330 183540
rect 236458 183540 236460 183560
rect 236460 183540 236512 183560
rect 236512 183540 236514 183560
rect 236458 183504 236514 183540
rect 236366 173884 236368 173904
rect 236368 173884 236420 173904
rect 236420 173884 236422 173904
rect 236366 173848 236422 173884
rect 236550 173848 236606 173904
rect 236274 164192 236330 164248
rect 236550 164192 236606 164248
rect 236274 135224 236330 135280
rect 241426 40316 241482 40352
rect 241426 40296 241428 40316
rect 241428 40296 241480 40316
rect 241480 40296 241482 40316
rect 241426 16768 241482 16824
rect 241426 16632 241482 16688
rect 244462 259392 244518 259448
rect 244646 259392 244702 259448
rect 244278 241440 244334 241496
rect 244462 241440 244518 241496
rect 244278 222128 244334 222184
rect 244462 222128 244518 222184
rect 244278 202816 244334 202872
rect 244462 202816 244518 202872
rect 244278 154536 244334 154592
rect 244462 154536 244518 154592
rect 244278 135224 244334 135280
rect 244462 135224 244518 135280
rect 244462 115912 244518 115968
rect 244646 115912 244702 115968
rect 244370 44104 244426 44160
rect 244554 44104 244610 44160
rect 245014 40024 245070 40080
rect 247130 144900 247186 144936
rect 247130 144880 247132 144900
rect 247132 144880 247184 144900
rect 247184 144880 247186 144900
rect 247314 144880 247370 144936
rect 247130 96736 247186 96792
rect 247130 96620 247186 96656
rect 247130 96600 247132 96620
rect 247132 96600 247184 96620
rect 247184 96600 247186 96620
rect 248418 29180 248420 29200
rect 248420 29180 248472 29200
rect 248472 29180 248474 29200
rect 248418 29144 248474 29180
rect 249246 336640 249302 336696
rect 249246 327120 249302 327176
rect 249246 321408 249302 321464
rect 249246 317600 249302 317656
rect 249246 298016 249302 298072
rect 249246 288496 249302 288552
rect 249246 288360 249302 288416
rect 249246 278976 249302 279032
rect 249430 277344 249486 277400
rect 249430 267824 249486 267880
rect 249246 212472 249302 212528
rect 249246 205400 249302 205456
rect 249614 202816 249670 202872
rect 249614 196560 249670 196616
rect 249246 191528 249302 191584
rect 249246 182144 249302 182200
rect 249430 180512 249486 180568
rect 249430 173848 249486 173904
rect 249798 75928 249854 75984
rect 250074 288360 250130 288416
rect 250350 288360 250406 288416
rect 250350 154672 250406 154728
rect 250074 154536 250130 154592
rect 250166 124072 250222 124128
rect 250350 124072 250406 124128
rect 250074 75928 250130 75984
rect 249982 6160 250038 6216
rect 251178 87100 251234 87136
rect 251178 87080 251180 87100
rect 251180 87080 251232 87100
rect 251232 87080 251234 87100
rect 251086 16652 251142 16688
rect 251086 16632 251088 16652
rect 251088 16632 251140 16652
rect 251140 16632 251142 16652
rect 251454 241440 251510 241496
rect 251638 241440 251694 241496
rect 251454 222128 251510 222184
rect 251638 222128 251694 222184
rect 251454 202816 251510 202872
rect 251638 202816 251694 202872
rect 251454 183504 251510 183560
rect 251638 183504 251694 183560
rect 251454 154536 251510 154592
rect 251638 154536 251694 154592
rect 251454 21392 251510 21448
rect 251362 8336 251418 8392
rect 253846 76084 253902 76120
rect 253846 76064 253848 76084
rect 253848 76064 253900 76084
rect 253900 76064 253902 76084
rect 253846 40060 253848 40080
rect 253848 40060 253900 40080
rect 253900 40060 253902 40080
rect 253846 40024 253902 40060
rect 257894 29280 257950 29336
rect 259366 75928 259422 75984
rect 259366 16652 259422 16688
rect 259366 16632 259368 16652
rect 259368 16632 259420 16652
rect 259420 16632 259422 16652
rect 259550 280200 259606 280256
rect 259918 280200 259974 280256
rect 259642 202816 259698 202872
rect 259918 202816 259974 202872
rect 259642 164212 259698 164248
rect 259642 164192 259644 164212
rect 259644 164192 259696 164212
rect 259696 164192 259698 164212
rect 259918 164192 259974 164248
rect 259734 116048 259790 116104
rect 259642 115912 259698 115968
rect 259550 96600 259606 96656
rect 259734 96600 259790 96656
rect 260654 87100 260710 87136
rect 260654 87080 260656 87100
rect 260656 87080 260708 87100
rect 260708 87080 260710 87100
rect 262586 202816 262642 202872
rect 262678 202680 262734 202736
rect 262586 183504 262642 183560
rect 262770 183504 262826 183560
rect 262862 40060 262864 40080
rect 262864 40060 262916 40080
rect 262916 40060 262918 40080
rect 262862 40024 262918 40060
rect 262862 29280 262918 29336
rect 262862 29008 262918 29064
rect 264978 248376 265034 248432
rect 264978 180784 265034 180840
rect 265254 277344 265310 277400
rect 265438 277344 265494 277400
rect 265162 259392 265218 259448
rect 265346 259392 265402 259448
rect 265162 248376 265218 248432
rect 265162 202816 265218 202872
rect 265346 202816 265402 202872
rect 265162 180804 265218 180840
rect 265162 180784 265164 180804
rect 265164 180784 265216 180804
rect 265216 180784 265218 180804
rect 265162 125588 265218 125624
rect 265162 125568 265164 125588
rect 265164 125568 265216 125588
rect 265216 125568 265218 125588
rect 265346 125588 265402 125624
rect 265346 125568 265348 125588
rect 265348 125568 265400 125588
rect 265400 125568 265402 125588
rect 265162 96328 265218 96384
rect 265254 88984 265310 89040
rect 266818 270544 266874 270600
rect 266634 270408 266690 270464
rect 267738 259428 267740 259448
rect 267740 259428 267792 259448
rect 267792 259428 267794 259448
rect 267738 259392 267794 259428
rect 267922 259392 267978 259448
rect 267738 248376 267794 248432
rect 268106 248376 268162 248432
rect 267830 82864 267886 82920
rect 268106 82864 268162 82920
rect 267830 81368 267886 81424
rect 268014 81368 268070 81424
rect 267830 62056 267886 62112
rect 268014 62056 268070 62112
rect 270498 162832 270554 162888
rect 270498 125568 270554 125624
rect 270406 110492 270462 110528
rect 270406 110472 270408 110492
rect 270408 110472 270460 110492
rect 270460 110472 270462 110492
rect 270774 293936 270830 293992
rect 270958 293936 271014 293992
rect 270682 240080 270738 240136
rect 270682 239944 270738 240000
rect 270682 202852 270684 202872
rect 270684 202852 270736 202872
rect 270736 202852 270738 202872
rect 270682 202816 270738 202852
rect 270682 202680 270738 202736
rect 270682 183540 270684 183560
rect 270684 183540 270736 183560
rect 270736 183540 270738 183560
rect 270682 183504 270738 183540
rect 270866 183368 270922 183424
rect 270682 162832 270738 162888
rect 270682 125588 270738 125624
rect 270682 125568 270684 125588
rect 270684 125568 270736 125588
rect 270736 125568 270738 125588
rect 272246 230424 272302 230480
rect 272430 230424 272486 230480
rect 272154 202816 272210 202872
rect 272246 190440 272302 190496
rect 272246 162832 272302 162888
rect 272430 162832 272486 162888
rect 272154 125588 272210 125624
rect 272154 125568 272156 125588
rect 272156 125568 272208 125588
rect 272208 125568 272210 125588
rect 272338 125568 272394 125624
rect 273166 63552 273222 63608
rect 278686 157664 278742 157720
rect 278686 157528 278742 157584
rect 278686 110492 278742 110528
rect 278686 110472 278688 110492
rect 278688 110472 278740 110492
rect 278740 110472 278742 110492
rect 278686 63708 278742 63744
rect 278686 63688 278688 63708
rect 278688 63688 278740 63708
rect 278740 63688 278742 63708
rect 280066 110744 280122 110800
rect 280066 110472 280122 110528
rect 282642 157412 282698 157448
rect 282642 157392 282644 157412
rect 282644 157392 282696 157412
rect 282696 157392 282698 157412
rect 282918 87216 282974 87272
rect 282826 87080 282882 87136
rect 282734 40160 282790 40216
rect 282918 40160 282974 40216
rect 283102 7520 283158 7576
rect 284758 306312 284814 306368
rect 284942 306312 284998 306368
rect 284666 296656 284722 296712
rect 284850 296692 284852 296712
rect 284852 296692 284904 296712
rect 284904 296692 284906 296712
rect 284850 296656 284906 296692
rect 284574 269048 284630 269104
rect 284758 269048 284814 269104
rect 284666 249736 284722 249792
rect 284942 249736 284998 249792
rect 284758 201456 284814 201512
rect 284942 201456 284998 201512
rect 284758 135496 284814 135552
rect 284666 135224 284722 135280
rect 284482 8880 284538 8936
rect 285770 202816 285826 202872
rect 285770 153176 285826 153232
rect 286046 261024 286102 261080
rect 285954 260888 286010 260944
rect 286046 249772 286048 249792
rect 286048 249772 286100 249792
rect 286100 249772 286102 249792
rect 286046 249736 286102 249772
rect 285954 249600 286010 249656
rect 285954 222128 286010 222184
rect 286138 222128 286194 222184
rect 285954 220768 286010 220824
rect 286138 220768 286194 220824
rect 285954 202852 285956 202872
rect 285956 202852 286008 202872
rect 286008 202852 286010 202872
rect 285954 202816 286010 202852
rect 285954 183504 286010 183560
rect 285954 183368 286010 183424
rect 285954 153196 286010 153232
rect 285954 153176 285956 153196
rect 285956 153176 286008 153196
rect 286008 153176 286010 153196
rect 286046 103672 286102 103728
rect 285954 103536 286010 103592
rect 288346 16768 288402 16824
rect 288346 16496 288402 16552
rect 288898 238856 288954 238912
rect 289082 238448 289138 238504
rect 288898 157412 288954 157448
rect 288898 157392 288900 157412
rect 288900 157392 288952 157412
rect 288952 157392 288954 157412
rect 290186 240080 290242 240136
rect 290370 240080 290426 240136
rect 290278 201592 290334 201648
rect 290186 201456 290242 201512
rect 289910 190440 289966 190496
rect 290094 190440 290150 190496
rect 290002 172624 290058 172680
rect 290002 172488 290058 172544
rect 291566 258168 291622 258224
rect 291474 258032 291530 258088
rect 291474 248376 291530 248432
rect 291842 248376 291898 248432
rect 291842 201592 291898 201648
rect 291658 201456 291714 201512
rect 291382 190440 291438 190496
rect 291566 190440 291622 190496
rect 291474 172624 291530 172680
rect 291474 172488 291530 172544
rect 294142 267724 294144 267744
rect 294144 267724 294196 267744
rect 294196 267724 294198 267744
rect 294142 267688 294198 267724
rect 294234 267552 294290 267608
rect 295246 248376 295302 248432
rect 295246 29552 295302 29608
rect 295246 29280 295302 29336
rect 295614 258032 295670 258088
rect 295798 258032 295854 258088
rect 295522 248396 295578 248432
rect 295522 248376 295524 248396
rect 295524 248376 295576 248396
rect 295576 248376 295578 248396
rect 295614 238740 295670 238776
rect 295614 238720 295616 238740
rect 295616 238720 295668 238740
rect 295668 238720 295670 238740
rect 295798 238720 295854 238776
rect 296626 63960 296682 64016
rect 296626 63552 296682 63608
rect 296626 29416 296682 29472
rect 296626 29280 296682 29336
rect 296810 258032 296866 258088
rect 296994 258032 297050 258088
rect 296902 151680 296958 151736
rect 297178 151680 297234 151736
rect 297178 142296 297234 142352
rect 296810 142160 296866 142216
rect 298006 16768 298062 16824
rect 298006 16496 298062 16552
rect 299846 249736 299902 249792
rect 299938 249600 299994 249656
rect 299846 200232 299902 200288
rect 299754 200116 299810 200152
rect 299754 200096 299756 200116
rect 299756 200096 299808 200116
rect 299808 200096 299810 200116
rect 301226 306348 301228 306368
rect 301228 306348 301280 306368
rect 301280 306348 301282 306368
rect 301226 306312 301282 306348
rect 301410 306312 301466 306368
rect 302514 285640 302570 285696
rect 302698 285640 302754 285696
rect 302514 266328 302570 266384
rect 302790 266328 302846 266384
rect 302514 258032 302570 258088
rect 302790 258032 302846 258088
rect 302422 143520 302478 143576
rect 302606 143520 302662 143576
rect 304262 87352 304318 87408
rect 304262 86944 304318 87000
rect 306286 157428 306288 157448
rect 306288 157428 306340 157448
rect 306340 157428 306342 157448
rect 306286 157392 306342 157428
rect 306286 110744 306342 110800
rect 306286 110472 306342 110528
rect 306286 29144 306342 29200
rect 306286 28872 306342 28928
rect 306654 266328 306710 266384
rect 306838 266328 306894 266384
rect 306746 200116 306802 200152
rect 306746 200096 306748 200116
rect 306748 200096 306800 200116
rect 306800 200096 306802 200116
rect 306930 200096 306986 200152
rect 306838 161472 306894 161528
rect 307022 161472 307078 161528
rect 307666 110744 307722 110800
rect 306838 93880 306894 93936
rect 307022 93880 307078 93936
rect 307666 28892 307722 28928
rect 307666 28872 307668 28892
rect 307668 28872 307720 28892
rect 307720 28872 307722 28892
rect 309046 76236 309048 76256
rect 309048 76236 309100 76256
rect 309100 76236 309102 76256
rect 309046 76200 309102 76236
rect 307390 3304 307446 3360
rect 310794 193160 310850 193216
rect 311070 193160 311126 193216
rect 310886 153312 310942 153368
rect 310794 153196 310850 153232
rect 310794 153176 310796 153196
rect 310796 153176 310848 153196
rect 310848 153176 310850 153196
rect 310794 67768 310850 67824
rect 310794 67632 310850 67688
rect 312082 4936 312138 4992
rect 314566 157428 314568 157448
rect 314568 157428 314620 157448
rect 314620 157428 314622 157448
rect 314566 157392 314622 157428
rect 315946 110472 316002 110528
rect 315946 28892 316002 28928
rect 315946 28872 315948 28892
rect 315948 28872 316000 28892
rect 316000 28872 316002 28892
rect 315946 16360 316002 16416
rect 315946 16088 316002 16144
rect 315946 4972 315948 4992
rect 315948 4972 316000 4992
rect 316000 4972 316002 4992
rect 315946 4936 316002 4972
rect 314658 4800 314714 4856
rect 317326 111016 317382 111072
rect 317326 110472 317382 110528
rect 317326 76236 317328 76256
rect 317328 76236 317380 76256
rect 317380 76236 317382 76256
rect 317326 76200 317382 76236
rect 317326 29280 317382 29336
rect 317326 28872 317382 28928
rect 317326 16632 317382 16688
rect 317326 16360 317382 16416
rect 318706 76200 318762 76256
rect 318706 75928 318762 75984
rect 322202 29280 322258 29336
rect 322202 29008 322258 29064
rect 322202 16632 322258 16688
rect 322202 16360 322258 16416
rect 323490 278740 323492 278760
rect 323492 278740 323544 278760
rect 323544 278740 323546 278760
rect 323490 278704 323546 278740
rect 323674 278704 323730 278760
rect 323214 259392 323270 259448
rect 323398 259392 323454 259448
rect 323306 193196 323308 193216
rect 323308 193196 323360 193216
rect 323360 193196 323362 193216
rect 323306 193160 323362 193196
rect 323490 193196 323492 193216
rect 323492 193196 323544 193216
rect 323544 193196 323546 193216
rect 323490 193160 323546 193196
rect 324502 182164 324558 182200
rect 324502 182144 324504 182164
rect 324504 182144 324556 182164
rect 324556 182144 324558 182164
rect 324870 182144 324926 182200
rect 324594 125588 324650 125624
rect 324594 125568 324596 125588
rect 324596 125568 324648 125588
rect 324648 125568 324650 125588
rect 324778 125588 324834 125624
rect 324778 125568 324780 125588
rect 324780 125568 324832 125588
rect 324832 125568 324834 125588
rect 324594 104760 324650 104816
rect 324778 104624 324834 104680
rect 325974 231784 326030 231840
rect 326066 231648 326122 231704
rect 325882 202816 325938 202872
rect 325974 202680 326030 202736
rect 325882 183504 325938 183560
rect 326066 183504 326122 183560
rect 325974 172488 326030 172544
rect 326250 172488 326306 172544
rect 325974 153176 326030 153232
rect 326158 153176 326214 153232
rect 325974 145016 326030 145072
rect 325882 144900 325938 144936
rect 325882 144880 325884 144900
rect 325884 144880 325936 144900
rect 325936 144880 325938 144900
rect 327170 144900 327226 144936
rect 327170 144880 327172 144900
rect 327172 144880 327224 144900
rect 327224 144880 327226 144900
rect 327354 144900 327410 144936
rect 327354 144880 327356 144900
rect 327356 144880 327408 144900
rect 327408 144880 327410 144900
rect 327262 113192 327318 113248
rect 327446 113192 327502 113248
rect 327170 103400 327226 103456
rect 327446 103264 327502 103320
rect 328458 110880 328514 110936
rect 328458 110608 328514 110664
rect 328274 16768 328330 16824
rect 328274 16496 328330 16552
rect 329930 248376 329986 248432
rect 329930 220768 329986 220824
rect 329930 202852 329932 202872
rect 329932 202852 329984 202872
rect 329984 202852 329986 202872
rect 329930 202816 329986 202852
rect 329930 153176 329986 153232
rect 329930 48320 329986 48376
rect 330114 296656 330170 296712
rect 330666 296656 330722 296712
rect 330206 269084 330208 269104
rect 330208 269084 330260 269104
rect 330260 269084 330262 269104
rect 330206 269048 330262 269084
rect 330390 269048 330446 269104
rect 330298 248376 330354 248432
rect 330206 220768 330262 220824
rect 330114 202852 330116 202872
rect 330116 202852 330168 202872
rect 330168 202852 330170 202872
rect 330114 202816 330170 202852
rect 330114 182144 330170 182200
rect 330298 182144 330354 182200
rect 330114 162852 330170 162888
rect 330114 162832 330116 162852
rect 330116 162832 330168 162852
rect 330168 162832 330170 162852
rect 330298 162832 330354 162888
rect 330206 153176 330262 153232
rect 330114 48320 330170 48376
rect 331402 222128 331458 222184
rect 331586 222128 331642 222184
rect 331402 202816 331458 202872
rect 331586 202816 331642 202872
rect 331402 183504 331458 183560
rect 331586 183504 331642 183560
rect 331862 29552 331918 29608
rect 331862 29280 331918 29336
rect 337106 287000 337162 287056
rect 337290 287000 337346 287056
rect 337014 256672 337070 256728
rect 337198 256672 337254 256728
rect 337106 201456 337162 201512
rect 337382 201456 337438 201512
rect 337106 135224 337162 135280
rect 337290 135224 337346 135280
rect 336738 16668 336740 16688
rect 336740 16668 336792 16688
rect 336792 16668 336794 16688
rect 336738 16632 336794 16668
rect 338210 16904 338266 16960
rect 338670 241440 338726 241496
rect 338854 241440 338910 241496
rect 338670 222128 338726 222184
rect 338854 222128 338910 222184
rect 338670 202816 338726 202872
rect 338854 202816 338910 202872
rect 338854 154672 338910 154728
rect 338854 154536 338910 154592
rect 341062 260888 341118 260944
rect 341430 260888 341486 260944
rect 341246 179424 341302 179480
rect 341430 179424 341486 179480
rect 341062 132504 341118 132560
rect 341246 132504 341302 132560
rect 350630 3848 350686 3904
rect 354126 3984 354182 4040
rect 354218 3884 354220 3904
rect 354220 3884 354272 3904
rect 354272 3884 354274 3904
rect 354218 3848 354274 3884
rect 353666 3032 353722 3088
rect 356242 3304 356298 3360
rect 357438 220768 357494 220824
rect 357622 220768 357678 220824
rect 357438 211112 357494 211168
rect 357714 211112 357770 211168
rect 357714 193160 357770 193216
rect 357898 193160 357954 193216
rect 357622 164328 357678 164384
rect 357530 164192 357586 164248
rect 357254 133864 357310 133920
rect 357438 133864 357494 133920
rect 358542 278704 358598 278760
rect 358726 278704 358782 278760
rect 358542 259392 358598 259448
rect 358726 259392 358782 259448
rect 358542 240080 358598 240136
rect 358726 240080 358782 240136
rect 358542 220768 358598 220824
rect 358726 220768 358782 220824
rect 358542 211112 358598 211168
rect 358726 211112 358782 211168
rect 358542 182144 358598 182200
rect 358726 182144 358782 182200
rect 358726 106528 358782 106584
rect 358726 106256 358782 106312
rect 358174 4020 358176 4040
rect 358176 4020 358228 4040
rect 358228 4020 358230 4040
rect 358174 3984 358230 4020
rect 356794 3032 356850 3088
rect 360934 327256 360990 327312
rect 360474 327120 360530 327176
rect 360106 157528 360162 157584
rect 360290 157528 360346 157584
rect 360382 96736 360438 96792
rect 360290 96620 360346 96656
rect 360290 96600 360292 96620
rect 360292 96600 360344 96620
rect 360344 96600 360346 96620
rect 360198 63824 360254 63880
rect 360106 63688 360162 63744
rect 360106 40160 360162 40216
rect 360290 40160 360346 40216
rect 366822 183504 366878 183560
rect 367006 241440 367062 241496
rect 367006 231920 367062 231976
rect 367006 183540 367008 183560
rect 367008 183540 367060 183560
rect 367060 183540 367062 183560
rect 367006 183504 367062 183540
rect 367006 173848 367062 173904
rect 367006 164192 367062 164248
rect 367006 96736 367062 96792
rect 367006 96620 367062 96656
rect 367006 96600 367008 96620
rect 367008 96600 367060 96620
rect 367060 96600 367062 96620
rect 367098 29044 367100 29064
rect 367100 29044 367152 29064
rect 367152 29044 367154 29064
rect 367098 29008 367154 29044
rect 372526 241440 372582 241496
rect 372710 241440 372766 241496
rect 372526 222128 372582 222184
rect 372710 222128 372766 222184
rect 372526 202816 372582 202872
rect 372710 202816 372766 202872
rect 372526 183504 372582 183560
rect 372710 183504 372766 183560
rect 374366 114688 374422 114744
rect 374274 114552 374330 114608
rect 376758 338020 376814 338056
rect 376758 338000 376760 338020
rect 376760 338000 376812 338020
rect 376812 338000 376814 338020
rect 376850 318824 376906 318880
rect 377126 318824 377182 318880
rect 376942 241440 376998 241496
rect 377126 241440 377182 241496
rect 376942 222128 376998 222184
rect 377126 222128 377182 222184
rect 376942 202816 376998 202872
rect 377126 202816 377182 202872
rect 376942 183504 376998 183560
rect 377126 183504 377182 183560
rect 376942 154536 376998 154592
rect 377126 154536 377182 154592
rect 376942 135224 376998 135280
rect 377126 135224 377182 135280
rect 376758 87100 376814 87136
rect 376758 87080 376760 87100
rect 376760 87080 376812 87100
rect 376812 87080 376814 87100
rect 376666 29280 376722 29336
rect 377126 29008 377182 29064
rect 377310 29008 377366 29064
rect 379334 338000 379390 338056
rect 386234 86944 386290 87000
rect 386418 86944 386474 87000
rect 388994 251096 389050 251152
rect 389178 251096 389234 251152
rect 389270 231784 389326 231840
rect 389454 231784 389510 231840
rect 389270 212472 389326 212528
rect 389454 212472 389510 212528
rect 389270 193160 389326 193216
rect 389454 193160 389510 193216
rect 389362 144880 389418 144936
rect 389638 144880 389694 144936
rect 389270 118768 389326 118824
rect 389454 108840 389510 108896
rect 389454 22208 389510 22264
rect 389362 17992 389418 18048
rect 395986 87080 396042 87136
rect 398654 76064 398710 76120
rect 398838 76064 398894 76120
rect 417882 157548 417938 157584
rect 417882 157528 417884 157548
rect 417884 157528 417936 157548
rect 417936 157528 417938 157548
rect 417882 110628 417938 110664
rect 417882 110608 417884 110628
rect 417884 110608 417936 110628
rect 417936 110608 417938 110628
rect 417882 87100 417938 87136
rect 417882 87080 417884 87100
rect 417884 87080 417936 87100
rect 417936 87080 417938 87100
rect 417882 76100 417884 76120
rect 417884 76100 417936 76120
rect 417936 76100 417938 76120
rect 417882 76064 417938 76100
rect 417882 63708 417938 63744
rect 417882 63688 417884 63708
rect 417884 63688 417936 63708
rect 417936 63688 417938 63708
rect 417882 40196 417884 40216
rect 417884 40196 417936 40216
rect 417936 40196 417938 40216
rect 417882 40160 417938 40196
rect 417882 29180 417884 29200
rect 417884 29180 417936 29200
rect 417936 29180 417938 29200
rect 417882 29144 417938 29180
rect 417882 16788 417938 16824
rect 417882 16768 417884 16788
rect 417884 16768 417936 16788
rect 417936 16768 417938 16788
rect 418158 157548 418214 157584
rect 418158 157528 418160 157548
rect 418160 157528 418212 157548
rect 418212 157528 418214 157548
rect 418158 110628 418214 110664
rect 418158 110608 418160 110628
rect 418160 110608 418212 110628
rect 418212 110608 418214 110628
rect 418158 87100 418214 87136
rect 418158 87080 418160 87100
rect 418160 87080 418212 87100
rect 418212 87080 418214 87100
rect 418158 63708 418214 63744
rect 418158 63688 418160 63708
rect 418160 63688 418212 63708
rect 418212 63688 418214 63708
rect 418802 29180 418804 29200
rect 418804 29180 418856 29200
rect 418856 29180 418858 29200
rect 418802 29144 418858 29180
rect 418158 16788 418214 16824
rect 418158 16768 418160 16788
rect 418160 16768 418212 16788
rect 418212 16768 418214 16788
rect 420366 76100 420368 76120
rect 420368 76100 420420 76120
rect 420420 76100 420422 76120
rect 420366 76064 420422 76100
rect 420366 40196 420368 40216
rect 420368 40196 420420 40216
rect 420420 40196 420422 40216
rect 420366 40160 420422 40196
rect 437202 157548 437258 157584
rect 437202 157528 437204 157548
rect 437204 157528 437256 157548
rect 437256 157528 437258 157548
rect 437202 110628 437258 110664
rect 437202 110608 437204 110628
rect 437204 110608 437256 110628
rect 437256 110608 437258 110628
rect 437202 87116 437204 87136
rect 437204 87116 437256 87136
rect 437256 87116 437258 87136
rect 437202 87080 437258 87116
rect 437202 76084 437258 76120
rect 437202 76064 437204 76084
rect 437204 76064 437256 76084
rect 437256 76064 437258 76084
rect 437202 63708 437258 63744
rect 437202 63688 437204 63708
rect 437204 63688 437256 63708
rect 437256 63688 437258 63708
rect 437202 40196 437204 40216
rect 437204 40196 437256 40216
rect 437256 40196 437258 40216
rect 437202 40160 437258 40196
rect 437202 29164 437258 29200
rect 437202 29144 437204 29164
rect 437204 29144 437256 29164
rect 437256 29144 437258 29164
rect 437202 16788 437258 16824
rect 437202 16768 437204 16788
rect 437204 16768 437256 16788
rect 437256 16768 437258 16788
rect 437478 157548 437534 157584
rect 437478 157528 437480 157548
rect 437480 157528 437532 157548
rect 437532 157528 437534 157548
rect 437478 110628 437534 110664
rect 437478 110608 437480 110628
rect 437480 110608 437532 110628
rect 437532 110608 437534 110628
rect 437478 87116 437480 87136
rect 437480 87116 437532 87136
rect 437532 87116 437534 87136
rect 437478 87080 437534 87116
rect 437478 76084 437534 76120
rect 437478 76064 437480 76084
rect 437480 76064 437532 76084
rect 437532 76064 437534 76084
rect 437478 63708 437534 63744
rect 437478 63688 437480 63708
rect 437480 63688 437532 63708
rect 437532 63688 437534 63708
rect 437478 40196 437480 40216
rect 437480 40196 437532 40216
rect 437532 40196 437534 40216
rect 437478 40160 437534 40196
rect 437478 29164 437534 29200
rect 437478 29144 437480 29164
rect 437480 29144 437532 29164
rect 437532 29144 437534 29164
rect 437478 16788 437534 16824
rect 437478 16768 437480 16788
rect 437480 16768 437532 16788
rect 437532 16768 437534 16788
rect 456522 157548 456578 157584
rect 456522 157528 456524 157548
rect 456524 157528 456576 157548
rect 456576 157528 456578 157548
rect 456522 110644 456524 110664
rect 456524 110644 456576 110664
rect 456576 110644 456578 110664
rect 456522 110608 456578 110644
rect 456522 87116 456524 87136
rect 456524 87116 456576 87136
rect 456576 87116 456578 87136
rect 456522 87080 456578 87116
rect 456522 76084 456578 76120
rect 456522 76064 456524 76084
rect 456524 76064 456576 76084
rect 456576 76064 456578 76084
rect 456522 63708 456578 63744
rect 456522 63688 456524 63708
rect 456524 63688 456576 63708
rect 456576 63688 456578 63708
rect 456522 40180 456578 40216
rect 456522 40160 456524 40180
rect 456524 40160 456576 40180
rect 456576 40160 456578 40180
rect 456522 29180 456524 29200
rect 456524 29180 456576 29200
rect 456576 29180 456578 29200
rect 456522 29144 456578 29180
rect 456522 16804 456524 16824
rect 456524 16804 456576 16824
rect 456576 16804 456578 16824
rect 456522 16768 456578 16804
rect 456890 157548 456946 157584
rect 456890 157528 456892 157548
rect 456892 157528 456944 157548
rect 456944 157528 456946 157548
rect 456982 87116 456984 87136
rect 456984 87116 457036 87136
rect 457036 87116 457038 87136
rect 456982 87080 457038 87116
rect 456798 76084 456854 76120
rect 456798 76064 456800 76084
rect 456800 76064 456852 76084
rect 456852 76064 456854 76084
rect 456890 63708 456946 63744
rect 456890 63688 456892 63708
rect 456892 63688 456944 63708
rect 456944 63688 456946 63708
rect 456890 40180 456946 40216
rect 456890 40160 456892 40180
rect 456892 40160 456944 40180
rect 456944 40160 456946 40180
rect 456982 29180 456984 29200
rect 456984 29180 457036 29200
rect 457036 29180 457038 29200
rect 456982 29144 457038 29180
rect 458822 110644 458824 110664
rect 458824 110644 458876 110664
rect 458876 110644 458878 110664
rect 458822 110608 458878 110644
rect 458822 16804 458824 16824
rect 458824 16804 458876 16824
rect 458876 16804 458878 16824
rect 458822 16768 458878 16804
rect 463790 231784 463846 231840
rect 463974 231784 464030 231840
rect 463790 212472 463846 212528
rect 463974 212472 464030 212528
rect 463790 193160 463846 193216
rect 463974 193160 464030 193216
rect 463882 154536 463938 154592
rect 464066 154536 464122 154592
rect 463882 125568 463938 125624
rect 464066 125568 464122 125624
rect 467562 337320 467618 337376
rect 467746 4800 467802 4856
rect 468758 3304 468814 3360
rect 580170 580760 580226 580816
rect 579710 557232 579766 557288
rect 579710 545536 579766 545592
rect 579710 533840 579766 533896
rect 579710 510312 579766 510368
rect 579710 498616 579766 498672
rect 579710 463392 579766 463448
rect 579802 451696 579858 451752
rect 579802 439864 579858 439920
rect 579802 416472 579858 416528
rect 579894 404776 579950 404832
rect 579894 392944 579950 393000
rect 579986 369552 580042 369608
rect 580078 357856 580134 357912
rect 579802 346024 579858 346080
rect 470506 337184 470562 337240
rect 470690 337184 470746 337240
rect 470414 231784 470470 231840
rect 470598 231784 470654 231840
rect 470414 212472 470470 212528
rect 470598 212472 470654 212528
rect 470414 193160 470470 193216
rect 470598 193160 470654 193216
rect 470414 173848 470470 173904
rect 470598 173848 470654 173904
rect 470414 164192 470470 164248
rect 470598 164192 470654 164248
rect 470414 144880 470470 144936
rect 470598 144880 470654 144936
rect 470414 125568 470470 125624
rect 470598 125568 470654 125624
rect 476026 87216 476082 87272
rect 476210 87080 476266 87136
rect 476026 29280 476082 29336
rect 476210 29144 476266 29200
rect 482926 111016 482982 111072
rect 482926 110608 482982 110664
rect 482926 76472 482982 76528
rect 482926 76064 482982 76120
rect 482926 17176 482982 17232
rect 482926 16768 482982 16824
rect 487802 110880 487858 110936
rect 487802 110472 487858 110528
rect 491206 87352 491262 87408
rect 491206 86944 491262 87000
rect 487802 76336 487858 76392
rect 487802 75928 487858 75984
rect 491206 29416 491262 29472
rect 491206 29008 491262 29064
rect 487802 17040 487858 17096
rect 487802 16632 487858 16688
rect 494610 86944 494666 87000
rect 492770 29044 492772 29064
rect 492772 29044 492824 29064
rect 492824 29044 492826 29064
rect 492770 29008 492826 29044
rect 502246 87216 502302 87272
rect 502246 29280 502302 29336
rect 512642 337320 512698 337376
rect 579986 325624 580042 325680
rect 580078 322632 580134 322688
rect 580170 310800 580226 310856
rect 580078 306348 580080 306368
rect 580080 306348 580132 306368
rect 580132 306348 580134 306368
rect 580078 306312 580134 306348
rect 580170 299104 580226 299160
rect 580170 275712 580226 275768
rect 579618 252184 579674 252240
rect 580906 325660 580908 325680
rect 580908 325660 580960 325680
rect 580960 325660 580962 325680
rect 580906 325624 580962 325660
rect 580906 306348 580908 306368
rect 580908 306348 580960 306368
rect 580960 306348 580962 306368
rect 580906 306312 580962 306348
rect 580814 263880 580870 263936
rect 580722 228792 580778 228848
rect 580630 216960 580686 217016
rect 580538 205264 580594 205320
rect 580446 181872 580502 181928
rect 580354 170040 580410 170096
rect 580262 134816 580318 134872
rect 576214 4800 576270 4856
rect 580998 3304 581054 3360
<< metal3 >>
rect 8109 700362 8175 700365
rect 378133 700362 378199 700365
rect 8109 700360 378199 700362
rect 8109 700304 8114 700360
rect 8170 700304 378138 700360
rect 378194 700304 378199 700360
rect 8109 700302 378199 700304
rect 8109 700299 8175 700302
rect 378133 700299 378199 700302
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 494881 686082 494947 686085
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 494237 685883 494303 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect 4889 583266 4955 583269
rect 460289 583266 460355 583269
rect 4889 583264 460355 583266
rect 4889 583208 4894 583264
rect 4950 583208 460294 583264
rect 460350 583208 460355 583264
rect 4889 583206 460355 583208
rect 4889 583203 4955 583206
rect 460289 583203 460355 583206
rect 293953 583130 294019 583133
rect 467230 583130 467236 583132
rect 293953 583128 467236 583130
rect 293953 583072 293958 583128
rect 294014 583072 467236 583128
rect 293953 583070 467236 583072
rect 293953 583067 294019 583070
rect 467230 583068 467236 583070
rect 467300 583068 467306 583132
rect 240910 582932 240916 582996
rect 240980 582994 240986 582996
rect 420269 582994 420335 582997
rect 240980 582992 420335 582994
rect 240980 582936 420274 582992
rect 420330 582936 420335 582992
rect 240980 582934 420335 582936
rect 240980 582932 240986 582934
rect 420269 582931 420335 582934
rect 240726 582796 240732 582860
rect 240796 582858 240802 582860
rect 426617 582858 426683 582861
rect 240796 582856 426683 582858
rect 240796 582800 426622 582856
rect 426678 582800 426683 582856
rect 240796 582798 426683 582800
rect 240796 582796 240802 582798
rect 426617 582795 426683 582798
rect 247677 582722 247743 582725
rect 467046 582722 467052 582724
rect 247677 582720 467052 582722
rect 247677 582664 247682 582720
rect 247738 582664 467052 582720
rect 247677 582662 467052 582664
rect 247677 582659 247743 582662
rect 467046 582660 467052 582662
rect 467116 582660 467122 582724
rect 24117 582586 24183 582589
rect 462405 582586 462471 582589
rect 24117 582584 462471 582586
rect 24117 582528 24122 582584
rect 24178 582528 462410 582584
rect 462466 582528 462471 582584
rect 24117 582526 462471 582528
rect 24117 582523 24183 582526
rect 462405 582523 462471 582526
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 231117 579322 231183 579325
rect 232957 579324 233023 579325
rect 231710 579322 231716 579324
rect 231117 579320 231716 579322
rect 231117 579264 231122 579320
rect 231178 579264 231716 579320
rect 231117 579262 231716 579264
rect 231117 579259 231183 579262
rect 231710 579260 231716 579262
rect 231780 579260 231786 579324
rect 232957 579320 233004 579324
rect 233068 579322 233074 579324
rect 235257 579322 235323 579325
rect 237189 579324 237255 579325
rect 235758 579322 235764 579324
rect 232957 579264 232962 579320
rect 232957 579260 233004 579264
rect 233068 579262 233114 579322
rect 235257 579320 235764 579322
rect 235257 579264 235262 579320
rect 235318 579264 235764 579320
rect 235257 579262 235764 579264
rect 233068 579260 233074 579262
rect 232957 579259 233023 579260
rect 235257 579259 235323 579262
rect 235758 579260 235764 579262
rect 235828 579260 235834 579324
rect 237189 579320 237236 579324
rect 237300 579322 237306 579324
rect 239397 579322 239463 579325
rect 239990 579322 239996 579324
rect 237189 579264 237194 579320
rect 237189 579260 237236 579264
rect 237300 579262 237346 579322
rect 239397 579320 239996 579322
rect 239397 579264 239402 579320
rect 239458 579264 239996 579320
rect 239397 579262 239996 579264
rect 237300 579260 237306 579262
rect 237189 579259 237255 579260
rect 239397 579259 239463 579262
rect 239990 579260 239996 579262
rect 240060 579260 240066 579324
rect 241278 579260 241284 579324
rect 241348 579322 241354 579324
rect 241421 579322 241487 579325
rect 241348 579320 241487 579322
rect 241348 579264 241426 579320
rect 241482 579264 241487 579320
rect 241348 579262 241487 579264
rect 241348 579260 241354 579262
rect 241421 579259 241487 579262
rect 243261 579324 243327 579325
rect 249517 579324 249583 579325
rect 243261 579320 243308 579324
rect 243372 579322 243378 579324
rect 243261 579264 243266 579320
rect 243261 579260 243308 579264
rect 243372 579262 243418 579322
rect 249517 579320 249564 579324
rect 249628 579322 249634 579324
rect 249517 579264 249522 579320
rect 243372 579260 243378 579262
rect 249517 579260 249564 579264
rect 249628 579262 249674 579322
rect 249628 579260 249634 579262
rect 465574 579260 465580 579324
rect 465644 579322 465650 579324
rect 468569 579322 468635 579325
rect 465644 579320 468635 579322
rect 465644 579264 468574 579320
rect 468630 579264 468635 579320
rect 465644 579262 468635 579264
rect 465644 579260 465650 579262
rect 243261 579259 243327 579260
rect 249517 579259 249583 579260
rect 468569 579259 468635 579262
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3049 567354 3115 567357
rect -960 567352 3115 567354
rect -960 567296 3054 567352
rect 3110 567296 3115 567352
rect -960 567294 3115 567296
rect -960 567204 480 567294
rect 3049 567291 3115 567294
rect 579705 557290 579771 557293
rect 583520 557290 584960 557380
rect 579705 557288 584960 557290
rect 579705 557232 579710 557288
rect 579766 557232 584960 557288
rect 579705 557230 584960 557232
rect 579705 557227 579771 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3049 553074 3115 553077
rect -960 553072 3115 553074
rect -960 553016 3054 553072
rect 3110 553016 3115 553072
rect -960 553014 3115 553016
rect -960 552924 480 553014
rect 3049 553011 3115 553014
rect 579705 545594 579771 545597
rect 583520 545594 584960 545684
rect 579705 545592 584960 545594
rect 579705 545536 579710 545592
rect 579766 545536 584960 545592
rect 579705 545534 584960 545536
rect 579705 545531 579771 545534
rect 583520 545444 584960 545534
rect -960 538658 480 538748
rect 3049 538658 3115 538661
rect -960 538656 3115 538658
rect -960 538600 3054 538656
rect 3110 538600 3115 538656
rect -960 538598 3115 538600
rect -960 538508 480 538598
rect 3049 538595 3115 538598
rect 579705 533898 579771 533901
rect 583520 533898 584960 533988
rect 579705 533896 584960 533898
rect 579705 533840 579710 533896
rect 579766 533840 584960 533896
rect 579705 533838 584960 533840
rect 579705 533835 579771 533838
rect 583520 533748 584960 533838
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 579705 510370 579771 510373
rect 583520 510370 584960 510460
rect 579705 510368 584960 510370
rect 579705 510312 579710 510368
rect 579766 510312 584960 510368
rect 579705 510310 584960 510312
rect 579705 510307 579771 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3049 509962 3115 509965
rect -960 509960 3115 509962
rect -960 509904 3054 509960
rect 3110 509904 3115 509960
rect -960 509902 3115 509904
rect -960 509812 480 509902
rect 3049 509899 3115 509902
rect 579705 498674 579771 498677
rect 583520 498674 584960 498764
rect 579705 498672 584960 498674
rect 579705 498616 579710 498672
rect 579766 498616 584960 498672
rect 579705 498614 584960 498616
rect 579705 498611 579771 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 2773 495546 2839 495549
rect -960 495544 2839 495546
rect -960 495488 2778 495544
rect 2834 495488 2839 495544
rect -960 495486 2839 495488
rect -960 495396 480 495486
rect 2773 495483 2839 495486
rect 583520 486842 584960 486932
rect 583342 486782 584960 486842
rect 467230 486100 467236 486164
rect 467300 486162 467306 486164
rect 467300 486102 470610 486162
rect 467300 486100 467306 486102
rect 470550 486026 470610 486102
rect 480302 486102 489930 486162
rect 470550 485966 480178 486026
rect 480118 485890 480178 485966
rect 480302 485890 480362 486102
rect 489870 486026 489930 486102
rect 499622 486102 509250 486162
rect 489870 485966 499498 486026
rect 480118 485830 480362 485890
rect 499438 485890 499498 485966
rect 499622 485890 499682 486102
rect 509190 486026 509250 486102
rect 518942 486102 528570 486162
rect 509190 485966 518818 486026
rect 499438 485830 499682 485890
rect 518758 485890 518818 485966
rect 518942 485890 519002 486102
rect 528510 486026 528570 486102
rect 538262 486102 547890 486162
rect 528510 485966 538138 486026
rect 518758 485830 519002 485890
rect 538078 485890 538138 485966
rect 538262 485890 538322 486102
rect 547830 486026 547890 486102
rect 557582 486102 567210 486162
rect 547830 485966 557458 486026
rect 538078 485830 538322 485890
rect 557398 485890 557458 485966
rect 557582 485890 557642 486102
rect 567150 486026 567210 486102
rect 583342 486026 583402 486782
rect 583520 486692 584960 486782
rect 567150 485966 576778 486026
rect 557398 485830 557642 485890
rect 576718 485890 576778 485966
rect 576902 485966 583402 486026
rect 576902 485890 576962 485966
rect 576718 485830 576962 485890
rect -960 481130 480 481220
rect 2957 481130 3023 481133
rect -960 481128 3023 481130
rect -960 481072 2962 481128
rect 3018 481072 3023 481128
rect -960 481070 3023 481072
rect -960 480980 480 481070
rect 2957 481067 3023 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 579705 463450 579771 463453
rect 583520 463450 584960 463540
rect 579705 463448 584960 463450
rect 579705 463392 579710 463448
rect 579766 463392 584960 463448
rect 579705 463390 584960 463392
rect 579705 463387 579771 463390
rect 583520 463300 584960 463390
rect -960 452434 480 452524
rect 3141 452434 3207 452437
rect -960 452432 3207 452434
rect -960 452376 3146 452432
rect 3202 452376 3207 452432
rect -960 452374 3207 452376
rect -960 452284 480 452374
rect 3141 452371 3207 452374
rect 579797 451754 579863 451757
rect 583520 451754 584960 451844
rect 579797 451752 584960 451754
rect 579797 451696 579802 451752
rect 579858 451696 584960 451752
rect 579797 451694 584960 451696
rect 579797 451691 579863 451694
rect 583520 451604 584960 451694
rect 579797 439922 579863 439925
rect 583520 439922 584960 440012
rect 579797 439920 584960 439922
rect 579797 439864 579802 439920
rect 579858 439864 584960 439920
rect 579797 439862 584960 439864
rect 579797 439859 579863 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3141 438018 3207 438021
rect -960 438016 3207 438018
rect -960 437960 3146 438016
rect 3202 437960 3207 438016
rect -960 437958 3207 437960
rect -960 437868 480 437958
rect 3141 437955 3207 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3141 423738 3207 423741
rect -960 423736 3207 423738
rect -960 423680 3146 423736
rect 3202 423680 3207 423736
rect -960 423678 3207 423680
rect -960 423588 480 423678
rect 3141 423675 3207 423678
rect 579797 416530 579863 416533
rect 583520 416530 584960 416620
rect 579797 416528 584960 416530
rect 579797 416472 579802 416528
rect 579858 416472 584960 416528
rect 579797 416470 584960 416472
rect 579797 416467 579863 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 579889 404834 579955 404837
rect 583520 404834 584960 404924
rect 579889 404832 584960 404834
rect 579889 404776 579894 404832
rect 579950 404776 584960 404832
rect 579889 404774 584960 404776
rect 579889 404771 579955 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 3233 395042 3299 395045
rect -960 395040 3299 395042
rect -960 394984 3238 395040
rect 3294 394984 3299 395040
rect -960 394982 3299 394984
rect -960 394892 480 394982
rect 3233 394979 3299 394982
rect 579889 393002 579955 393005
rect 583520 393002 584960 393092
rect 579889 393000 584960 393002
rect 579889 392944 579894 393000
rect 579950 392944 584960 393000
rect 579889 392942 584960 392944
rect 579889 392939 579955 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3233 380626 3299 380629
rect -960 380624 3299 380626
rect -960 380568 3238 380624
rect 3294 380568 3299 380624
rect -960 380566 3299 380568
rect -960 380476 480 380566
rect 3233 380563 3299 380566
rect 579981 369610 580047 369613
rect 583520 369610 584960 369700
rect 579981 369608 584960 369610
rect 579981 369552 579986 369608
rect 580042 369552 584960 369608
rect 579981 369550 584960 369552
rect 579981 369547 580047 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 3325 366210 3391 366213
rect -960 366208 3391 366210
rect -960 366152 3330 366208
rect 3386 366152 3391 366208
rect -960 366150 3391 366152
rect -960 366060 480 366150
rect 3325 366147 3391 366150
rect 580073 357914 580139 357917
rect 583520 357914 584960 358004
rect 580073 357912 584960 357914
rect 580073 357856 580078 357912
rect 580134 357856 584960 357912
rect 580073 357854 584960 357856
rect 580073 357851 580139 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 579797 346082 579863 346085
rect 583520 346082 584960 346172
rect 579797 346080 584960 346082
rect 579797 346024 579802 346080
rect 579858 346024 584960 346080
rect 579797 346022 584960 346024
rect 579797 346019 579863 346022
rect 583520 345932 584960 346022
rect 242934 340580 242940 340644
rect 243004 340642 243010 340644
rect 249558 340642 249564 340644
rect 243004 340582 249564 340642
rect 243004 340580 243010 340582
rect 249558 340580 249564 340582
rect 249628 340580 249634 340644
rect 240910 338058 240916 338060
rect 614 337998 240916 338058
rect -960 337514 480 337604
rect 614 337514 674 337998
rect 240910 337996 240916 337998
rect 240980 337996 240986 338060
rect 376753 338058 376819 338061
rect 379329 338058 379395 338061
rect 376753 338056 379395 338058
rect 376753 338000 376758 338056
rect 376814 338000 379334 338056
rect 379390 338000 379395 338056
rect 376753 337998 379395 338000
rect 376753 337995 376819 337998
rect 379329 337995 379395 337998
rect -960 337454 674 337514
rect -960 337364 480 337454
rect 10317 337378 10383 337381
rect 231945 337378 232011 337381
rect 10317 337376 232011 337378
rect 10317 337320 10322 337376
rect 10378 337320 231950 337376
rect 232006 337320 232011 337376
rect 10317 337318 232011 337320
rect 10317 337315 10383 337318
rect 231945 337315 232011 337318
rect 467557 337378 467623 337381
rect 512637 337378 512703 337381
rect 467557 337376 512703 337378
rect 467557 337320 467562 337376
rect 467618 337320 512642 337376
rect 512698 337320 512703 337376
rect 467557 337318 512703 337320
rect 467557 337315 467623 337318
rect 512637 337315 512703 337318
rect 132493 337242 132559 337245
rect 142061 337242 142127 337245
rect 132493 337240 142127 337242
rect 132493 337184 132498 337240
rect 132554 337184 142066 337240
rect 142122 337184 142127 337240
rect 132493 337182 142127 337184
rect 132493 337179 132559 337182
rect 142061 337179 142127 337182
rect 151813 337242 151879 337245
rect 161381 337242 161447 337245
rect 151813 337240 161447 337242
rect 151813 337184 151818 337240
rect 151874 337184 161386 337240
rect 161442 337184 161447 337240
rect 151813 337182 161447 337184
rect 151813 337179 151879 337182
rect 161381 337179 161447 337182
rect 171133 337242 171199 337245
rect 180701 337242 180767 337245
rect 171133 337240 180767 337242
rect 171133 337184 171138 337240
rect 171194 337184 180706 337240
rect 180762 337184 180767 337240
rect 171133 337182 180767 337184
rect 171133 337179 171199 337182
rect 180701 337179 180767 337182
rect 190453 337242 190519 337245
rect 200021 337242 200087 337245
rect 190453 337240 200087 337242
rect 190453 337184 190458 337240
rect 190514 337184 200026 337240
rect 200082 337184 200087 337240
rect 190453 337182 200087 337184
rect 190453 337179 190519 337182
rect 200021 337179 200087 337182
rect 209773 337242 209839 337245
rect 219341 337242 219407 337245
rect 209773 337240 219407 337242
rect 209773 337184 209778 337240
rect 209834 337184 219346 337240
rect 219402 337184 219407 337240
rect 209773 337182 219407 337184
rect 209773 337179 209839 337182
rect 219341 337179 219407 337182
rect 229185 337242 229251 337245
rect 234613 337242 234679 337245
rect 229185 337240 234679 337242
rect 229185 337184 229190 337240
rect 229246 337184 234618 337240
rect 234674 337184 234679 337240
rect 229185 337182 234679 337184
rect 229185 337179 229251 337182
rect 234613 337179 234679 337182
rect 470501 337242 470567 337245
rect 470685 337242 470751 337245
rect 470501 337240 470751 337242
rect 470501 337184 470506 337240
rect 470562 337184 470690 337240
rect 470746 337184 470751 337240
rect 470501 337182 470751 337184
rect 470501 337179 470567 337182
rect 470685 337179 470751 337182
rect 249241 336698 249307 336701
rect 249558 336698 249564 336700
rect 249241 336696 249564 336698
rect 249241 336640 249246 336696
rect 249302 336640 249564 336696
rect 249241 336638 249564 336640
rect 249241 336635 249307 336638
rect 249558 336636 249564 336638
rect 249628 336636 249634 336700
rect 583520 334236 584960 334476
rect 360929 327314 360995 327317
rect 360334 327312 360995 327314
rect 360334 327256 360934 327312
rect 360990 327256 360995 327312
rect 360334 327254 360995 327256
rect 249241 327178 249307 327181
rect 249374 327178 249380 327180
rect 249241 327176 249380 327178
rect 249241 327120 249246 327176
rect 249302 327120 249380 327176
rect 249241 327118 249380 327120
rect 249241 327115 249307 327118
rect 249374 327116 249380 327118
rect 249444 327116 249450 327180
rect 360334 327178 360394 327254
rect 360929 327251 360995 327254
rect 360469 327178 360535 327181
rect 360334 327176 360535 327178
rect 360334 327120 360474 327176
rect 360530 327120 360535 327176
rect 360334 327118 360535 327120
rect 360469 327115 360535 327118
rect 579981 325682 580047 325685
rect 580901 325682 580967 325685
rect 579981 325680 580967 325682
rect 579981 325624 579986 325680
rect 580042 325624 580906 325680
rect 580962 325624 580967 325680
rect 579981 325622 580967 325624
rect 579981 325619 580047 325622
rect 580901 325619 580967 325622
rect -960 323098 480 323188
rect 3325 323098 3391 323101
rect -960 323096 3391 323098
rect -960 323040 3330 323096
rect 3386 323040 3391 323096
rect -960 323038 3391 323040
rect -960 322948 480 323038
rect 3325 323035 3391 323038
rect 580073 322690 580139 322693
rect 583520 322690 584960 322780
rect 580073 322688 584960 322690
rect 580073 322632 580078 322688
rect 580134 322632 584960 322688
rect 580073 322630 584960 322632
rect 580073 322627 580139 322630
rect 583520 322540 584960 322630
rect 249241 321466 249307 321469
rect 249374 321466 249380 321468
rect 249241 321464 249380 321466
rect 249241 321408 249246 321464
rect 249302 321408 249380 321464
rect 249241 321406 249380 321408
rect 249241 321403 249307 321406
rect 249374 321404 249380 321406
rect 249444 321404 249450 321468
rect 376845 318882 376911 318885
rect 377121 318882 377187 318885
rect 376845 318880 377187 318882
rect 376845 318824 376850 318880
rect 376906 318824 377126 318880
rect 377182 318824 377187 318880
rect 376845 318822 377187 318824
rect 376845 318819 376911 318822
rect 377121 318819 377187 318822
rect 249241 317658 249307 317661
rect 249014 317656 249307 317658
rect 249014 317600 249246 317656
rect 249302 317600 249307 317656
rect 249014 317598 249307 317600
rect 249014 317524 249074 317598
rect 249241 317595 249307 317598
rect 249006 317460 249012 317524
rect 249076 317460 249082 317524
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect 249006 309164 249012 309228
rect 249076 309164 249082 309228
rect 249014 308954 249074 309164
rect 249190 308954 249196 308956
rect -960 308818 480 308908
rect 249014 308894 249196 308954
rect 249190 308892 249196 308894
rect 249260 308892 249266 308956
rect 2773 308818 2839 308821
rect -960 308816 2839 308818
rect -960 308760 2778 308816
rect 2834 308760 2839 308816
rect -960 308758 2839 308760
rect -960 308668 480 308758
rect 2773 308755 2839 308758
rect 284753 306370 284819 306373
rect 284937 306370 285003 306373
rect 284753 306368 285003 306370
rect 284753 306312 284758 306368
rect 284814 306312 284942 306368
rect 284998 306312 285003 306368
rect 284753 306310 285003 306312
rect 284753 306307 284819 306310
rect 284937 306307 285003 306310
rect 301221 306370 301287 306373
rect 301405 306370 301471 306373
rect 301221 306368 301471 306370
rect 301221 306312 301226 306368
rect 301282 306312 301410 306368
rect 301466 306312 301471 306368
rect 301221 306310 301471 306312
rect 301221 306307 301287 306310
rect 301405 306307 301471 306310
rect 580073 306370 580139 306373
rect 580901 306370 580967 306373
rect 580073 306368 580967 306370
rect 580073 306312 580078 306368
rect 580134 306312 580906 306368
rect 580962 306312 580967 306368
rect 580073 306310 580967 306312
rect 580073 306307 580139 306310
rect 580901 306307 580967 306310
rect 249190 302228 249196 302292
rect 249260 302228 249266 302292
rect 249198 302156 249258 302228
rect 249190 302092 249196 302156
rect 249260 302092 249266 302156
rect 580165 299162 580231 299165
rect 583520 299162 584960 299252
rect 580165 299160 584960 299162
rect 580165 299104 580170 299160
rect 580226 299104 584960 299160
rect 580165 299102 584960 299104
rect 580165 299099 580231 299102
rect 583520 299012 584960 299102
rect 249241 298076 249307 298077
rect 249190 298074 249196 298076
rect 249150 298014 249196 298074
rect 249260 298072 249307 298076
rect 249302 298016 249307 298072
rect 249190 298012 249196 298014
rect 249260 298012 249307 298016
rect 249241 298011 249307 298012
rect 284661 296714 284727 296717
rect 284845 296714 284911 296717
rect 284661 296712 284911 296714
rect 284661 296656 284666 296712
rect 284722 296656 284850 296712
rect 284906 296656 284911 296712
rect 284661 296654 284911 296656
rect 284661 296651 284727 296654
rect 284845 296651 284911 296654
rect 330109 296714 330175 296717
rect 330661 296714 330727 296717
rect 330109 296712 330727 296714
rect 330109 296656 330114 296712
rect 330170 296656 330666 296712
rect 330722 296656 330727 296712
rect 330109 296654 330727 296656
rect 330109 296651 330175 296654
rect 330661 296651 330727 296654
rect 2957 295218 3023 295221
rect 240726 295218 240732 295220
rect 2957 295216 240732 295218
rect 2957 295160 2962 295216
rect 3018 295160 240732 295216
rect 2957 295158 240732 295160
rect 2957 295155 3023 295158
rect 240726 295156 240732 295158
rect 240796 295156 240802 295220
rect -960 294402 480 294492
rect 2957 294402 3023 294405
rect -960 294400 3023 294402
rect -960 294344 2962 294400
rect 3018 294344 3023 294400
rect -960 294342 3023 294344
rect -960 294252 480 294342
rect 2957 294339 3023 294342
rect 270769 293994 270835 293997
rect 270953 293994 271019 293997
rect 270769 293992 271019 293994
rect 270769 293936 270774 293992
rect 270830 293936 270958 293992
rect 271014 293936 271019 293992
rect 270769 293934 271019 293936
rect 270769 293931 270835 293934
rect 270953 293931 271019 293934
rect 249241 288554 249307 288557
rect 249374 288554 249380 288556
rect 249241 288552 249380 288554
rect 249241 288496 249246 288552
rect 249302 288496 249380 288552
rect 249241 288494 249380 288496
rect 249241 288491 249307 288494
rect 249374 288492 249380 288494
rect 249444 288492 249450 288556
rect 249241 288418 249307 288421
rect 249374 288418 249380 288420
rect 249241 288416 249380 288418
rect 249241 288360 249246 288416
rect 249302 288360 249380 288416
rect 249241 288358 249380 288360
rect 249241 288355 249307 288358
rect 249374 288356 249380 288358
rect 249444 288356 249450 288420
rect 250069 288418 250135 288421
rect 250345 288418 250411 288421
rect 250069 288416 250411 288418
rect 250069 288360 250074 288416
rect 250130 288360 250350 288416
rect 250406 288360 250411 288416
rect 250069 288358 250411 288360
rect 250069 288355 250135 288358
rect 250345 288355 250411 288358
rect 583520 287316 584960 287556
rect 337101 287058 337167 287061
rect 337285 287058 337351 287061
rect 337101 287056 337351 287058
rect 337101 287000 337106 287056
rect 337162 287000 337290 287056
rect 337346 287000 337351 287056
rect 337101 286998 337351 287000
rect 337101 286995 337167 286998
rect 337285 286995 337351 286998
rect 302509 285698 302575 285701
rect 302693 285698 302759 285701
rect 302509 285696 302759 285698
rect 302509 285640 302514 285696
rect 302570 285640 302698 285696
rect 302754 285640 302759 285696
rect 302509 285638 302759 285640
rect 302509 285635 302575 285638
rect 302693 285635 302759 285638
rect 259545 280258 259611 280261
rect 259913 280258 259979 280261
rect 259545 280256 259979 280258
rect -960 280122 480 280212
rect 259545 280200 259550 280256
rect 259606 280200 259918 280256
rect 259974 280200 259979 280256
rect 259545 280198 259979 280200
rect 259545 280195 259611 280198
rect 259913 280195 259979 280198
rect 4061 280122 4127 280125
rect -960 280120 4127 280122
rect -960 280064 4066 280120
rect 4122 280064 4127 280120
rect -960 280062 4127 280064
rect -960 279972 480 280062
rect 4061 280059 4127 280062
rect 249241 279036 249307 279037
rect 249190 279034 249196 279036
rect 249150 278974 249196 279034
rect 249260 279032 249307 279036
rect 249302 278976 249307 279032
rect 249190 278972 249196 278974
rect 249260 278972 249307 278976
rect 249241 278971 249307 278972
rect 323485 278762 323551 278765
rect 323669 278762 323735 278765
rect 323485 278760 323735 278762
rect 323485 278704 323490 278760
rect 323546 278704 323674 278760
rect 323730 278704 323735 278760
rect 323485 278702 323735 278704
rect 323485 278699 323551 278702
rect 323669 278699 323735 278702
rect 358537 278762 358603 278765
rect 358721 278762 358787 278765
rect 358537 278760 358787 278762
rect 358537 278704 358542 278760
rect 358598 278704 358726 278760
rect 358782 278704 358787 278760
rect 358537 278702 358787 278704
rect 358537 278699 358603 278702
rect 358721 278699 358787 278702
rect 249190 277340 249196 277404
rect 249260 277402 249266 277404
rect 249425 277402 249491 277405
rect 249260 277400 249491 277402
rect 249260 277344 249430 277400
rect 249486 277344 249491 277400
rect 249260 277342 249491 277344
rect 249260 277340 249266 277342
rect 249425 277339 249491 277342
rect 265249 277402 265315 277405
rect 265433 277402 265499 277405
rect 265249 277400 265499 277402
rect 265249 277344 265254 277400
rect 265310 277344 265438 277400
rect 265494 277344 265499 277400
rect 265249 277342 265499 277344
rect 265249 277339 265315 277342
rect 265433 277339 265499 277342
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 266813 270602 266879 270605
rect 266678 270600 266879 270602
rect 266678 270544 266818 270600
rect 266874 270544 266879 270600
rect 266678 270542 266879 270544
rect 266678 270469 266738 270542
rect 266813 270539 266879 270542
rect 266629 270464 266738 270469
rect 266629 270408 266634 270464
rect 266690 270408 266738 270464
rect 266629 270406 266738 270408
rect 266629 270403 266695 270406
rect 284569 269106 284635 269109
rect 284753 269106 284819 269109
rect 284569 269104 284819 269106
rect 284569 269048 284574 269104
rect 284630 269048 284758 269104
rect 284814 269048 284819 269104
rect 284569 269046 284819 269048
rect 284569 269043 284635 269046
rect 284753 269043 284819 269046
rect 330201 269106 330267 269109
rect 330385 269106 330451 269109
rect 330201 269104 330451 269106
rect 330201 269048 330206 269104
rect 330262 269048 330390 269104
rect 330446 269048 330451 269104
rect 330201 269046 330451 269048
rect 330201 269043 330267 269046
rect 330385 269043 330451 269046
rect 249425 267884 249491 267885
rect 249374 267820 249380 267884
rect 249444 267882 249491 267884
rect 249444 267880 249536 267882
rect 249486 267824 249536 267880
rect 249444 267822 249536 267824
rect 249444 267820 249491 267822
rect 249425 267819 249491 267820
rect 294137 267746 294203 267749
rect 294094 267744 294203 267746
rect 294094 267688 294142 267744
rect 294198 267688 294203 267744
rect 294094 267683 294203 267688
rect 294094 267610 294154 267683
rect 294229 267610 294295 267613
rect 294094 267608 294295 267610
rect 294094 267552 294234 267608
rect 294290 267552 294295 267608
rect 294094 267550 294295 267552
rect 294229 267547 294295 267550
rect 302509 266386 302575 266389
rect 302785 266386 302851 266389
rect 302509 266384 302851 266386
rect 302509 266328 302514 266384
rect 302570 266328 302790 266384
rect 302846 266328 302851 266384
rect 302509 266326 302851 266328
rect 302509 266323 302575 266326
rect 302785 266323 302851 266326
rect 306649 266386 306715 266389
rect 306833 266386 306899 266389
rect 306649 266384 306899 266386
rect 306649 266328 306654 266384
rect 306710 266328 306838 266384
rect 306894 266328 306899 266384
rect 306649 266326 306899 266328
rect 306649 266323 306715 266326
rect 306833 266323 306899 266326
rect -960 265706 480 265796
rect 3969 265706 4035 265709
rect -960 265704 4035 265706
rect -960 265648 3974 265704
rect 4030 265648 4035 265704
rect -960 265646 4035 265648
rect -960 265556 480 265646
rect 3969 265643 4035 265646
rect 580809 263938 580875 263941
rect 583520 263938 584960 264028
rect 580809 263936 584960 263938
rect 580809 263880 580814 263936
rect 580870 263880 584960 263936
rect 580809 263878 584960 263880
rect 580809 263875 580875 263878
rect 249374 263802 249380 263804
rect 249198 263742 249380 263802
rect 249198 263532 249258 263742
rect 249374 263740 249380 263742
rect 249444 263740 249450 263804
rect 583520 263788 584960 263878
rect 249190 263468 249196 263532
rect 249260 263468 249266 263532
rect 286041 261082 286107 261085
rect 285814 261080 286107 261082
rect 285814 261024 286046 261080
rect 286102 261024 286107 261080
rect 285814 261022 286107 261024
rect 285814 260946 285874 261022
rect 286041 261019 286107 261022
rect 285949 260946 286015 260949
rect 285814 260944 286015 260946
rect 285814 260888 285954 260944
rect 286010 260888 286015 260944
rect 285814 260886 286015 260888
rect 285949 260883 286015 260886
rect 341057 260946 341123 260949
rect 341425 260946 341491 260949
rect 341057 260944 341491 260946
rect 341057 260888 341062 260944
rect 341118 260888 341430 260944
rect 341486 260888 341491 260944
rect 341057 260886 341491 260888
rect 341057 260883 341123 260886
rect 341425 260883 341491 260886
rect 244457 259450 244523 259453
rect 244641 259450 244707 259453
rect 244457 259448 244707 259450
rect 244457 259392 244462 259448
rect 244518 259392 244646 259448
rect 244702 259392 244707 259448
rect 244457 259390 244707 259392
rect 244457 259387 244523 259390
rect 244641 259387 244707 259390
rect 265157 259450 265223 259453
rect 265341 259450 265407 259453
rect 265157 259448 265407 259450
rect 265157 259392 265162 259448
rect 265218 259392 265346 259448
rect 265402 259392 265407 259448
rect 265157 259390 265407 259392
rect 265157 259387 265223 259390
rect 265341 259387 265407 259390
rect 267733 259450 267799 259453
rect 267917 259450 267983 259453
rect 267733 259448 267983 259450
rect 267733 259392 267738 259448
rect 267794 259392 267922 259448
rect 267978 259392 267983 259448
rect 267733 259390 267983 259392
rect 267733 259387 267799 259390
rect 267917 259387 267983 259390
rect 323209 259450 323275 259453
rect 323393 259450 323459 259453
rect 323209 259448 323459 259450
rect 323209 259392 323214 259448
rect 323270 259392 323398 259448
rect 323454 259392 323459 259448
rect 323209 259390 323459 259392
rect 323209 259387 323275 259390
rect 323393 259387 323459 259390
rect 358537 259450 358603 259453
rect 358721 259450 358787 259453
rect 358537 259448 358787 259450
rect 358537 259392 358542 259448
rect 358598 259392 358726 259448
rect 358782 259392 358787 259448
rect 358537 259390 358787 259392
rect 358537 259387 358603 259390
rect 358721 259387 358787 259390
rect 291561 258226 291627 258229
rect 291518 258224 291627 258226
rect 291518 258168 291566 258224
rect 291622 258168 291627 258224
rect 291518 258163 291627 258168
rect 291518 258093 291578 258163
rect 291469 258088 291578 258093
rect 291469 258032 291474 258088
rect 291530 258032 291578 258088
rect 291469 258030 291578 258032
rect 295609 258090 295675 258093
rect 295793 258090 295859 258093
rect 295609 258088 295859 258090
rect 295609 258032 295614 258088
rect 295670 258032 295798 258088
rect 295854 258032 295859 258088
rect 295609 258030 295859 258032
rect 291469 258027 291535 258030
rect 295609 258027 295675 258030
rect 295793 258027 295859 258030
rect 296805 258090 296871 258093
rect 296989 258090 297055 258093
rect 296805 258088 297055 258090
rect 296805 258032 296810 258088
rect 296866 258032 296994 258088
rect 297050 258032 297055 258088
rect 296805 258030 297055 258032
rect 296805 258027 296871 258030
rect 296989 258027 297055 258030
rect 302509 258090 302575 258093
rect 302785 258090 302851 258093
rect 302509 258088 302851 258090
rect 302509 258032 302514 258088
rect 302570 258032 302790 258088
rect 302846 258032 302851 258088
rect 302509 258030 302851 258032
rect 302509 258027 302575 258030
rect 302785 258027 302851 258030
rect 337009 256730 337075 256733
rect 337193 256730 337259 256733
rect 337009 256728 337259 256730
rect 337009 256672 337014 256728
rect 337070 256672 337198 256728
rect 337254 256672 337259 256728
rect 337009 256670 337259 256672
rect 337009 256667 337075 256670
rect 337193 256667 337259 256670
rect 579613 252242 579679 252245
rect 583520 252242 584960 252332
rect 579613 252240 584960 252242
rect 579613 252184 579618 252240
rect 579674 252184 584960 252240
rect 579613 252182 584960 252184
rect 579613 252179 579679 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 2773 251290 2839 251293
rect -960 251288 2839 251290
rect -960 251232 2778 251288
rect 2834 251232 2839 251288
rect -960 251230 2839 251232
rect -960 251140 480 251230
rect 2773 251227 2839 251230
rect 236269 251154 236335 251157
rect 236453 251154 236519 251157
rect 236269 251152 236519 251154
rect 236269 251096 236274 251152
rect 236330 251096 236458 251152
rect 236514 251096 236519 251152
rect 236269 251094 236519 251096
rect 236269 251091 236335 251094
rect 236453 251091 236519 251094
rect 388989 251154 389055 251157
rect 389173 251154 389239 251157
rect 388989 251152 389239 251154
rect 388989 251096 388994 251152
rect 389050 251096 389178 251152
rect 389234 251096 389239 251152
rect 388989 251094 389239 251096
rect 388989 251091 389055 251094
rect 389173 251091 389239 251094
rect 284661 249794 284727 249797
rect 284937 249794 285003 249797
rect 286041 249794 286107 249797
rect 299841 249794 299907 249797
rect 284661 249792 285003 249794
rect 284661 249736 284666 249792
rect 284722 249736 284942 249792
rect 284998 249736 285003 249792
rect 284661 249734 285003 249736
rect 284661 249731 284727 249734
rect 284937 249731 285003 249734
rect 285998 249792 286107 249794
rect 285998 249736 286046 249792
rect 286102 249736 286107 249792
rect 285998 249731 286107 249736
rect 299798 249792 299907 249794
rect 299798 249736 299846 249792
rect 299902 249736 299907 249792
rect 299798 249731 299907 249736
rect 285998 249661 286058 249731
rect 285949 249656 286058 249661
rect 285949 249600 285954 249656
rect 286010 249600 286058 249656
rect 285949 249598 286058 249600
rect 299798 249658 299858 249731
rect 299933 249658 299999 249661
rect 299798 249656 299999 249658
rect 299798 249600 299938 249656
rect 299994 249600 299999 249656
rect 299798 249598 299999 249600
rect 285949 249595 286015 249598
rect 299933 249595 299999 249598
rect 264973 248434 265039 248437
rect 265157 248434 265223 248437
rect 264973 248432 265223 248434
rect 264973 248376 264978 248432
rect 265034 248376 265162 248432
rect 265218 248376 265223 248432
rect 264973 248374 265223 248376
rect 264973 248371 265039 248374
rect 265157 248371 265223 248374
rect 267733 248434 267799 248437
rect 268101 248434 268167 248437
rect 267733 248432 268167 248434
rect 267733 248376 267738 248432
rect 267794 248376 268106 248432
rect 268162 248376 268167 248432
rect 267733 248374 268167 248376
rect 267733 248371 267799 248374
rect 268101 248371 268167 248374
rect 291469 248434 291535 248437
rect 291837 248434 291903 248437
rect 291469 248432 291903 248434
rect 291469 248376 291474 248432
rect 291530 248376 291842 248432
rect 291898 248376 291903 248432
rect 291469 248374 291903 248376
rect 291469 248371 291535 248374
rect 291837 248371 291903 248374
rect 295241 248434 295307 248437
rect 295517 248434 295583 248437
rect 295241 248432 295583 248434
rect 295241 248376 295246 248432
rect 295302 248376 295522 248432
rect 295578 248376 295583 248432
rect 295241 248374 295583 248376
rect 295241 248371 295307 248374
rect 295517 248371 295583 248374
rect 329925 248434 329991 248437
rect 330293 248434 330359 248437
rect 329925 248432 330359 248434
rect 329925 248376 329930 248432
rect 329986 248376 330298 248432
rect 330354 248376 330359 248432
rect 329925 248374 330359 248376
rect 329925 248371 329991 248374
rect 330293 248371 330359 248374
rect 249374 241906 249380 241908
rect 249198 241846 249380 241906
rect 249198 241772 249258 241846
rect 249374 241844 249380 241846
rect 249444 241844 249450 241908
rect 249190 241708 249196 241772
rect 249260 241708 249266 241772
rect 244273 241498 244339 241501
rect 244457 241498 244523 241501
rect 244273 241496 244523 241498
rect 244273 241440 244278 241496
rect 244334 241440 244462 241496
rect 244518 241440 244523 241496
rect 244273 241438 244523 241440
rect 244273 241435 244339 241438
rect 244457 241435 244523 241438
rect 249190 241436 249196 241500
rect 249260 241436 249266 241500
rect 251449 241498 251515 241501
rect 251633 241498 251699 241501
rect 251449 241496 251699 241498
rect 251449 241440 251454 241496
rect 251510 241440 251638 241496
rect 251694 241440 251699 241496
rect 251449 241438 251699 241440
rect 249198 240954 249258 241436
rect 251449 241435 251515 241438
rect 251633 241435 251699 241438
rect 338665 241498 338731 241501
rect 338849 241498 338915 241501
rect 367001 241500 367067 241501
rect 366950 241498 366956 241500
rect 338665 241496 338915 241498
rect 338665 241440 338670 241496
rect 338726 241440 338854 241496
rect 338910 241440 338915 241496
rect 338665 241438 338915 241440
rect 366910 241438 366956 241498
rect 367020 241496 367067 241500
rect 367062 241440 367067 241496
rect 338665 241435 338731 241438
rect 338849 241435 338915 241438
rect 366950 241436 366956 241438
rect 367020 241436 367067 241440
rect 367001 241435 367067 241436
rect 372521 241498 372587 241501
rect 372705 241498 372771 241501
rect 372521 241496 372771 241498
rect 372521 241440 372526 241496
rect 372582 241440 372710 241496
rect 372766 241440 372771 241496
rect 372521 241438 372771 241440
rect 372521 241435 372587 241438
rect 372705 241435 372771 241438
rect 376937 241498 377003 241501
rect 377121 241498 377187 241501
rect 376937 241496 377187 241498
rect 376937 241440 376942 241496
rect 376998 241440 377126 241496
rect 377182 241440 377187 241496
rect 376937 241438 377187 241440
rect 376937 241435 377003 241438
rect 377121 241435 377187 241438
rect 249374 240954 249380 240956
rect 249198 240894 249380 240954
rect 249374 240892 249380 240894
rect 249444 240892 249450 240956
rect 583520 240396 584960 240636
rect 270677 240138 270743 240141
rect 270542 240136 270743 240138
rect 270542 240080 270682 240136
rect 270738 240080 270743 240136
rect 270542 240078 270743 240080
rect 270542 240002 270602 240078
rect 270677 240075 270743 240078
rect 290181 240138 290247 240141
rect 290365 240138 290431 240141
rect 290181 240136 290431 240138
rect 290181 240080 290186 240136
rect 290242 240080 290370 240136
rect 290426 240080 290431 240136
rect 290181 240078 290431 240080
rect 290181 240075 290247 240078
rect 290365 240075 290431 240078
rect 358537 240138 358603 240141
rect 358721 240138 358787 240141
rect 358537 240136 358787 240138
rect 358537 240080 358542 240136
rect 358598 240080 358726 240136
rect 358782 240080 358787 240136
rect 358537 240078 358787 240080
rect 358537 240075 358603 240078
rect 358721 240075 358787 240078
rect 270677 240002 270743 240005
rect 270542 240000 270743 240002
rect 270542 239944 270682 240000
rect 270738 239944 270743 240000
rect 270542 239942 270743 239944
rect 270677 239939 270743 239942
rect 288893 238912 288959 238917
rect 288893 238856 288898 238912
rect 288954 238856 288959 238912
rect 288893 238851 288959 238856
rect 288896 238506 288956 238851
rect 295609 238778 295675 238781
rect 295793 238778 295859 238781
rect 295609 238776 295859 238778
rect 295609 238720 295614 238776
rect 295670 238720 295798 238776
rect 295854 238720 295859 238776
rect 295609 238718 295859 238720
rect 295609 238715 295675 238718
rect 295793 238715 295859 238718
rect 289077 238506 289143 238509
rect 288896 238504 289143 238506
rect 288896 238448 289082 238504
rect 289138 238448 289143 238504
rect 288896 238446 289143 238448
rect 289077 238443 289143 238446
rect -960 237010 480 237100
rect 3049 237010 3115 237013
rect -960 237008 3115 237010
rect -960 236952 3054 237008
rect 3110 236952 3115 237008
rect -960 236950 3115 236952
rect -960 236860 480 236950
rect 3049 236947 3115 236950
rect 367001 231980 367067 231981
rect 366950 231978 366956 231980
rect 366910 231918 366956 231978
rect 367020 231976 367067 231980
rect 367062 231920 367067 231976
rect 366950 231916 366956 231918
rect 367020 231916 367067 231920
rect 367001 231915 367067 231916
rect 236269 231842 236335 231845
rect 236453 231842 236519 231845
rect 325969 231842 326035 231845
rect 236269 231840 236519 231842
rect 236269 231784 236274 231840
rect 236330 231784 236458 231840
rect 236514 231784 236519 231840
rect 236269 231782 236519 231784
rect 236269 231779 236335 231782
rect 236453 231779 236519 231782
rect 325926 231840 326035 231842
rect 325926 231784 325974 231840
rect 326030 231784 326035 231840
rect 325926 231779 326035 231784
rect 389265 231842 389331 231845
rect 389449 231842 389515 231845
rect 389265 231840 389515 231842
rect 389265 231784 389270 231840
rect 389326 231784 389454 231840
rect 389510 231784 389515 231840
rect 389265 231782 389515 231784
rect 389265 231779 389331 231782
rect 389449 231779 389515 231782
rect 463785 231842 463851 231845
rect 463969 231842 464035 231845
rect 463785 231840 464035 231842
rect 463785 231784 463790 231840
rect 463846 231784 463974 231840
rect 464030 231784 464035 231840
rect 463785 231782 464035 231784
rect 463785 231779 463851 231782
rect 463969 231779 464035 231782
rect 470409 231842 470475 231845
rect 470593 231842 470659 231845
rect 470409 231840 470659 231842
rect 470409 231784 470414 231840
rect 470470 231784 470598 231840
rect 470654 231784 470659 231840
rect 470409 231782 470659 231784
rect 470409 231779 470475 231782
rect 470593 231779 470659 231782
rect 325926 231706 325986 231779
rect 326061 231706 326127 231709
rect 325926 231704 326127 231706
rect 325926 231648 326066 231704
rect 326122 231648 326127 231704
rect 325926 231646 326127 231648
rect 326061 231643 326127 231646
rect 272241 230482 272307 230485
rect 272425 230482 272491 230485
rect 272241 230480 272491 230482
rect 272241 230424 272246 230480
rect 272302 230424 272430 230480
rect 272486 230424 272491 230480
rect 272241 230422 272491 230424
rect 272241 230419 272307 230422
rect 272425 230419 272491 230422
rect 580717 228850 580783 228853
rect 583520 228850 584960 228940
rect 580717 228848 584960 228850
rect 580717 228792 580722 228848
rect 580778 228792 584960 228848
rect 580717 228790 584960 228792
rect 580717 228787 580783 228790
rect 583520 228700 584960 228790
rect 249374 224980 249380 225044
rect 249444 224980 249450 225044
rect 249382 224770 249442 224980
rect 249558 224770 249564 224772
rect 249382 224710 249564 224770
rect 249558 224708 249564 224710
rect 249628 224708 249634 224772
rect -960 222594 480 222684
rect 3877 222594 3943 222597
rect -960 222592 3943 222594
rect -960 222536 3882 222592
rect 3938 222536 3943 222592
rect -960 222534 3943 222536
rect -960 222444 480 222534
rect 3877 222531 3943 222534
rect 244273 222186 244339 222189
rect 244457 222186 244523 222189
rect 244273 222184 244523 222186
rect 244273 222128 244278 222184
rect 244334 222128 244462 222184
rect 244518 222128 244523 222184
rect 244273 222126 244523 222128
rect 244273 222123 244339 222126
rect 244457 222123 244523 222126
rect 251449 222186 251515 222189
rect 251633 222186 251699 222189
rect 251449 222184 251699 222186
rect 251449 222128 251454 222184
rect 251510 222128 251638 222184
rect 251694 222128 251699 222184
rect 251449 222126 251699 222128
rect 251449 222123 251515 222126
rect 251633 222123 251699 222126
rect 285949 222186 286015 222189
rect 286133 222186 286199 222189
rect 285949 222184 286199 222186
rect 285949 222128 285954 222184
rect 286010 222128 286138 222184
rect 286194 222128 286199 222184
rect 285949 222126 286199 222128
rect 285949 222123 286015 222126
rect 286133 222123 286199 222126
rect 331397 222186 331463 222189
rect 331581 222186 331647 222189
rect 331397 222184 331647 222186
rect 331397 222128 331402 222184
rect 331458 222128 331586 222184
rect 331642 222128 331647 222184
rect 331397 222126 331647 222128
rect 331397 222123 331463 222126
rect 331581 222123 331647 222126
rect 338665 222186 338731 222189
rect 338849 222186 338915 222189
rect 338665 222184 338915 222186
rect 338665 222128 338670 222184
rect 338726 222128 338854 222184
rect 338910 222128 338915 222184
rect 338665 222126 338915 222128
rect 338665 222123 338731 222126
rect 338849 222123 338915 222126
rect 372521 222186 372587 222189
rect 372705 222186 372771 222189
rect 372521 222184 372771 222186
rect 372521 222128 372526 222184
rect 372582 222128 372710 222184
rect 372766 222128 372771 222184
rect 372521 222126 372771 222128
rect 372521 222123 372587 222126
rect 372705 222123 372771 222126
rect 376937 222186 377003 222189
rect 377121 222186 377187 222189
rect 376937 222184 377187 222186
rect 376937 222128 376942 222184
rect 376998 222128 377126 222184
rect 377182 222128 377187 222184
rect 376937 222126 377187 222128
rect 376937 222123 377003 222126
rect 377121 222123 377187 222126
rect 285949 220826 286015 220829
rect 286133 220826 286199 220829
rect 285949 220824 286199 220826
rect 285949 220768 285954 220824
rect 286010 220768 286138 220824
rect 286194 220768 286199 220824
rect 285949 220766 286199 220768
rect 285949 220763 286015 220766
rect 286133 220763 286199 220766
rect 329925 220826 329991 220829
rect 330201 220826 330267 220829
rect 329925 220824 330267 220826
rect 329925 220768 329930 220824
rect 329986 220768 330206 220824
rect 330262 220768 330267 220824
rect 329925 220766 330267 220768
rect 329925 220763 329991 220766
rect 330201 220763 330267 220766
rect 357433 220826 357499 220829
rect 357617 220826 357683 220829
rect 357433 220824 357683 220826
rect 357433 220768 357438 220824
rect 357494 220768 357622 220824
rect 357678 220768 357683 220824
rect 357433 220766 357683 220768
rect 357433 220763 357499 220766
rect 357617 220763 357683 220766
rect 358537 220826 358603 220829
rect 358721 220826 358787 220829
rect 358537 220824 358787 220826
rect 358537 220768 358542 220824
rect 358598 220768 358726 220824
rect 358782 220768 358787 220824
rect 358537 220766 358787 220768
rect 358537 220763 358603 220766
rect 358721 220763 358787 220766
rect 249190 217364 249196 217428
rect 249260 217426 249266 217428
rect 249558 217426 249564 217428
rect 249260 217366 249564 217426
rect 249260 217364 249266 217366
rect 249558 217364 249564 217366
rect 249628 217364 249634 217428
rect 580625 217018 580691 217021
rect 583520 217018 584960 217108
rect 580625 217016 584960 217018
rect 580625 216960 580630 217016
rect 580686 216960 584960 217016
rect 580625 216958 584960 216960
rect 580625 216955 580691 216958
rect 583520 216868 584960 216958
rect 236269 212530 236335 212533
rect 236453 212530 236519 212533
rect 249241 212532 249307 212533
rect 249190 212530 249196 212532
rect 236269 212528 236519 212530
rect 236269 212472 236274 212528
rect 236330 212472 236458 212528
rect 236514 212472 236519 212528
rect 236269 212470 236519 212472
rect 249150 212470 249196 212530
rect 249260 212528 249307 212532
rect 249302 212472 249307 212528
rect 236269 212467 236335 212470
rect 236453 212467 236519 212470
rect 249190 212468 249196 212470
rect 249260 212468 249307 212472
rect 249241 212467 249307 212468
rect 389265 212530 389331 212533
rect 389449 212530 389515 212533
rect 389265 212528 389515 212530
rect 389265 212472 389270 212528
rect 389326 212472 389454 212528
rect 389510 212472 389515 212528
rect 389265 212470 389515 212472
rect 389265 212467 389331 212470
rect 389449 212467 389515 212470
rect 463785 212530 463851 212533
rect 463969 212530 464035 212533
rect 463785 212528 464035 212530
rect 463785 212472 463790 212528
rect 463846 212472 463974 212528
rect 464030 212472 464035 212528
rect 463785 212470 464035 212472
rect 463785 212467 463851 212470
rect 463969 212467 464035 212470
rect 470409 212530 470475 212533
rect 470593 212530 470659 212533
rect 470409 212528 470659 212530
rect 470409 212472 470414 212528
rect 470470 212472 470598 212528
rect 470654 212472 470659 212528
rect 470409 212470 470659 212472
rect 470409 212467 470475 212470
rect 470593 212467 470659 212470
rect 357433 211170 357499 211173
rect 357709 211170 357775 211173
rect 357433 211168 357775 211170
rect 357433 211112 357438 211168
rect 357494 211112 357714 211168
rect 357770 211112 357775 211168
rect 357433 211110 357775 211112
rect 357433 211107 357499 211110
rect 357709 211107 357775 211110
rect 358537 211170 358603 211173
rect 358721 211170 358787 211173
rect 358537 211168 358787 211170
rect 358537 211112 358542 211168
rect 358598 211112 358726 211168
rect 358782 211112 358787 211168
rect 358537 211110 358787 211112
rect 358537 211107 358603 211110
rect 358721 211107 358787 211110
rect -960 208178 480 208268
rect 3785 208178 3851 208181
rect -960 208176 3851 208178
rect -960 208120 3790 208176
rect 3846 208120 3851 208176
rect -960 208118 3851 208120
rect -960 208028 480 208118
rect 3785 208115 3851 208118
rect 249241 205458 249307 205461
rect 249558 205458 249564 205460
rect 249241 205456 249564 205458
rect 249241 205400 249246 205456
rect 249302 205400 249564 205456
rect 249241 205398 249564 205400
rect 249241 205395 249307 205398
rect 249558 205396 249564 205398
rect 249628 205396 249634 205460
rect 580533 205322 580599 205325
rect 583520 205322 584960 205412
rect 580533 205320 584960 205322
rect 580533 205264 580538 205320
rect 580594 205264 584960 205320
rect 580533 205262 584960 205264
rect 580533 205259 580599 205262
rect 583520 205172 584960 205262
rect 230749 202874 230815 202877
rect 231025 202874 231091 202877
rect 230749 202872 231091 202874
rect 230749 202816 230754 202872
rect 230810 202816 231030 202872
rect 231086 202816 231091 202872
rect 230749 202814 231091 202816
rect 230749 202811 230815 202814
rect 231025 202811 231091 202814
rect 232221 202874 232287 202877
rect 244273 202874 244339 202877
rect 244457 202874 244523 202877
rect 249609 202876 249675 202877
rect 232221 202872 232330 202874
rect 232221 202816 232226 202872
rect 232282 202816 232330 202872
rect 232221 202811 232330 202816
rect 244273 202872 244523 202874
rect 244273 202816 244278 202872
rect 244334 202816 244462 202872
rect 244518 202816 244523 202872
rect 244273 202814 244523 202816
rect 244273 202811 244339 202814
rect 244457 202811 244523 202814
rect 249558 202812 249564 202876
rect 249628 202874 249675 202876
rect 251449 202874 251515 202877
rect 251633 202874 251699 202877
rect 249628 202872 249720 202874
rect 249670 202816 249720 202872
rect 249628 202814 249720 202816
rect 251449 202872 251699 202874
rect 251449 202816 251454 202872
rect 251510 202816 251638 202872
rect 251694 202816 251699 202872
rect 251449 202814 251699 202816
rect 249628 202812 249675 202814
rect 249609 202811 249675 202812
rect 251449 202811 251515 202814
rect 251633 202811 251699 202814
rect 259637 202874 259703 202877
rect 259913 202874 259979 202877
rect 259637 202872 259979 202874
rect 259637 202816 259642 202872
rect 259698 202816 259918 202872
rect 259974 202816 259979 202872
rect 259637 202814 259979 202816
rect 259637 202811 259703 202814
rect 259913 202811 259979 202814
rect 262581 202874 262647 202877
rect 265157 202874 265223 202877
rect 265341 202874 265407 202877
rect 270677 202874 270743 202877
rect 272149 202876 272215 202877
rect 272149 202874 272196 202876
rect 262581 202872 262690 202874
rect 262581 202816 262586 202872
rect 262642 202816 262690 202872
rect 262581 202811 262690 202816
rect 265157 202872 265407 202874
rect 265157 202816 265162 202872
rect 265218 202816 265346 202872
rect 265402 202816 265407 202872
rect 265157 202814 265407 202816
rect 265157 202811 265223 202814
rect 265341 202811 265407 202814
rect 270542 202872 270743 202874
rect 270542 202816 270682 202872
rect 270738 202816 270743 202872
rect 270542 202814 270743 202816
rect 272104 202872 272196 202874
rect 272104 202816 272154 202872
rect 272104 202814 272196 202816
rect 232270 202741 232330 202811
rect 262630 202741 262690 202811
rect 232270 202736 232379 202741
rect 232270 202680 232318 202736
rect 232374 202680 232379 202736
rect 232270 202678 232379 202680
rect 262630 202736 262739 202741
rect 262630 202680 262678 202736
rect 262734 202680 262739 202736
rect 262630 202678 262739 202680
rect 270542 202738 270602 202814
rect 270677 202811 270743 202814
rect 272149 202812 272196 202814
rect 272260 202812 272266 202876
rect 285765 202874 285831 202877
rect 285949 202874 286015 202877
rect 285765 202872 286015 202874
rect 285765 202816 285770 202872
rect 285826 202816 285954 202872
rect 286010 202816 286015 202872
rect 285765 202814 286015 202816
rect 272149 202811 272215 202812
rect 285765 202811 285831 202814
rect 285949 202811 286015 202814
rect 325877 202874 325943 202877
rect 329925 202874 329991 202877
rect 330109 202874 330175 202877
rect 325877 202872 325986 202874
rect 325877 202816 325882 202872
rect 325938 202816 325986 202872
rect 325877 202811 325986 202816
rect 329925 202872 330175 202874
rect 329925 202816 329930 202872
rect 329986 202816 330114 202872
rect 330170 202816 330175 202872
rect 329925 202814 330175 202816
rect 329925 202811 329991 202814
rect 330109 202811 330175 202814
rect 331397 202874 331463 202877
rect 331581 202874 331647 202877
rect 331397 202872 331647 202874
rect 331397 202816 331402 202872
rect 331458 202816 331586 202872
rect 331642 202816 331647 202872
rect 331397 202814 331647 202816
rect 331397 202811 331463 202814
rect 331581 202811 331647 202814
rect 338665 202874 338731 202877
rect 338849 202874 338915 202877
rect 338665 202872 338915 202874
rect 338665 202816 338670 202872
rect 338726 202816 338854 202872
rect 338910 202816 338915 202872
rect 338665 202814 338915 202816
rect 338665 202811 338731 202814
rect 338849 202811 338915 202814
rect 372521 202874 372587 202877
rect 372705 202874 372771 202877
rect 372521 202872 372771 202874
rect 372521 202816 372526 202872
rect 372582 202816 372710 202872
rect 372766 202816 372771 202872
rect 372521 202814 372771 202816
rect 372521 202811 372587 202814
rect 372705 202811 372771 202814
rect 376937 202874 377003 202877
rect 377121 202874 377187 202877
rect 376937 202872 377187 202874
rect 376937 202816 376942 202872
rect 376998 202816 377126 202872
rect 377182 202816 377187 202872
rect 376937 202814 377187 202816
rect 376937 202811 377003 202814
rect 377121 202811 377187 202814
rect 325926 202741 325986 202811
rect 270677 202738 270743 202741
rect 270542 202736 270743 202738
rect 270542 202680 270682 202736
rect 270738 202680 270743 202736
rect 270542 202678 270743 202680
rect 325926 202736 326035 202741
rect 325926 202680 325974 202736
rect 326030 202680 326035 202736
rect 325926 202678 326035 202680
rect 232313 202675 232379 202678
rect 262673 202675 262739 202678
rect 270677 202675 270743 202678
rect 325969 202675 326035 202678
rect 290273 201650 290339 201653
rect 291837 201650 291903 201653
rect 290046 201648 290339 201650
rect 290046 201592 290278 201648
rect 290334 201592 290339 201648
rect 290046 201590 290339 201592
rect 284753 201514 284819 201517
rect 284937 201514 285003 201517
rect 284753 201512 285003 201514
rect 284753 201456 284758 201512
rect 284814 201456 284942 201512
rect 284998 201456 285003 201512
rect 284753 201454 285003 201456
rect 290046 201514 290106 201590
rect 290273 201587 290339 201590
rect 291518 201648 291903 201650
rect 291518 201592 291842 201648
rect 291898 201592 291903 201648
rect 291518 201590 291903 201592
rect 290181 201514 290247 201517
rect 290046 201512 290247 201514
rect 290046 201456 290186 201512
rect 290242 201456 290247 201512
rect 290046 201454 290247 201456
rect 291518 201514 291578 201590
rect 291837 201587 291903 201590
rect 291653 201514 291719 201517
rect 291518 201512 291719 201514
rect 291518 201456 291658 201512
rect 291714 201456 291719 201512
rect 291518 201454 291719 201456
rect 284753 201451 284819 201454
rect 284937 201451 285003 201454
rect 290181 201451 290247 201454
rect 291653 201451 291719 201454
rect 337101 201514 337167 201517
rect 337377 201514 337443 201517
rect 337101 201512 337443 201514
rect 337101 201456 337106 201512
rect 337162 201456 337382 201512
rect 337438 201456 337443 201512
rect 337101 201454 337443 201456
rect 337101 201451 337167 201454
rect 337377 201451 337443 201454
rect 299841 200290 299907 200293
rect 299798 200288 299907 200290
rect 299798 200232 299846 200288
rect 299902 200232 299907 200288
rect 299798 200227 299907 200232
rect 299798 200157 299858 200227
rect 299749 200152 299858 200157
rect 299749 200096 299754 200152
rect 299810 200096 299858 200152
rect 299749 200094 299858 200096
rect 306741 200154 306807 200157
rect 306925 200154 306991 200157
rect 306741 200152 306991 200154
rect 306741 200096 306746 200152
rect 306802 200096 306930 200152
rect 306986 200096 306991 200152
rect 306741 200094 306991 200096
rect 299749 200091 299815 200094
rect 306741 200091 306807 200094
rect 306925 200091 306991 200094
rect 249374 196556 249380 196620
rect 249444 196618 249450 196620
rect 249609 196618 249675 196621
rect 249444 196616 249675 196618
rect 249444 196560 249614 196616
rect 249670 196560 249675 196616
rect 249444 196558 249675 196560
rect 249444 196556 249450 196558
rect 249609 196555 249675 196558
rect -960 193898 480 193988
rect 3693 193898 3759 193901
rect -960 193896 3759 193898
rect -960 193840 3698 193896
rect 3754 193840 3759 193896
rect -960 193838 3759 193840
rect -960 193748 480 193838
rect 3693 193835 3759 193838
rect 583520 193476 584960 193716
rect 236269 193218 236335 193221
rect 236453 193218 236519 193221
rect 236269 193216 236519 193218
rect 236269 193160 236274 193216
rect 236330 193160 236458 193216
rect 236514 193160 236519 193216
rect 236269 193158 236519 193160
rect 236269 193155 236335 193158
rect 236453 193155 236519 193158
rect 310789 193218 310855 193221
rect 311065 193218 311131 193221
rect 310789 193216 311131 193218
rect 310789 193160 310794 193216
rect 310850 193160 311070 193216
rect 311126 193160 311131 193216
rect 310789 193158 311131 193160
rect 310789 193155 310855 193158
rect 311065 193155 311131 193158
rect 323301 193218 323367 193221
rect 323485 193218 323551 193221
rect 323301 193216 323551 193218
rect 323301 193160 323306 193216
rect 323362 193160 323490 193216
rect 323546 193160 323551 193216
rect 323301 193158 323551 193160
rect 323301 193155 323367 193158
rect 323485 193155 323551 193158
rect 357709 193218 357775 193221
rect 357893 193218 357959 193221
rect 357709 193216 357959 193218
rect 357709 193160 357714 193216
rect 357770 193160 357898 193216
rect 357954 193160 357959 193216
rect 357709 193158 357959 193160
rect 357709 193155 357775 193158
rect 357893 193155 357959 193158
rect 389265 193218 389331 193221
rect 389449 193218 389515 193221
rect 389265 193216 389515 193218
rect 389265 193160 389270 193216
rect 389326 193160 389454 193216
rect 389510 193160 389515 193216
rect 389265 193158 389515 193160
rect 389265 193155 389331 193158
rect 389449 193155 389515 193158
rect 463785 193218 463851 193221
rect 463969 193218 464035 193221
rect 463785 193216 464035 193218
rect 463785 193160 463790 193216
rect 463846 193160 463974 193216
rect 464030 193160 464035 193216
rect 463785 193158 464035 193160
rect 463785 193155 463851 193158
rect 463969 193155 464035 193158
rect 470409 193218 470475 193221
rect 470593 193218 470659 193221
rect 470409 193216 470659 193218
rect 470409 193160 470414 193216
rect 470470 193160 470598 193216
rect 470654 193160 470659 193216
rect 470409 193158 470659 193160
rect 470409 193155 470475 193158
rect 470593 193155 470659 193158
rect 249374 191824 249380 191826
rect 249198 191764 249380 191824
rect 249198 191589 249258 191764
rect 249374 191762 249380 191764
rect 249444 191762 249450 191826
rect 249198 191584 249307 191589
rect 249198 191528 249246 191584
rect 249302 191528 249307 191584
rect 249198 191526 249307 191528
rect 249241 191523 249307 191526
rect 272241 190500 272307 190501
rect 272190 190498 272196 190500
rect 272150 190438 272196 190498
rect 272260 190496 272307 190500
rect 272302 190440 272307 190496
rect 272190 190436 272196 190438
rect 272260 190436 272307 190440
rect 272241 190435 272307 190436
rect 289905 190498 289971 190501
rect 290089 190498 290155 190501
rect 289905 190496 290155 190498
rect 289905 190440 289910 190496
rect 289966 190440 290094 190496
rect 290150 190440 290155 190496
rect 289905 190438 290155 190440
rect 289905 190435 289971 190438
rect 290089 190435 290155 190438
rect 291377 190498 291443 190501
rect 291561 190498 291627 190501
rect 291377 190496 291627 190498
rect 291377 190440 291382 190496
rect 291438 190440 291566 190496
rect 291622 190440 291627 190496
rect 291377 190438 291627 190440
rect 291377 190435 291443 190438
rect 291561 190435 291627 190438
rect 230749 183562 230815 183565
rect 231025 183562 231091 183565
rect 230749 183560 231091 183562
rect 230749 183504 230754 183560
rect 230810 183504 231030 183560
rect 231086 183504 231091 183560
rect 230749 183502 231091 183504
rect 230749 183499 230815 183502
rect 231025 183499 231091 183502
rect 232221 183562 232287 183565
rect 236269 183562 236335 183565
rect 236453 183562 236519 183565
rect 232221 183560 232330 183562
rect 232221 183504 232226 183560
rect 232282 183504 232330 183560
rect 232221 183499 232330 183504
rect 236269 183560 236519 183562
rect 236269 183504 236274 183560
rect 236330 183504 236458 183560
rect 236514 183504 236519 183560
rect 236269 183502 236519 183504
rect 236269 183499 236335 183502
rect 236453 183499 236519 183502
rect 251449 183562 251515 183565
rect 251633 183562 251699 183565
rect 251449 183560 251699 183562
rect 251449 183504 251454 183560
rect 251510 183504 251638 183560
rect 251694 183504 251699 183560
rect 251449 183502 251699 183504
rect 251449 183499 251515 183502
rect 251633 183499 251699 183502
rect 262581 183562 262647 183565
rect 262765 183562 262831 183565
rect 270677 183562 270743 183565
rect 262581 183560 262831 183562
rect 262581 183504 262586 183560
rect 262642 183504 262770 183560
rect 262826 183504 262831 183560
rect 262581 183502 262831 183504
rect 262581 183499 262647 183502
rect 262765 183499 262831 183502
rect 270542 183560 270743 183562
rect 270542 183504 270682 183560
rect 270738 183504 270743 183560
rect 270542 183502 270743 183504
rect 232270 183429 232330 183499
rect 232270 183424 232379 183429
rect 232270 183368 232318 183424
rect 232374 183368 232379 183424
rect 232270 183366 232379 183368
rect 270542 183426 270602 183502
rect 270677 183499 270743 183502
rect 285949 183562 286015 183565
rect 325877 183562 325943 183565
rect 326061 183562 326127 183565
rect 285949 183560 286058 183562
rect 285949 183504 285954 183560
rect 286010 183504 286058 183560
rect 285949 183499 286058 183504
rect 325877 183560 326127 183562
rect 325877 183504 325882 183560
rect 325938 183504 326066 183560
rect 326122 183504 326127 183560
rect 325877 183502 326127 183504
rect 325877 183499 325943 183502
rect 326061 183499 326127 183502
rect 331397 183562 331463 183565
rect 331581 183562 331647 183565
rect 331397 183560 331647 183562
rect 331397 183504 331402 183560
rect 331458 183504 331586 183560
rect 331642 183504 331647 183560
rect 331397 183502 331647 183504
rect 331397 183499 331463 183502
rect 331581 183499 331647 183502
rect 366817 183562 366883 183565
rect 367001 183562 367067 183565
rect 366817 183560 367067 183562
rect 366817 183504 366822 183560
rect 366878 183504 367006 183560
rect 367062 183504 367067 183560
rect 366817 183502 367067 183504
rect 366817 183499 366883 183502
rect 367001 183499 367067 183502
rect 372521 183562 372587 183565
rect 372705 183562 372771 183565
rect 372521 183560 372771 183562
rect 372521 183504 372526 183560
rect 372582 183504 372710 183560
rect 372766 183504 372771 183560
rect 372521 183502 372771 183504
rect 372521 183499 372587 183502
rect 372705 183499 372771 183502
rect 376937 183562 377003 183565
rect 377121 183562 377187 183565
rect 376937 183560 377187 183562
rect 376937 183504 376942 183560
rect 376998 183504 377126 183560
rect 377182 183504 377187 183560
rect 376937 183502 377187 183504
rect 376937 183499 377003 183502
rect 377121 183499 377187 183502
rect 285998 183429 286058 183499
rect 270861 183426 270927 183429
rect 270542 183424 270927 183426
rect 270542 183368 270866 183424
rect 270922 183368 270927 183424
rect 270542 183366 270927 183368
rect 232313 183363 232379 183366
rect 270861 183363 270927 183366
rect 285949 183424 286058 183429
rect 285949 183368 285954 183424
rect 286010 183368 286058 183424
rect 285949 183366 286058 183368
rect 285949 183363 286015 183366
rect 249241 182204 249307 182205
rect 249190 182202 249196 182204
rect 249150 182142 249196 182202
rect 249260 182200 249307 182204
rect 249302 182144 249307 182200
rect 249190 182140 249196 182142
rect 249260 182140 249307 182144
rect 249241 182139 249307 182140
rect 324497 182202 324563 182205
rect 324865 182202 324931 182205
rect 324497 182200 324931 182202
rect 324497 182144 324502 182200
rect 324558 182144 324870 182200
rect 324926 182144 324931 182200
rect 324497 182142 324931 182144
rect 324497 182139 324563 182142
rect 324865 182139 324931 182142
rect 330109 182202 330175 182205
rect 330293 182202 330359 182205
rect 330109 182200 330359 182202
rect 330109 182144 330114 182200
rect 330170 182144 330298 182200
rect 330354 182144 330359 182200
rect 330109 182142 330359 182144
rect 330109 182139 330175 182142
rect 330293 182139 330359 182142
rect 358537 182202 358603 182205
rect 358721 182202 358787 182205
rect 358537 182200 358787 182202
rect 358537 182144 358542 182200
rect 358598 182144 358726 182200
rect 358782 182144 358787 182200
rect 358537 182142 358787 182144
rect 358537 182139 358603 182142
rect 358721 182139 358787 182142
rect 580441 181930 580507 181933
rect 583520 181930 584960 182020
rect 580441 181928 584960 181930
rect 580441 181872 580446 181928
rect 580502 181872 584960 181928
rect 580441 181870 584960 181872
rect 580441 181867 580507 181870
rect 583520 181780 584960 181870
rect 264973 180842 265039 180845
rect 265157 180842 265223 180845
rect 264973 180840 265223 180842
rect 264973 180784 264978 180840
rect 265034 180784 265162 180840
rect 265218 180784 265223 180840
rect 264973 180782 265223 180784
rect 264973 180779 265039 180782
rect 265157 180779 265223 180782
rect 249190 180644 249196 180708
rect 249260 180644 249266 180708
rect 249198 180570 249258 180644
rect 249425 180570 249491 180573
rect 249198 180568 249491 180570
rect 249198 180512 249430 180568
rect 249486 180512 249491 180568
rect 249198 180510 249491 180512
rect 249425 180507 249491 180510
rect -960 179482 480 179572
rect 3601 179482 3667 179485
rect -960 179480 3667 179482
rect -960 179424 3606 179480
rect 3662 179424 3667 179480
rect -960 179422 3667 179424
rect -960 179332 480 179422
rect 3601 179419 3667 179422
rect 341241 179482 341307 179485
rect 341425 179482 341491 179485
rect 341241 179480 341491 179482
rect 341241 179424 341246 179480
rect 341302 179424 341430 179480
rect 341486 179424 341491 179480
rect 341241 179422 341491 179424
rect 341241 179419 341307 179422
rect 341425 179419 341491 179422
rect 236361 173906 236427 173909
rect 236545 173906 236611 173909
rect 236361 173904 236611 173906
rect 236361 173848 236366 173904
rect 236422 173848 236550 173904
rect 236606 173848 236611 173904
rect 236361 173846 236611 173848
rect 236361 173843 236427 173846
rect 236545 173843 236611 173846
rect 249425 173906 249491 173909
rect 367001 173908 367067 173909
rect 249742 173906 249748 173908
rect 249425 173904 249748 173906
rect 249425 173848 249430 173904
rect 249486 173848 249748 173904
rect 249425 173846 249748 173848
rect 249425 173843 249491 173846
rect 249742 173844 249748 173846
rect 249812 173844 249818 173908
rect 366950 173906 366956 173908
rect 366910 173846 366956 173906
rect 367020 173904 367067 173908
rect 367062 173848 367067 173904
rect 366950 173844 366956 173846
rect 367020 173844 367067 173848
rect 367001 173843 367067 173844
rect 470409 173906 470475 173909
rect 470593 173906 470659 173909
rect 470409 173904 470659 173906
rect 470409 173848 470414 173904
rect 470470 173848 470598 173904
rect 470654 173848 470659 173904
rect 470409 173846 470659 173848
rect 470409 173843 470475 173846
rect 470593 173843 470659 173846
rect 289997 172682 290063 172685
rect 291469 172682 291535 172685
rect 289862 172680 290063 172682
rect 289862 172624 290002 172680
rect 290058 172624 290063 172680
rect 289862 172622 290063 172624
rect 289862 172546 289922 172622
rect 289997 172619 290063 172622
rect 291334 172680 291535 172682
rect 291334 172624 291474 172680
rect 291530 172624 291535 172680
rect 291334 172622 291535 172624
rect 289997 172546 290063 172549
rect 289862 172544 290063 172546
rect 289862 172488 290002 172544
rect 290058 172488 290063 172544
rect 289862 172486 290063 172488
rect 291334 172546 291394 172622
rect 291469 172619 291535 172622
rect 291469 172546 291535 172549
rect 291334 172544 291535 172546
rect 291334 172488 291474 172544
rect 291530 172488 291535 172544
rect 291334 172486 291535 172488
rect 289997 172483 290063 172486
rect 291469 172483 291535 172486
rect 325969 172546 326035 172549
rect 326245 172546 326311 172549
rect 325969 172544 326311 172546
rect 325969 172488 325974 172544
rect 326030 172488 326250 172544
rect 326306 172488 326311 172544
rect 325969 172486 326311 172488
rect 325969 172483 326035 172486
rect 326245 172483 326311 172486
rect 580349 170098 580415 170101
rect 583520 170098 584960 170188
rect 580349 170096 584960 170098
rect 580349 170040 580354 170096
rect 580410 170040 584960 170096
rect 580349 170038 584960 170040
rect 580349 170035 580415 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 2773 165066 2839 165069
rect -960 165064 2839 165066
rect -960 165008 2778 165064
rect 2834 165008 2839 165064
rect -960 165006 2839 165008
rect -960 164916 480 165006
rect 2773 165003 2839 165006
rect 357617 164386 357683 164389
rect 357390 164384 357683 164386
rect 357390 164328 357622 164384
rect 357678 164328 357683 164384
rect 357390 164326 357683 164328
rect 236269 164250 236335 164253
rect 236545 164250 236611 164253
rect 236269 164248 236611 164250
rect 236269 164192 236274 164248
rect 236330 164192 236550 164248
rect 236606 164192 236611 164248
rect 236269 164190 236611 164192
rect 236269 164187 236335 164190
rect 236545 164187 236611 164190
rect 249374 164188 249380 164252
rect 249444 164250 249450 164252
rect 249742 164250 249748 164252
rect 249444 164190 249748 164250
rect 249444 164188 249450 164190
rect 249742 164188 249748 164190
rect 249812 164188 249818 164252
rect 259637 164250 259703 164253
rect 259913 164250 259979 164253
rect 259637 164248 259979 164250
rect 259637 164192 259642 164248
rect 259698 164192 259918 164248
rect 259974 164192 259979 164248
rect 259637 164190 259979 164192
rect 357390 164250 357450 164326
rect 357617 164323 357683 164326
rect 357525 164250 357591 164253
rect 367001 164252 367067 164253
rect 366950 164250 366956 164252
rect 357390 164248 357591 164250
rect 357390 164192 357530 164248
rect 357586 164192 357591 164248
rect 357390 164190 357591 164192
rect 366910 164190 366956 164250
rect 367020 164248 367067 164252
rect 367062 164192 367067 164248
rect 259637 164187 259703 164190
rect 259913 164187 259979 164190
rect 357525 164187 357591 164190
rect 366950 164188 366956 164190
rect 367020 164188 367067 164192
rect 367001 164187 367067 164188
rect 470409 164250 470475 164253
rect 470593 164250 470659 164253
rect 470409 164248 470659 164250
rect 470409 164192 470414 164248
rect 470470 164192 470598 164248
rect 470654 164192 470659 164248
rect 470409 164190 470659 164192
rect 470409 164187 470475 164190
rect 470593 164187 470659 164190
rect 270493 162890 270559 162893
rect 270677 162890 270743 162893
rect 270493 162888 270743 162890
rect 270493 162832 270498 162888
rect 270554 162832 270682 162888
rect 270738 162832 270743 162888
rect 270493 162830 270743 162832
rect 270493 162827 270559 162830
rect 270677 162827 270743 162830
rect 272241 162890 272307 162893
rect 272425 162890 272491 162893
rect 272241 162888 272491 162890
rect 272241 162832 272246 162888
rect 272302 162832 272430 162888
rect 272486 162832 272491 162888
rect 272241 162830 272491 162832
rect 272241 162827 272307 162830
rect 272425 162827 272491 162830
rect 330109 162890 330175 162893
rect 330293 162890 330359 162893
rect 330109 162888 330359 162890
rect 330109 162832 330114 162888
rect 330170 162832 330298 162888
rect 330354 162832 330359 162888
rect 330109 162830 330359 162832
rect 330109 162827 330175 162830
rect 330293 162827 330359 162830
rect 306833 161530 306899 161533
rect 307017 161530 307083 161533
rect 306833 161528 307083 161530
rect 306833 161472 306838 161528
rect 306894 161472 307022 161528
rect 307078 161472 307083 161528
rect 306833 161470 307083 161472
rect 306833 161467 306899 161470
rect 307017 161467 307083 161470
rect 583520 158402 584960 158492
rect 583342 158342 584960 158402
rect 405406 157858 405412 157860
rect 398606 157798 405412 157858
rect 278681 157722 278747 157725
rect 269254 157720 278747 157722
rect 269254 157664 278686 157720
rect 278742 157664 278747 157720
rect 269254 157662 278747 157664
rect 269254 157586 269314 157662
rect 278681 157659 278747 157662
rect 324262 157660 324268 157724
rect 324332 157722 324338 157724
rect 324332 157662 340890 157722
rect 324332 157660 324338 157662
rect 253614 157526 254410 157586
rect 249374 157388 249380 157452
rect 249444 157450 249450 157452
rect 253614 157450 253674 157526
rect 249444 157390 253674 157450
rect 254350 157450 254410 157526
rect 256190 157526 264346 157586
rect 256190 157450 256250 157526
rect 254350 157390 256250 157450
rect 264286 157450 264346 157526
rect 269070 157526 269314 157586
rect 278681 157586 278747 157589
rect 278681 157584 278882 157586
rect 278681 157528 278686 157584
rect 278742 157528 278882 157584
rect 278681 157526 278882 157528
rect 269070 157450 269130 157526
rect 278681 157523 278747 157526
rect 264286 157390 269130 157450
rect 278822 157450 278882 157526
rect 282637 157450 282703 157453
rect 278822 157448 282703 157450
rect 278822 157392 282642 157448
rect 282698 157392 282703 157448
rect 278822 157390 282703 157392
rect 249444 157388 249450 157390
rect 282637 157387 282703 157390
rect 288893 157450 288959 157453
rect 306281 157450 306347 157453
rect 288893 157448 306347 157450
rect 288893 157392 288898 157448
rect 288954 157392 306286 157448
rect 306342 157392 306347 157448
rect 288893 157390 306347 157392
rect 288893 157387 288959 157390
rect 306281 157387 306347 157390
rect 314561 157450 314627 157453
rect 324262 157450 324268 157452
rect 314561 157448 324268 157450
rect 314561 157392 314566 157448
rect 314622 157392 324268 157448
rect 314561 157390 324268 157392
rect 314561 157387 314627 157390
rect 324262 157388 324268 157390
rect 324332 157388 324338 157452
rect 340830 157450 340890 157662
rect 360101 157586 360167 157589
rect 350582 157584 360167 157586
rect 350582 157528 360106 157584
rect 360162 157528 360167 157584
rect 350582 157526 360167 157528
rect 350582 157450 350642 157526
rect 360101 157523 360167 157526
rect 360285 157586 360351 157589
rect 398606 157586 398666 157798
rect 405406 157796 405412 157798
rect 405476 157796 405482 157860
rect 470550 157662 480178 157722
rect 417877 157586 417943 157589
rect 360285 157584 369778 157586
rect 360285 157528 360290 157584
rect 360346 157528 369778 157584
rect 360285 157526 369778 157528
rect 360285 157523 360351 157526
rect 340830 157390 350642 157450
rect 369718 157450 369778 157526
rect 389222 157526 398666 157586
rect 408542 157584 417943 157586
rect 408542 157528 417882 157584
rect 417938 157528 417943 157584
rect 408542 157526 417943 157528
rect 389222 157450 389282 157526
rect 369718 157390 389282 157450
rect 405590 157388 405596 157452
rect 405660 157450 405666 157452
rect 408542 157450 408602 157526
rect 417877 157523 417943 157526
rect 418153 157586 418219 157589
rect 437197 157586 437263 157589
rect 418153 157584 424978 157586
rect 418153 157528 418158 157584
rect 418214 157528 424978 157584
rect 418153 157526 424978 157528
rect 418153 157523 418219 157526
rect 405660 157390 408602 157450
rect 424918 157450 424978 157526
rect 427862 157584 437263 157586
rect 427862 157528 437202 157584
rect 437258 157528 437263 157584
rect 427862 157526 437263 157528
rect 427862 157450 427922 157526
rect 437197 157523 437263 157526
rect 437473 157586 437539 157589
rect 456517 157586 456583 157589
rect 437473 157584 444298 157586
rect 437473 157528 437478 157584
rect 437534 157528 444298 157584
rect 437473 157526 444298 157528
rect 437473 157523 437539 157526
rect 424918 157390 427922 157450
rect 444238 157450 444298 157526
rect 447182 157584 456583 157586
rect 447182 157528 456522 157584
rect 456578 157528 456583 157584
rect 447182 157526 456583 157528
rect 447182 157450 447242 157526
rect 456517 157523 456583 157526
rect 456885 157586 456951 157589
rect 456885 157584 466378 157586
rect 456885 157528 456890 157584
rect 456946 157528 466378 157584
rect 456885 157526 466378 157528
rect 456885 157523 456951 157526
rect 444238 157390 447242 157450
rect 466318 157450 466378 157526
rect 470550 157450 470610 157662
rect 466318 157390 470610 157450
rect 480118 157450 480178 157662
rect 480302 157662 489930 157722
rect 480302 157450 480362 157662
rect 489870 157586 489930 157662
rect 499622 157662 509250 157722
rect 489870 157526 499498 157586
rect 480118 157390 480362 157450
rect 499438 157450 499498 157526
rect 499622 157450 499682 157662
rect 509190 157586 509250 157662
rect 518942 157662 528570 157722
rect 509190 157526 518818 157586
rect 499438 157390 499682 157450
rect 518758 157450 518818 157526
rect 518942 157450 519002 157662
rect 528510 157586 528570 157662
rect 538262 157662 547890 157722
rect 528510 157526 538138 157586
rect 518758 157390 519002 157450
rect 538078 157450 538138 157526
rect 538262 157450 538322 157662
rect 547830 157586 547890 157662
rect 557582 157662 567210 157722
rect 547830 157526 557458 157586
rect 538078 157390 538322 157450
rect 557398 157450 557458 157526
rect 557582 157450 557642 157662
rect 567150 157586 567210 157662
rect 583342 157586 583402 158342
rect 583520 158252 584960 158342
rect 567150 157526 576778 157586
rect 557398 157390 557642 157450
rect 576718 157450 576778 157526
rect 576902 157526 583402 157586
rect 576902 157450 576962 157526
rect 576718 157390 576962 157450
rect 405660 157388 405666 157390
rect 250345 154730 250411 154733
rect 249934 154728 250411 154730
rect 249934 154672 250350 154728
rect 250406 154672 250411 154728
rect 249934 154670 250411 154672
rect 244273 154594 244339 154597
rect 244457 154594 244523 154597
rect 244273 154592 244523 154594
rect 244273 154536 244278 154592
rect 244334 154536 244462 154592
rect 244518 154536 244523 154592
rect 244273 154534 244523 154536
rect 249934 154594 249994 154670
rect 250345 154667 250411 154670
rect 338849 154730 338915 154733
rect 338849 154728 339050 154730
rect 338849 154672 338854 154728
rect 338910 154672 339050 154728
rect 338849 154670 339050 154672
rect 338849 154667 338915 154670
rect 250069 154594 250135 154597
rect 249934 154592 250135 154594
rect 249934 154536 250074 154592
rect 250130 154536 250135 154592
rect 249934 154534 250135 154536
rect 244273 154531 244339 154534
rect 244457 154531 244523 154534
rect 250069 154531 250135 154534
rect 251449 154594 251515 154597
rect 251633 154594 251699 154597
rect 251449 154592 251699 154594
rect 251449 154536 251454 154592
rect 251510 154536 251638 154592
rect 251694 154536 251699 154592
rect 251449 154534 251699 154536
rect 251449 154531 251515 154534
rect 251633 154531 251699 154534
rect 338849 154594 338915 154597
rect 338990 154594 339050 154670
rect 338849 154592 339050 154594
rect 338849 154536 338854 154592
rect 338910 154536 339050 154592
rect 338849 154534 339050 154536
rect 376937 154594 377003 154597
rect 377121 154594 377187 154597
rect 376937 154592 377187 154594
rect 376937 154536 376942 154592
rect 376998 154536 377126 154592
rect 377182 154536 377187 154592
rect 376937 154534 377187 154536
rect 338849 154531 338915 154534
rect 376937 154531 377003 154534
rect 377121 154531 377187 154534
rect 463877 154594 463943 154597
rect 464061 154594 464127 154597
rect 463877 154592 464127 154594
rect 463877 154536 463882 154592
rect 463938 154536 464066 154592
rect 464122 154536 464127 154592
rect 463877 154534 464127 154536
rect 463877 154531 463943 154534
rect 464061 154531 464127 154534
rect 310881 153370 310947 153373
rect 310838 153368 310947 153370
rect 310838 153312 310886 153368
rect 310942 153312 310947 153368
rect 310838 153307 310947 153312
rect 310838 153237 310898 153307
rect 285765 153234 285831 153237
rect 285949 153234 286015 153237
rect 285765 153232 286015 153234
rect 285765 153176 285770 153232
rect 285826 153176 285954 153232
rect 286010 153176 286015 153232
rect 285765 153174 286015 153176
rect 285765 153171 285831 153174
rect 285949 153171 286015 153174
rect 310789 153232 310898 153237
rect 310789 153176 310794 153232
rect 310850 153176 310898 153232
rect 310789 153174 310898 153176
rect 325969 153234 326035 153237
rect 326153 153234 326219 153237
rect 325969 153232 326219 153234
rect 325969 153176 325974 153232
rect 326030 153176 326158 153232
rect 326214 153176 326219 153232
rect 325969 153174 326219 153176
rect 310789 153171 310855 153174
rect 325969 153171 326035 153174
rect 326153 153171 326219 153174
rect 329925 153234 329991 153237
rect 330201 153234 330267 153237
rect 329925 153232 330267 153234
rect 329925 153176 329930 153232
rect 329986 153176 330206 153232
rect 330262 153176 330267 153232
rect 329925 153174 330267 153176
rect 329925 153171 329991 153174
rect 330201 153171 330267 153174
rect 296897 151738 296963 151741
rect 297173 151738 297239 151741
rect 296897 151736 297239 151738
rect 296897 151680 296902 151736
rect 296958 151680 297178 151736
rect 297234 151680 297239 151736
rect 296897 151678 297239 151680
rect 296897 151675 296963 151678
rect 297173 151675 297239 151678
rect -960 150786 480 150876
rect 3325 150786 3391 150789
rect -960 150784 3391 150786
rect -960 150728 3330 150784
rect 3386 150728 3391 150784
rect -960 150726 3391 150728
rect -960 150636 480 150726
rect 3325 150723 3391 150726
rect 583520 146556 584960 146796
rect 325969 145074 326035 145077
rect 325926 145072 326035 145074
rect 325926 145016 325974 145072
rect 326030 145016 326035 145072
rect 325926 145011 326035 145016
rect 325926 144941 325986 145011
rect 247125 144938 247191 144941
rect 247309 144938 247375 144941
rect 247125 144936 247375 144938
rect 247125 144880 247130 144936
rect 247186 144880 247314 144936
rect 247370 144880 247375 144936
rect 247125 144878 247375 144880
rect 247125 144875 247191 144878
rect 247309 144875 247375 144878
rect 325877 144936 325986 144941
rect 325877 144880 325882 144936
rect 325938 144880 325986 144936
rect 325877 144878 325986 144880
rect 327165 144938 327231 144941
rect 327349 144938 327415 144941
rect 327165 144936 327415 144938
rect 327165 144880 327170 144936
rect 327226 144880 327354 144936
rect 327410 144880 327415 144936
rect 327165 144878 327415 144880
rect 325877 144875 325943 144878
rect 327165 144875 327231 144878
rect 327349 144875 327415 144878
rect 389357 144938 389423 144941
rect 389633 144938 389699 144941
rect 389357 144936 389699 144938
rect 389357 144880 389362 144936
rect 389418 144880 389638 144936
rect 389694 144880 389699 144936
rect 389357 144878 389699 144880
rect 389357 144875 389423 144878
rect 389633 144875 389699 144878
rect 470409 144938 470475 144941
rect 470593 144938 470659 144941
rect 470409 144936 470659 144938
rect 470409 144880 470414 144936
rect 470470 144880 470598 144936
rect 470654 144880 470659 144936
rect 470409 144878 470659 144880
rect 470409 144875 470475 144878
rect 470593 144875 470659 144878
rect 302417 143578 302483 143581
rect 302601 143578 302667 143581
rect 302417 143576 302667 143578
rect 302417 143520 302422 143576
rect 302478 143520 302606 143576
rect 302662 143520 302667 143576
rect 302417 143518 302667 143520
rect 302417 143515 302483 143518
rect 302601 143515 302667 143518
rect 297173 142354 297239 142357
rect 296670 142352 297239 142354
rect 296670 142296 297178 142352
rect 297234 142296 297239 142352
rect 296670 142294 297239 142296
rect 296670 142218 296730 142294
rect 297173 142291 297239 142294
rect 296805 142218 296871 142221
rect 296670 142216 296871 142218
rect 296670 142160 296810 142216
rect 296866 142160 296871 142216
rect 296670 142158 296871 142160
rect 296805 142155 296871 142158
rect -960 136370 480 136460
rect 2773 136370 2839 136373
rect -960 136368 2839 136370
rect -960 136312 2778 136368
rect 2834 136312 2839 136368
rect -960 136310 2839 136312
rect -960 136220 480 136310
rect 2773 136307 2839 136310
rect 284753 135554 284819 135557
rect 284526 135552 284819 135554
rect 284526 135496 284758 135552
rect 284814 135496 284819 135552
rect 284526 135494 284819 135496
rect 234889 135282 234955 135285
rect 235165 135282 235231 135285
rect 234889 135280 235231 135282
rect 234889 135224 234894 135280
rect 234950 135224 235170 135280
rect 235226 135224 235231 135280
rect 234889 135222 235231 135224
rect 234889 135219 234955 135222
rect 235165 135219 235231 135222
rect 235993 135282 236059 135285
rect 236269 135282 236335 135285
rect 235993 135280 236335 135282
rect 235993 135224 235998 135280
rect 236054 135224 236274 135280
rect 236330 135224 236335 135280
rect 235993 135222 236335 135224
rect 235993 135219 236059 135222
rect 236269 135219 236335 135222
rect 244273 135282 244339 135285
rect 244457 135282 244523 135285
rect 244273 135280 244523 135282
rect 244273 135224 244278 135280
rect 244334 135224 244462 135280
rect 244518 135224 244523 135280
rect 244273 135222 244523 135224
rect 284526 135282 284586 135494
rect 284753 135491 284819 135494
rect 284661 135282 284727 135285
rect 284526 135280 284727 135282
rect 284526 135224 284666 135280
rect 284722 135224 284727 135280
rect 284526 135222 284727 135224
rect 244273 135219 244339 135222
rect 244457 135219 244523 135222
rect 284661 135219 284727 135222
rect 337101 135282 337167 135285
rect 337285 135282 337351 135285
rect 337101 135280 337351 135282
rect 337101 135224 337106 135280
rect 337162 135224 337290 135280
rect 337346 135224 337351 135280
rect 337101 135222 337351 135224
rect 337101 135219 337167 135222
rect 337285 135219 337351 135222
rect 376937 135282 377003 135285
rect 377121 135282 377187 135285
rect 376937 135280 377187 135282
rect 376937 135224 376942 135280
rect 376998 135224 377126 135280
rect 377182 135224 377187 135280
rect 376937 135222 377187 135224
rect 376937 135219 377003 135222
rect 377121 135219 377187 135222
rect 580257 134874 580323 134877
rect 583520 134874 584960 134964
rect 580257 134872 584960 134874
rect 580257 134816 580262 134872
rect 580318 134816 584960 134872
rect 580257 134814 584960 134816
rect 580257 134811 580323 134814
rect 583520 134724 584960 134814
rect 357249 133922 357315 133925
rect 357433 133922 357499 133925
rect 357249 133920 357499 133922
rect 357249 133864 357254 133920
rect 357310 133864 357438 133920
rect 357494 133864 357499 133920
rect 357249 133862 357499 133864
rect 357249 133859 357315 133862
rect 357433 133859 357499 133862
rect 341057 132562 341123 132565
rect 341241 132562 341307 132565
rect 341057 132560 341307 132562
rect 341057 132504 341062 132560
rect 341118 132504 341246 132560
rect 341302 132504 341307 132560
rect 341057 132502 341307 132504
rect 341057 132499 341123 132502
rect 341241 132499 341307 132502
rect 265157 125626 265223 125629
rect 265341 125626 265407 125629
rect 265157 125624 265407 125626
rect 265157 125568 265162 125624
rect 265218 125568 265346 125624
rect 265402 125568 265407 125624
rect 265157 125566 265407 125568
rect 265157 125563 265223 125566
rect 265341 125563 265407 125566
rect 270493 125626 270559 125629
rect 270677 125626 270743 125629
rect 270493 125624 270743 125626
rect 270493 125568 270498 125624
rect 270554 125568 270682 125624
rect 270738 125568 270743 125624
rect 270493 125566 270743 125568
rect 270493 125563 270559 125566
rect 270677 125563 270743 125566
rect 272149 125626 272215 125629
rect 272333 125626 272399 125629
rect 272149 125624 272399 125626
rect 272149 125568 272154 125624
rect 272210 125568 272338 125624
rect 272394 125568 272399 125624
rect 272149 125566 272399 125568
rect 272149 125563 272215 125566
rect 272333 125563 272399 125566
rect 324589 125626 324655 125629
rect 324773 125626 324839 125629
rect 324589 125624 324839 125626
rect 324589 125568 324594 125624
rect 324650 125568 324778 125624
rect 324834 125568 324839 125624
rect 324589 125566 324839 125568
rect 324589 125563 324655 125566
rect 324773 125563 324839 125566
rect 463877 125626 463943 125629
rect 464061 125626 464127 125629
rect 463877 125624 464127 125626
rect 463877 125568 463882 125624
rect 463938 125568 464066 125624
rect 464122 125568 464127 125624
rect 463877 125566 464127 125568
rect 463877 125563 463943 125566
rect 464061 125563 464127 125566
rect 470409 125626 470475 125629
rect 470593 125626 470659 125629
rect 470409 125624 470659 125626
rect 470409 125568 470414 125624
rect 470470 125568 470598 125624
rect 470654 125568 470659 125624
rect 470409 125566 470659 125568
rect 470409 125563 470475 125566
rect 470593 125563 470659 125566
rect 250161 124130 250227 124133
rect 250345 124130 250411 124133
rect 250161 124128 250411 124130
rect 250161 124072 250166 124128
rect 250222 124072 250350 124128
rect 250406 124072 250411 124128
rect 250161 124070 250411 124072
rect 250161 124067 250227 124070
rect 250345 124067 250411 124070
rect 467046 123116 467052 123180
rect 467116 123178 467122 123180
rect 583520 123178 584960 123268
rect 467116 123118 470610 123178
rect 467116 123116 467122 123118
rect 470550 123042 470610 123118
rect 480302 123118 489930 123178
rect 470550 122982 480178 123042
rect 480118 122906 480178 122982
rect 480302 122906 480362 123118
rect 489870 123042 489930 123118
rect 499622 123118 509250 123178
rect 489870 122982 499498 123042
rect 480118 122846 480362 122906
rect 499438 122906 499498 122982
rect 499622 122906 499682 123118
rect 509190 123042 509250 123118
rect 518942 123118 528570 123178
rect 509190 122982 518818 123042
rect 499438 122846 499682 122906
rect 518758 122906 518818 122982
rect 518942 122906 519002 123118
rect 528510 123042 528570 123118
rect 538262 123118 547890 123178
rect 528510 122982 538138 123042
rect 518758 122846 519002 122906
rect 538078 122906 538138 122982
rect 538262 122906 538322 123118
rect 547830 123042 547890 123118
rect 557582 123118 567210 123178
rect 547830 122982 557458 123042
rect 538078 122846 538322 122906
rect 557398 122906 557458 122982
rect 557582 122906 557642 123118
rect 567150 123042 567210 123118
rect 583342 123118 584960 123178
rect 583342 123042 583402 123118
rect 567150 122982 576778 123042
rect 557398 122846 557642 122906
rect 576718 122906 576778 122982
rect 576902 122982 583402 123042
rect 583520 123028 584960 123118
rect 576902 122906 576962 122982
rect 576718 122846 576962 122906
rect -960 122090 480 122180
rect 2773 122090 2839 122093
rect -960 122088 2839 122090
rect -960 122032 2778 122088
rect 2834 122032 2839 122088
rect -960 122030 2839 122032
rect -960 121940 480 122030
rect 2773 122027 2839 122030
rect 389265 118826 389331 118829
rect 389398 118826 389404 118828
rect 389265 118824 389404 118826
rect 389265 118768 389270 118824
rect 389326 118768 389404 118824
rect 389265 118766 389404 118768
rect 389265 118763 389331 118766
rect 389398 118764 389404 118766
rect 389468 118764 389474 118828
rect 259729 116106 259795 116109
rect 259686 116104 259795 116106
rect 259686 116048 259734 116104
rect 259790 116048 259795 116104
rect 259686 116043 259795 116048
rect 259686 115973 259746 116043
rect 244457 115970 244523 115973
rect 244641 115970 244707 115973
rect 244457 115968 244707 115970
rect 244457 115912 244462 115968
rect 244518 115912 244646 115968
rect 244702 115912 244707 115968
rect 244457 115910 244707 115912
rect 244457 115907 244523 115910
rect 244641 115907 244707 115910
rect 259637 115968 259746 115973
rect 259637 115912 259642 115968
rect 259698 115912 259746 115968
rect 259637 115910 259746 115912
rect 259637 115907 259703 115910
rect 374361 114746 374427 114749
rect 374318 114744 374427 114746
rect 374318 114688 374366 114744
rect 374422 114688 374427 114744
rect 374318 114683 374427 114688
rect 374318 114613 374378 114683
rect 374269 114608 374378 114613
rect 374269 114552 374274 114608
rect 374330 114552 374378 114608
rect 374269 114550 374378 114552
rect 374269 114547 374335 114550
rect 327257 113250 327323 113253
rect 327441 113250 327507 113253
rect 327257 113248 327507 113250
rect 327257 113192 327262 113248
rect 327318 113192 327446 113248
rect 327502 113192 327507 113248
rect 327257 113190 327507 113192
rect 327257 113187 327323 113190
rect 327441 113187 327507 113190
rect 583520 111482 584960 111572
rect 583342 111422 584960 111482
rect 317321 111074 317387 111077
rect 317321 111072 318810 111074
rect 317321 111016 317326 111072
rect 317382 111016 318810 111072
rect 317321 111014 318810 111016
rect 317321 111011 317387 111014
rect 318750 110938 318810 111014
rect 473302 111012 473308 111076
rect 473372 111074 473378 111076
rect 482921 111074 482987 111077
rect 473372 111072 482987 111074
rect 473372 111016 482926 111072
rect 482982 111016 482987 111072
rect 473372 111014 482987 111016
rect 473372 111012 473378 111014
rect 482921 111011 482987 111014
rect 328453 110938 328519 110941
rect 405406 110938 405412 110940
rect 318750 110878 321754 110938
rect 280061 110804 280127 110805
rect 243302 110740 243308 110804
rect 243372 110802 243378 110804
rect 243372 110742 254042 110802
rect 243372 110740 243378 110742
rect 253982 110666 254042 110742
rect 280061 110800 280108 110804
rect 280172 110802 280178 110804
rect 296662 110802 296668 110804
rect 280061 110744 280066 110800
rect 280061 110740 280108 110744
rect 280172 110742 280254 110802
rect 291886 110742 296668 110802
rect 280172 110740 280178 110742
rect 280061 110739 280127 110740
rect 291886 110666 291946 110742
rect 296662 110740 296668 110742
rect 296732 110740 296738 110804
rect 306281 110802 306347 110805
rect 307661 110802 307727 110805
rect 306281 110800 307727 110802
rect 306281 110744 306286 110800
rect 306342 110744 307666 110800
rect 307722 110744 307727 110800
rect 306281 110742 307727 110744
rect 306281 110739 306347 110742
rect 307661 110739 307727 110742
rect 253982 110606 265634 110666
rect 265574 110530 265634 110606
rect 285078 110606 291946 110666
rect 321694 110666 321754 110878
rect 328453 110936 328562 110938
rect 328453 110880 328458 110936
rect 328514 110880 328562 110936
rect 328453 110875 328562 110880
rect 328502 110802 328562 110875
rect 398606 110878 405412 110938
rect 328502 110742 340890 110802
rect 328453 110666 328519 110669
rect 321694 110664 328519 110666
rect 321694 110608 328458 110664
rect 328514 110608 328519 110664
rect 321694 110606 328519 110608
rect 270401 110530 270467 110533
rect 265574 110528 270467 110530
rect 265574 110472 270406 110528
rect 270462 110472 270467 110528
rect 265574 110470 270467 110472
rect 270401 110467 270467 110470
rect 278681 110530 278747 110533
rect 280061 110532 280127 110533
rect 280061 110530 280108 110532
rect 278681 110528 280108 110530
rect 280172 110530 280178 110532
rect 285078 110530 285138 110606
rect 328453 110603 328519 110606
rect 278681 110472 278686 110528
rect 278742 110472 280066 110528
rect 278681 110470 280108 110472
rect 278681 110467 278747 110470
rect 280061 110468 280108 110470
rect 280172 110470 285138 110530
rect 280172 110468 280178 110470
rect 296662 110468 296668 110532
rect 296732 110530 296738 110532
rect 306281 110530 306347 110533
rect 296732 110528 306347 110530
rect 296732 110472 306286 110528
rect 306342 110472 306347 110528
rect 296732 110470 306347 110472
rect 296732 110468 296738 110470
rect 280061 110467 280127 110468
rect 306281 110467 306347 110470
rect 315941 110530 316007 110533
rect 317321 110530 317387 110533
rect 315941 110528 317387 110530
rect 315941 110472 315946 110528
rect 316002 110472 317326 110528
rect 317382 110472 317387 110528
rect 315941 110470 317387 110472
rect 340830 110530 340890 110742
rect 365662 110740 365668 110804
rect 365732 110802 365738 110804
rect 365732 110742 379530 110802
rect 365732 110740 365738 110742
rect 357382 110666 357388 110668
rect 350582 110606 357388 110666
rect 350582 110530 350642 110606
rect 357382 110604 357388 110606
rect 357452 110604 357458 110668
rect 340830 110470 350642 110530
rect 379470 110530 379530 110742
rect 398606 110666 398666 110878
rect 405406 110876 405412 110878
rect 405476 110876 405482 110940
rect 487797 110938 487863 110941
rect 483062 110936 487863 110938
rect 483062 110880 487802 110936
rect 487858 110880 487863 110936
rect 483062 110878 487863 110880
rect 473302 110802 473308 110804
rect 466502 110742 473308 110802
rect 417877 110666 417943 110669
rect 389222 110606 398666 110666
rect 408542 110664 417943 110666
rect 408542 110608 417882 110664
rect 417938 110608 417943 110664
rect 408542 110606 417943 110608
rect 389222 110530 389282 110606
rect 379470 110470 389282 110530
rect 315941 110467 316007 110470
rect 317321 110467 317387 110470
rect 405590 110468 405596 110532
rect 405660 110530 405666 110532
rect 408542 110530 408602 110606
rect 417877 110603 417943 110606
rect 418153 110666 418219 110669
rect 437197 110666 437263 110669
rect 418153 110664 424978 110666
rect 418153 110608 418158 110664
rect 418214 110608 424978 110664
rect 418153 110606 424978 110608
rect 418153 110603 418219 110606
rect 405660 110470 408602 110530
rect 424918 110530 424978 110606
rect 427862 110664 437263 110666
rect 427862 110608 437202 110664
rect 437258 110608 437263 110664
rect 427862 110606 437263 110608
rect 427862 110530 427922 110606
rect 437197 110603 437263 110606
rect 437473 110666 437539 110669
rect 456517 110666 456583 110669
rect 437473 110664 444298 110666
rect 437473 110608 437478 110664
rect 437534 110608 444298 110664
rect 437473 110606 444298 110608
rect 437473 110603 437539 110606
rect 424918 110470 427922 110530
rect 444238 110530 444298 110606
rect 447182 110664 456583 110666
rect 447182 110608 456522 110664
rect 456578 110608 456583 110664
rect 447182 110606 456583 110608
rect 447182 110530 447242 110606
rect 456517 110603 456583 110606
rect 458817 110666 458883 110669
rect 458817 110664 463618 110666
rect 458817 110608 458822 110664
rect 458878 110608 463618 110664
rect 458817 110606 463618 110608
rect 458817 110603 458883 110606
rect 444238 110470 447242 110530
rect 463558 110530 463618 110606
rect 466502 110530 466562 110742
rect 473302 110740 473308 110742
rect 473372 110740 473378 110804
rect 482921 110666 482987 110669
rect 483062 110666 483122 110878
rect 487797 110875 487863 110878
rect 492622 110740 492628 110804
rect 492692 110802 492698 110804
rect 492692 110742 509250 110802
rect 492692 110740 492698 110742
rect 482921 110664 483122 110666
rect 482921 110608 482926 110664
rect 482982 110608 483122 110664
rect 482921 110606 483122 110608
rect 509190 110666 509250 110742
rect 518942 110742 528570 110802
rect 509190 110606 518818 110666
rect 482921 110603 482987 110606
rect 463558 110470 466562 110530
rect 487797 110530 487863 110533
rect 492622 110530 492628 110532
rect 487797 110528 492628 110530
rect 487797 110472 487802 110528
rect 487858 110472 492628 110528
rect 487797 110470 492628 110472
rect 405660 110468 405666 110470
rect 487797 110467 487863 110470
rect 492622 110468 492628 110470
rect 492692 110468 492698 110532
rect 518758 110530 518818 110606
rect 518942 110530 519002 110742
rect 528510 110666 528570 110742
rect 538262 110742 547890 110802
rect 528510 110606 538138 110666
rect 518758 110470 519002 110530
rect 538078 110530 538138 110606
rect 538262 110530 538322 110742
rect 547830 110666 547890 110742
rect 557582 110742 567210 110802
rect 547830 110606 557458 110666
rect 538078 110470 538322 110530
rect 557398 110530 557458 110606
rect 557582 110530 557642 110742
rect 567150 110666 567210 110742
rect 583342 110666 583402 111422
rect 583520 111332 584960 111422
rect 567150 110606 576778 110666
rect 557398 110470 557642 110530
rect 576718 110530 576778 110606
rect 576902 110606 583402 110666
rect 576902 110530 576962 110606
rect 576718 110470 576962 110530
rect 357382 110332 357388 110396
rect 357452 110394 357458 110396
rect 365662 110394 365668 110396
rect 357452 110334 365668 110394
rect 357452 110332 357458 110334
rect 365662 110332 365668 110334
rect 365732 110332 365738 110396
rect 389449 108900 389515 108901
rect 389398 108898 389404 108900
rect 389358 108838 389404 108898
rect 389468 108896 389515 108900
rect 389510 108840 389515 108896
rect 389398 108836 389404 108838
rect 389468 108836 389515 108840
rect 389449 108835 389515 108836
rect -960 107674 480 107764
rect 3509 107674 3575 107677
rect -960 107672 3575 107674
rect -960 107616 3514 107672
rect 3570 107616 3575 107672
rect -960 107614 3575 107616
rect -960 107524 480 107614
rect 3509 107611 3575 107614
rect 358721 106586 358787 106589
rect 358678 106584 358787 106586
rect 358678 106528 358726 106584
rect 358782 106528 358787 106584
rect 358678 106523 358787 106528
rect 358678 106317 358738 106523
rect 358678 106312 358787 106317
rect 358678 106256 358726 106312
rect 358782 106256 358787 106312
rect 358678 106254 358787 106256
rect 358721 106251 358787 106254
rect 324589 104818 324655 104821
rect 324454 104816 324655 104818
rect 324454 104760 324594 104816
rect 324650 104760 324655 104816
rect 324454 104758 324655 104760
rect 324454 104682 324514 104758
rect 324589 104755 324655 104758
rect 324773 104682 324839 104685
rect 324454 104680 324839 104682
rect 324454 104624 324778 104680
rect 324834 104624 324839 104680
rect 324454 104622 324839 104624
rect 324773 104619 324839 104622
rect 286041 103730 286107 103733
rect 285814 103728 286107 103730
rect 285814 103672 286046 103728
rect 286102 103672 286107 103728
rect 285814 103670 286107 103672
rect 285814 103594 285874 103670
rect 286041 103667 286107 103670
rect 285949 103594 286015 103597
rect 285814 103592 286015 103594
rect 285814 103536 285954 103592
rect 286010 103536 286015 103592
rect 285814 103534 286015 103536
rect 285949 103531 286015 103534
rect 327165 103458 327231 103461
rect 327030 103456 327231 103458
rect 327030 103400 327170 103456
rect 327226 103400 327231 103456
rect 327030 103398 327231 103400
rect 327030 103322 327090 103398
rect 327165 103395 327231 103398
rect 327441 103322 327507 103325
rect 327030 103320 327507 103322
rect 327030 103264 327446 103320
rect 327502 103264 327507 103320
rect 327030 103262 327507 103264
rect 327441 103259 327507 103262
rect 583520 99636 584960 99876
rect 247125 96794 247191 96797
rect 360377 96794 360443 96797
rect 367001 96794 367067 96797
rect 246990 96792 247191 96794
rect 246990 96736 247130 96792
rect 247186 96736 247191 96792
rect 246990 96734 247191 96736
rect 235073 96658 235139 96661
rect 235257 96658 235323 96661
rect 235073 96656 235323 96658
rect 235073 96600 235078 96656
rect 235134 96600 235262 96656
rect 235318 96600 235323 96656
rect 235073 96598 235323 96600
rect 246990 96658 247050 96734
rect 247125 96731 247191 96734
rect 360334 96792 360443 96794
rect 360334 96736 360382 96792
rect 360438 96736 360443 96792
rect 360334 96731 360443 96736
rect 366958 96792 367067 96794
rect 366958 96736 367006 96792
rect 367062 96736 367067 96792
rect 366958 96731 367067 96736
rect 360334 96661 360394 96731
rect 247125 96658 247191 96661
rect 246990 96656 247191 96658
rect 246990 96600 247130 96656
rect 247186 96600 247191 96656
rect 246990 96598 247191 96600
rect 235073 96595 235139 96598
rect 235257 96595 235323 96598
rect 247125 96595 247191 96598
rect 259545 96658 259611 96661
rect 259729 96658 259795 96661
rect 259545 96656 259795 96658
rect 259545 96600 259550 96656
rect 259606 96600 259734 96656
rect 259790 96600 259795 96656
rect 259545 96598 259795 96600
rect 259545 96595 259611 96598
rect 259729 96595 259795 96598
rect 360285 96656 360394 96661
rect 360285 96600 360290 96656
rect 360346 96600 360394 96656
rect 360285 96598 360394 96600
rect 366958 96661 367018 96731
rect 366958 96656 367067 96661
rect 366958 96600 367006 96656
rect 367062 96600 367067 96656
rect 366958 96598 367067 96600
rect 360285 96595 360351 96598
rect 367001 96595 367067 96598
rect 265157 96388 265223 96389
rect 265157 96386 265204 96388
rect 265112 96384 265204 96386
rect 265112 96328 265162 96384
rect 265112 96326 265204 96328
rect 265157 96324 265204 96326
rect 265268 96324 265274 96388
rect 265157 96323 265223 96324
rect 306833 93938 306899 93941
rect 307017 93938 307083 93941
rect 306833 93936 307083 93938
rect 306833 93880 306838 93936
rect 306894 93880 307022 93936
rect 307078 93880 307083 93936
rect 306833 93878 307083 93880
rect 306833 93875 306899 93878
rect 307017 93875 307083 93878
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 265249 89044 265315 89045
rect 265198 89042 265204 89044
rect 265158 88982 265204 89042
rect 265268 89040 265315 89044
rect 265310 88984 265315 89040
rect 265198 88980 265204 88982
rect 265268 88980 265315 88984
rect 265249 88979 265315 88980
rect 583520 87954 584960 88044
rect 583342 87894 584960 87954
rect 396022 87484 396028 87548
rect 396092 87546 396098 87548
rect 405590 87546 405596 87548
rect 396092 87486 405596 87546
rect 396092 87484 396098 87486
rect 405590 87484 405596 87486
rect 405660 87484 405666 87548
rect 299422 87348 299428 87412
rect 299492 87410 299498 87412
rect 304257 87410 304323 87413
rect 299492 87408 304323 87410
rect 299492 87352 304262 87408
rect 304318 87352 304323 87408
rect 299492 87350 304323 87352
rect 299492 87348 299498 87350
rect 304257 87347 304323 87350
rect 481582 87348 481588 87412
rect 481652 87410 481658 87412
rect 491201 87410 491267 87413
rect 481652 87408 491267 87410
rect 481652 87352 491206 87408
rect 491262 87352 491267 87408
rect 481652 87350 491267 87352
rect 481652 87348 481658 87350
rect 491201 87347 491267 87350
rect 251214 87274 251220 87276
rect 244414 87214 251220 87274
rect 244414 87138 244474 87214
rect 251214 87212 251220 87214
rect 251284 87212 251290 87276
rect 282913 87274 282979 87277
rect 282913 87272 283114 87274
rect 282913 87216 282918 87272
rect 282974 87216 283114 87272
rect 282913 87214 283114 87216
rect 282913 87211 282979 87214
rect 241654 87104 244106 87138
rect 244230 87104 244474 87138
rect 241470 87078 244474 87104
rect 251173 87140 251239 87141
rect 251173 87136 251220 87140
rect 251284 87138 251290 87140
rect 260649 87138 260715 87141
rect 282821 87138 282887 87141
rect 251173 87080 251178 87136
rect 241470 87044 241714 87078
rect 244046 87044 244290 87078
rect 251173 87076 251220 87080
rect 251284 87078 251330 87138
rect 260649 87136 282887 87138
rect 260649 87080 260654 87136
rect 260710 87080 282826 87136
rect 282882 87080 282887 87136
rect 260649 87078 282887 87080
rect 283054 87138 283114 87214
rect 307702 87212 307708 87276
rect 307772 87274 307778 87276
rect 476021 87274 476087 87277
rect 307772 87214 323594 87274
rect 307772 87212 307778 87214
rect 299422 87138 299428 87140
rect 283054 87078 299428 87138
rect 251284 87076 251290 87078
rect 251173 87075 251239 87076
rect 260649 87075 260715 87078
rect 282821 87075 282887 87078
rect 299422 87076 299428 87078
rect 299492 87076 299498 87140
rect 323534 87138 323594 87214
rect 328502 87214 340890 87274
rect 328502 87138 328562 87214
rect 323534 87078 328562 87138
rect 239990 86940 239996 87004
rect 240060 87002 240066 87004
rect 241470 87002 241530 87044
rect 240060 86942 241530 87002
rect 304257 87002 304323 87005
rect 307702 87002 307708 87004
rect 304257 87000 307708 87002
rect 304257 86944 304262 87000
rect 304318 86944 307708 87000
rect 304257 86942 307708 86944
rect 240060 86940 240066 86942
rect 304257 86939 304323 86942
rect 307702 86940 307708 86942
rect 307772 86940 307778 87004
rect 340830 87002 340890 87214
rect 466502 87272 476087 87274
rect 466502 87216 476026 87272
rect 476082 87216 476087 87272
rect 466502 87214 476087 87216
rect 357382 87138 357388 87140
rect 350582 87078 357388 87138
rect 350582 87002 350642 87078
rect 357382 87076 357388 87078
rect 357452 87076 357458 87140
rect 376753 87138 376819 87141
rect 369902 87136 376819 87138
rect 369902 87080 376758 87136
rect 376814 87080 376819 87136
rect 369902 87078 376819 87080
rect 340830 86942 350642 87002
rect 357566 86940 357572 87004
rect 357636 87002 357642 87004
rect 369902 87002 369962 87078
rect 376753 87075 376819 87078
rect 395981 87140 396047 87141
rect 395981 87136 396028 87140
rect 396092 87138 396098 87140
rect 417877 87138 417943 87141
rect 395981 87080 395986 87136
rect 395981 87076 396028 87080
rect 396092 87078 396174 87138
rect 408542 87136 417943 87138
rect 408542 87080 417882 87136
rect 417938 87080 417943 87136
rect 408542 87078 417943 87080
rect 396092 87076 396098 87078
rect 395981 87075 396047 87076
rect 357636 86942 369962 87002
rect 386229 87002 386295 87005
rect 386413 87002 386479 87005
rect 386229 87000 386479 87002
rect 386229 86944 386234 87000
rect 386290 86944 386418 87000
rect 386474 86944 386479 87000
rect 386229 86942 386479 86944
rect 357636 86940 357642 86942
rect 386229 86939 386295 86942
rect 386413 86939 386479 86942
rect 405590 86940 405596 87004
rect 405660 87002 405666 87004
rect 408542 87002 408602 87078
rect 417877 87075 417943 87078
rect 418153 87138 418219 87141
rect 437197 87138 437263 87141
rect 418153 87136 424978 87138
rect 418153 87080 418158 87136
rect 418214 87080 424978 87136
rect 418153 87078 424978 87080
rect 418153 87075 418219 87078
rect 405660 86942 408602 87002
rect 424918 87002 424978 87078
rect 427862 87136 437263 87138
rect 427862 87080 437202 87136
rect 437258 87080 437263 87136
rect 427862 87078 437263 87080
rect 427862 87002 427922 87078
rect 437197 87075 437263 87078
rect 437473 87138 437539 87141
rect 456517 87138 456583 87141
rect 437473 87136 444298 87138
rect 437473 87080 437478 87136
rect 437534 87080 444298 87136
rect 437473 87078 444298 87080
rect 437473 87075 437539 87078
rect 424918 86942 427922 87002
rect 444238 87002 444298 87078
rect 447182 87136 456583 87138
rect 447182 87080 456522 87136
rect 456578 87080 456583 87136
rect 447182 87078 456583 87080
rect 447182 87002 447242 87078
rect 456517 87075 456583 87078
rect 456977 87138 457043 87141
rect 456977 87136 463618 87138
rect 456977 87080 456982 87136
rect 457038 87080 463618 87136
rect 456977 87078 463618 87080
rect 456977 87075 457043 87078
rect 444238 86942 447242 87002
rect 463558 87002 463618 87078
rect 466502 87002 466562 87214
rect 476021 87211 476087 87214
rect 502241 87274 502307 87277
rect 502241 87272 509250 87274
rect 502241 87216 502246 87272
rect 502302 87216 509250 87272
rect 502241 87214 509250 87216
rect 502241 87211 502307 87214
rect 476205 87138 476271 87141
rect 481582 87138 481588 87140
rect 476205 87136 481588 87138
rect 476205 87080 476210 87136
rect 476266 87080 481588 87136
rect 476205 87078 481588 87080
rect 476205 87075 476271 87078
rect 481582 87076 481588 87078
rect 481652 87076 481658 87140
rect 509190 87138 509250 87214
rect 518942 87214 528570 87274
rect 509190 87078 518818 87138
rect 463558 86942 466562 87002
rect 491201 87002 491267 87005
rect 494605 87002 494671 87005
rect 491201 87000 494671 87002
rect 491201 86944 491206 87000
rect 491262 86944 494610 87000
rect 494666 86944 494671 87000
rect 491201 86942 494671 86944
rect 518758 87002 518818 87078
rect 518942 87002 519002 87214
rect 528510 87138 528570 87214
rect 538262 87214 547890 87274
rect 528510 87078 538138 87138
rect 518758 86942 519002 87002
rect 538078 87002 538138 87078
rect 538262 87002 538322 87214
rect 547830 87138 547890 87214
rect 557582 87214 567210 87274
rect 547830 87078 557458 87138
rect 538078 86942 538322 87002
rect 557398 87002 557458 87078
rect 557582 87002 557642 87214
rect 567150 87138 567210 87214
rect 583342 87138 583402 87894
rect 583520 87804 584960 87894
rect 567150 87078 576778 87138
rect 557398 86942 557642 87002
rect 576718 87002 576778 87078
rect 576902 87078 583402 87138
rect 576902 87002 576962 87078
rect 576718 86942 576962 87002
rect 405660 86940 405666 86942
rect 491201 86939 491267 86942
rect 494605 86939 494671 86942
rect 267825 82922 267891 82925
rect 268101 82922 268167 82925
rect 267825 82920 268167 82922
rect 267825 82864 267830 82920
rect 267886 82864 268106 82920
rect 268162 82864 268167 82920
rect 267825 82862 268167 82864
rect 267825 82859 267891 82862
rect 268101 82859 268167 82862
rect 267825 81426 267891 81429
rect 268009 81426 268075 81429
rect 267825 81424 268075 81426
rect 267825 81368 267830 81424
rect 267886 81368 268014 81424
rect 268070 81368 268075 81424
rect 267825 81366 268075 81368
rect 267825 81363 267891 81366
rect 268009 81363 268075 81366
rect -960 78978 480 79068
rect 2773 78978 2839 78981
rect -960 78976 2839 78978
rect -960 78920 2778 78976
rect 2834 78920 2839 78976
rect -960 78918 2839 78920
rect -960 78828 480 78918
rect 2773 78915 2839 78918
rect 376702 76468 376708 76532
rect 376772 76530 376778 76532
rect 395838 76530 395844 76532
rect 376772 76470 395844 76530
rect 376772 76468 376778 76470
rect 395838 76468 395844 76470
rect 395908 76468 395914 76532
rect 473302 76468 473308 76532
rect 473372 76530 473378 76532
rect 482921 76530 482987 76533
rect 473372 76528 482987 76530
rect 473372 76472 482926 76528
rect 482982 76472 482987 76528
rect 473372 76470 482987 76472
rect 473372 76468 473378 76470
rect 482921 76467 482987 76470
rect 487797 76394 487863 76397
rect 483062 76392 487863 76394
rect 483062 76336 487802 76392
rect 487858 76336 487863 76392
rect 483062 76334 487863 76336
rect 309041 76258 309107 76261
rect 299614 76256 309107 76258
rect 299614 76200 309046 76256
rect 309102 76200 309107 76256
rect 299614 76198 309107 76200
rect 241278 76060 241284 76124
rect 241348 76122 241354 76124
rect 253841 76122 253907 76125
rect 299614 76122 299674 76198
rect 309041 76195 309107 76198
rect 317321 76258 317387 76261
rect 318701 76258 318767 76261
rect 473302 76258 473308 76260
rect 317321 76256 318767 76258
rect 317321 76200 317326 76256
rect 317382 76200 318706 76256
rect 318762 76200 318767 76256
rect 317321 76198 318767 76200
rect 317321 76195 317387 76198
rect 318701 76195 318767 76198
rect 331078 76198 340890 76258
rect 241348 76120 253907 76122
rect 241348 76064 253846 76120
rect 253902 76064 253907 76120
rect 241348 76062 253907 76064
rect 241348 76060 241354 76062
rect 253841 76059 253907 76062
rect 299430 76062 299674 76122
rect 249793 75986 249859 75989
rect 250069 75986 250135 75989
rect 249793 75984 250135 75986
rect 249793 75928 249798 75984
rect 249854 75928 250074 75984
rect 250130 75928 250135 75984
rect 249793 75926 250135 75928
rect 249793 75923 249859 75926
rect 250069 75923 250135 75926
rect 259361 75986 259427 75989
rect 299430 75986 299490 76062
rect 259361 75984 282746 75986
rect 259361 75928 259366 75984
rect 259422 75928 282746 75984
rect 259361 75926 282746 75928
rect 259361 75923 259427 75926
rect 282686 75884 282746 75926
rect 283054 75926 299490 75986
rect 318701 75986 318767 75989
rect 331078 75986 331138 76198
rect 318701 75984 331138 75986
rect 318701 75928 318706 75984
rect 318762 75928 331138 75984
rect 318701 75926 331138 75928
rect 340830 75986 340890 76198
rect 466502 76198 473308 76258
rect 376702 76122 376708 76124
rect 350582 76062 369778 76122
rect 350582 75986 350642 76062
rect 340830 75926 350642 75986
rect 369718 75986 369778 76062
rect 369902 76062 376708 76122
rect 369902 75986 369962 76062
rect 376702 76060 376708 76062
rect 376772 76060 376778 76124
rect 395838 76060 395844 76124
rect 395908 76122 395914 76124
rect 398649 76122 398715 76125
rect 395908 76120 398715 76122
rect 395908 76064 398654 76120
rect 398710 76064 398715 76120
rect 395908 76062 398715 76064
rect 395908 76060 395914 76062
rect 398649 76059 398715 76062
rect 398833 76122 398899 76125
rect 417877 76122 417943 76125
rect 398833 76120 405658 76122
rect 398833 76064 398838 76120
rect 398894 76064 405658 76120
rect 398833 76062 405658 76064
rect 398833 76059 398899 76062
rect 369718 75926 369962 75986
rect 405598 75986 405658 76062
rect 408542 76120 417943 76122
rect 408542 76064 417882 76120
rect 417938 76064 417943 76120
rect 408542 76062 417943 76064
rect 408542 75986 408602 76062
rect 417877 76059 417943 76062
rect 420361 76122 420427 76125
rect 437197 76122 437263 76125
rect 420361 76120 424978 76122
rect 420361 76064 420366 76120
rect 420422 76064 424978 76120
rect 420361 76062 424978 76064
rect 420361 76059 420427 76062
rect 405598 75926 408602 75986
rect 424918 75986 424978 76062
rect 427862 76120 437263 76122
rect 427862 76064 437202 76120
rect 437258 76064 437263 76120
rect 427862 76062 437263 76064
rect 427862 75986 427922 76062
rect 437197 76059 437263 76062
rect 437473 76122 437539 76125
rect 456517 76122 456583 76125
rect 437473 76120 444298 76122
rect 437473 76064 437478 76120
rect 437534 76064 444298 76120
rect 437473 76062 444298 76064
rect 437473 76059 437539 76062
rect 424918 75926 427922 75986
rect 444238 75986 444298 76062
rect 447182 76120 456583 76122
rect 447182 76064 456522 76120
rect 456578 76064 456583 76120
rect 447182 76062 456583 76064
rect 447182 75986 447242 76062
rect 456517 76059 456583 76062
rect 456793 76122 456859 76125
rect 456793 76120 463618 76122
rect 456793 76064 456798 76120
rect 456854 76064 463618 76120
rect 456793 76062 463618 76064
rect 456793 76059 456859 76062
rect 444238 75926 447242 75986
rect 463558 75986 463618 76062
rect 466502 75986 466562 76198
rect 473302 76196 473308 76198
rect 473372 76196 473378 76260
rect 482921 76122 482987 76125
rect 483062 76122 483122 76334
rect 487797 76331 487863 76334
rect 492622 76196 492628 76260
rect 492692 76258 492698 76260
rect 583520 76258 584960 76348
rect 492692 76198 509250 76258
rect 492692 76196 492698 76198
rect 482921 76120 483122 76122
rect 482921 76064 482926 76120
rect 482982 76064 483122 76120
rect 482921 76062 483122 76064
rect 509190 76122 509250 76198
rect 518942 76198 528570 76258
rect 509190 76062 518818 76122
rect 482921 76059 482987 76062
rect 463558 75926 466562 75986
rect 487797 75986 487863 75989
rect 492622 75986 492628 75988
rect 487797 75984 492628 75986
rect 487797 75928 487802 75984
rect 487858 75928 492628 75984
rect 487797 75926 492628 75928
rect 283054 75884 283114 75926
rect 318701 75923 318767 75926
rect 487797 75923 487863 75926
rect 492622 75924 492628 75926
rect 492692 75924 492698 75988
rect 518758 75986 518818 76062
rect 518942 75986 519002 76198
rect 528510 76122 528570 76198
rect 538262 76198 547890 76258
rect 528510 76062 538138 76122
rect 518758 75926 519002 75986
rect 538078 75986 538138 76062
rect 538262 75986 538322 76198
rect 547830 76122 547890 76198
rect 557582 76198 567210 76258
rect 547830 76062 557458 76122
rect 538078 75926 538322 75986
rect 557398 75986 557458 76062
rect 557582 75986 557642 76198
rect 567150 76122 567210 76198
rect 583342 76198 584960 76258
rect 583342 76122 583402 76198
rect 567150 76062 576778 76122
rect 557398 75926 557642 75986
rect 576718 75986 576778 76062
rect 576902 76062 583402 76122
rect 583520 76108 584960 76198
rect 576902 75986 576962 76062
rect 576718 75926 576962 75986
rect 282686 75824 283114 75884
rect 310789 67826 310855 67829
rect 310654 67824 310855 67826
rect 310654 67768 310794 67824
rect 310850 67768 310855 67824
rect 310654 67766 310855 67768
rect 310654 67690 310714 67766
rect 310789 67763 310855 67766
rect 310789 67690 310855 67693
rect 310654 67688 310855 67690
rect 310654 67632 310794 67688
rect 310850 67632 310855 67688
rect 310654 67630 310855 67632
rect 310789 67627 310855 67630
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect 583520 64562 584960 64652
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 583342 64502 584960 64562
rect 287094 63956 287100 64020
rect 287164 64018 287170 64020
rect 296621 64018 296687 64021
rect 405406 64018 405412 64020
rect 287164 64016 296687 64018
rect 287164 63960 296626 64016
rect 296682 63960 296687 64016
rect 287164 63958 296687 63960
rect 287164 63956 287170 63958
rect 296621 63955 296687 63958
rect 398606 63958 405412 64018
rect 327022 63820 327028 63884
rect 327092 63882 327098 63884
rect 360193 63882 360259 63885
rect 327092 63822 340890 63882
rect 327092 63820 327098 63822
rect 278681 63746 278747 63749
rect 287094 63746 287100 63748
rect 278681 63744 287100 63746
rect 278681 63688 278686 63744
rect 278742 63688 287100 63744
rect 278681 63686 287100 63688
rect 278681 63683 278747 63686
rect 287094 63684 287100 63686
rect 287164 63684 287170 63748
rect 237230 63548 237236 63612
rect 237300 63610 237306 63612
rect 273161 63610 273227 63613
rect 237300 63608 273227 63610
rect 237300 63552 273166 63608
rect 273222 63552 273227 63608
rect 237300 63550 273227 63552
rect 237300 63548 237306 63550
rect 273161 63547 273227 63550
rect 296621 63610 296687 63613
rect 327022 63610 327028 63612
rect 296621 63608 307770 63610
rect 296621 63552 296626 63608
rect 296682 63552 307770 63608
rect 296621 63550 307770 63552
rect 296621 63547 296687 63550
rect 307710 63338 307770 63550
rect 317278 63550 327028 63610
rect 317278 63338 317338 63550
rect 327022 63548 327028 63550
rect 327092 63548 327098 63612
rect 340830 63610 340890 63822
rect 360193 63880 360394 63882
rect 360193 63824 360198 63880
rect 360254 63824 360394 63880
rect 360193 63822 360394 63824
rect 360193 63819 360259 63822
rect 360101 63746 360167 63749
rect 350582 63744 360167 63746
rect 350582 63688 360106 63744
rect 360162 63688 360167 63744
rect 350582 63686 360167 63688
rect 360334 63746 360394 63822
rect 398606 63746 398666 63958
rect 405406 63956 405412 63958
rect 405476 63956 405482 64020
rect 470550 63822 480178 63882
rect 417877 63746 417943 63749
rect 360334 63686 369778 63746
rect 350582 63610 350642 63686
rect 360101 63683 360167 63686
rect 340830 63550 350642 63610
rect 369718 63610 369778 63686
rect 389222 63686 398666 63746
rect 408542 63744 417943 63746
rect 408542 63688 417882 63744
rect 417938 63688 417943 63744
rect 408542 63686 417943 63688
rect 389222 63610 389282 63686
rect 369718 63550 389282 63610
rect 405590 63548 405596 63612
rect 405660 63610 405666 63612
rect 408542 63610 408602 63686
rect 417877 63683 417943 63686
rect 418153 63746 418219 63749
rect 437197 63746 437263 63749
rect 418153 63744 424978 63746
rect 418153 63688 418158 63744
rect 418214 63688 424978 63744
rect 418153 63686 424978 63688
rect 418153 63683 418219 63686
rect 405660 63550 408602 63610
rect 424918 63610 424978 63686
rect 427862 63744 437263 63746
rect 427862 63688 437202 63744
rect 437258 63688 437263 63744
rect 427862 63686 437263 63688
rect 427862 63610 427922 63686
rect 437197 63683 437263 63686
rect 437473 63746 437539 63749
rect 456517 63746 456583 63749
rect 437473 63744 444298 63746
rect 437473 63688 437478 63744
rect 437534 63688 444298 63744
rect 437473 63686 444298 63688
rect 437473 63683 437539 63686
rect 424918 63550 427922 63610
rect 444238 63610 444298 63686
rect 447182 63744 456583 63746
rect 447182 63688 456522 63744
rect 456578 63688 456583 63744
rect 447182 63686 456583 63688
rect 447182 63610 447242 63686
rect 456517 63683 456583 63686
rect 456885 63746 456951 63749
rect 456885 63744 466378 63746
rect 456885 63688 456890 63744
rect 456946 63688 466378 63744
rect 456885 63686 466378 63688
rect 456885 63683 456951 63686
rect 444238 63550 447242 63610
rect 466318 63610 466378 63686
rect 470550 63610 470610 63822
rect 466318 63550 470610 63610
rect 480118 63610 480178 63822
rect 480302 63822 489930 63882
rect 480302 63610 480362 63822
rect 489870 63746 489930 63822
rect 499622 63822 509250 63882
rect 489870 63686 499498 63746
rect 480118 63550 480362 63610
rect 499438 63610 499498 63686
rect 499622 63610 499682 63822
rect 509190 63746 509250 63822
rect 518942 63822 528570 63882
rect 509190 63686 518818 63746
rect 499438 63550 499682 63610
rect 518758 63610 518818 63686
rect 518942 63610 519002 63822
rect 528510 63746 528570 63822
rect 538262 63822 547890 63882
rect 528510 63686 538138 63746
rect 518758 63550 519002 63610
rect 538078 63610 538138 63686
rect 538262 63610 538322 63822
rect 547830 63746 547890 63822
rect 557582 63822 567210 63882
rect 547830 63686 557458 63746
rect 538078 63550 538322 63610
rect 557398 63610 557458 63686
rect 557582 63610 557642 63822
rect 567150 63746 567210 63822
rect 583342 63746 583402 64502
rect 583520 64412 584960 64502
rect 567150 63686 576778 63746
rect 557398 63550 557642 63610
rect 576718 63610 576778 63686
rect 576902 63686 583402 63746
rect 576902 63610 576962 63686
rect 576718 63550 576962 63610
rect 405660 63548 405666 63550
rect 307710 63278 317338 63338
rect 267825 62114 267891 62117
rect 268009 62114 268075 62117
rect 267825 62112 268075 62114
rect 267825 62056 267830 62112
rect 267886 62056 268014 62112
rect 268070 62056 268075 62112
rect 267825 62054 268075 62056
rect 267825 62051 267891 62054
rect 268009 62051 268075 62054
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 2773 50146 2839 50149
rect -960 50144 2839 50146
rect -960 50088 2778 50144
rect 2834 50088 2839 50144
rect -960 50086 2839 50088
rect -960 49996 480 50086
rect 2773 50083 2839 50086
rect 329925 48378 329991 48381
rect 330109 48378 330175 48381
rect 329925 48376 330175 48378
rect 329925 48320 329930 48376
rect 329986 48320 330114 48376
rect 330170 48320 330175 48376
rect 329925 48318 330175 48320
rect 329925 48315 329991 48318
rect 330109 48315 330175 48318
rect 244365 44162 244431 44165
rect 244549 44162 244615 44165
rect 244365 44160 244615 44162
rect 244365 44104 244370 44160
rect 244426 44104 244554 44160
rect 244610 44104 244615 44160
rect 244365 44102 244615 44104
rect 244365 44099 244431 44102
rect 244549 44099 244615 44102
rect 583520 41034 584960 41124
rect 583342 40974 584960 41034
rect 396030 40430 405658 40490
rect 241421 40354 241487 40357
rect 239998 40352 241487 40354
rect 239998 40296 241426 40352
rect 241482 40296 241487 40352
rect 239998 40294 241487 40296
rect 232998 40156 233004 40220
rect 233068 40218 233074 40220
rect 239998 40218 240058 40294
rect 241421 40291 241487 40294
rect 327022 40292 327028 40356
rect 327092 40354 327098 40356
rect 327092 40294 340890 40354
rect 327092 40292 327098 40294
rect 282729 40218 282795 40221
rect 233068 40158 240058 40218
rect 271094 40216 282795 40218
rect 271094 40160 282734 40216
rect 282790 40160 282795 40216
rect 271094 40158 282795 40160
rect 233068 40156 233074 40158
rect 245009 40082 245075 40085
rect 253841 40082 253907 40085
rect 245009 40080 253907 40082
rect 245009 40024 245014 40080
rect 245070 40024 253846 40080
rect 253902 40024 253907 40080
rect 245009 40022 253907 40024
rect 245009 40019 245075 40022
rect 253841 40019 253907 40022
rect 262857 40082 262923 40085
rect 271094 40082 271154 40158
rect 282729 40155 282795 40158
rect 282913 40218 282979 40221
rect 282913 40216 312002 40218
rect 282913 40160 282918 40216
rect 282974 40160 312002 40216
rect 282913 40158 312002 40160
rect 282913 40155 282979 40158
rect 262857 40080 271154 40082
rect 262857 40024 262862 40080
rect 262918 40024 271154 40080
rect 262857 40022 271154 40024
rect 311942 40082 312002 40158
rect 327022 40082 327028 40084
rect 311942 40022 327028 40082
rect 262857 40019 262923 40022
rect 327022 40020 327028 40022
rect 327092 40020 327098 40084
rect 340830 40082 340890 40294
rect 360101 40218 360167 40221
rect 350582 40216 360167 40218
rect 350582 40160 360106 40216
rect 360162 40160 360167 40216
rect 350582 40158 360167 40160
rect 350582 40082 350642 40158
rect 360101 40155 360167 40158
rect 360285 40218 360351 40221
rect 396030 40218 396090 40430
rect 405598 40356 405658 40430
rect 405590 40292 405596 40356
rect 405660 40292 405666 40356
rect 470550 40294 480178 40354
rect 417877 40218 417943 40221
rect 360285 40216 369778 40218
rect 360285 40160 360290 40216
rect 360346 40160 369778 40216
rect 360285 40158 369778 40160
rect 360285 40155 360351 40158
rect 340830 40022 350642 40082
rect 369718 40082 369778 40158
rect 389222 40158 396090 40218
rect 408542 40216 417943 40218
rect 408542 40160 417882 40216
rect 417938 40160 417943 40216
rect 408542 40158 417943 40160
rect 389222 40082 389282 40158
rect 369718 40022 389282 40082
rect 405590 40020 405596 40084
rect 405660 40082 405666 40084
rect 408542 40082 408602 40158
rect 417877 40155 417943 40158
rect 420361 40218 420427 40221
rect 437197 40218 437263 40221
rect 420361 40216 424978 40218
rect 420361 40160 420366 40216
rect 420422 40160 424978 40216
rect 420361 40158 424978 40160
rect 420361 40155 420427 40158
rect 405660 40022 408602 40082
rect 424918 40082 424978 40158
rect 427862 40216 437263 40218
rect 427862 40160 437202 40216
rect 437258 40160 437263 40216
rect 427862 40158 437263 40160
rect 427862 40082 427922 40158
rect 437197 40155 437263 40158
rect 437473 40218 437539 40221
rect 456517 40218 456583 40221
rect 437473 40216 444298 40218
rect 437473 40160 437478 40216
rect 437534 40160 444298 40216
rect 437473 40158 444298 40160
rect 437473 40155 437539 40158
rect 424918 40022 427922 40082
rect 444238 40082 444298 40158
rect 447182 40216 456583 40218
rect 447182 40160 456522 40216
rect 456578 40160 456583 40216
rect 447182 40158 456583 40160
rect 447182 40082 447242 40158
rect 456517 40155 456583 40158
rect 456885 40218 456951 40221
rect 456885 40216 466378 40218
rect 456885 40160 456890 40216
rect 456946 40160 466378 40216
rect 456885 40158 466378 40160
rect 456885 40155 456951 40158
rect 444238 40022 447242 40082
rect 466318 40082 466378 40158
rect 470550 40082 470610 40294
rect 466318 40022 470610 40082
rect 480118 40082 480178 40294
rect 480302 40294 489930 40354
rect 480302 40082 480362 40294
rect 489870 40218 489930 40294
rect 499622 40294 509250 40354
rect 489870 40158 499498 40218
rect 480118 40022 480362 40082
rect 499438 40082 499498 40158
rect 499622 40082 499682 40294
rect 509190 40218 509250 40294
rect 518942 40294 528570 40354
rect 509190 40158 518818 40218
rect 499438 40022 499682 40082
rect 518758 40082 518818 40158
rect 518942 40082 519002 40294
rect 528510 40218 528570 40294
rect 538262 40294 547890 40354
rect 528510 40158 538138 40218
rect 518758 40022 519002 40082
rect 538078 40082 538138 40158
rect 538262 40082 538322 40294
rect 547830 40218 547890 40294
rect 557582 40294 567210 40354
rect 547830 40158 557458 40218
rect 538078 40022 538322 40082
rect 557398 40082 557458 40158
rect 557582 40082 557642 40294
rect 567150 40218 567210 40294
rect 583342 40218 583402 40974
rect 583520 40884 584960 40974
rect 567150 40158 576778 40218
rect 557398 40022 557642 40082
rect 576718 40082 576778 40158
rect 576902 40158 583402 40218
rect 576902 40082 576962 40158
rect 576718 40022 576962 40082
rect 405660 40020 405666 40022
rect -960 35866 480 35956
rect 3141 35866 3207 35869
rect -960 35864 3207 35866
rect -960 35808 3146 35864
rect 3202 35808 3207 35864
rect -960 35806 3207 35808
rect -960 35716 480 35806
rect 3141 35803 3207 35806
rect 285622 29548 285628 29612
rect 285692 29610 285698 29612
rect 295241 29610 295307 29613
rect 331857 29610 331923 29613
rect 285692 29608 295307 29610
rect 285692 29552 295246 29608
rect 295302 29552 295307 29608
rect 285692 29550 295307 29552
rect 285692 29548 285698 29550
rect 295241 29547 295307 29550
rect 327030 29608 331923 29610
rect 327030 29552 331862 29608
rect 331918 29552 331923 29608
rect 327030 29550 331923 29552
rect 296621 29476 296687 29477
rect 296621 29472 296668 29476
rect 296732 29474 296738 29476
rect 296621 29416 296626 29472
rect 296621 29412 296668 29416
rect 296732 29414 296814 29474
rect 296732 29412 296738 29414
rect 296621 29411 296687 29412
rect 257889 29338 257955 29341
rect 258022 29338 258028 29340
rect 257889 29336 258028 29338
rect 257889 29280 257894 29336
rect 257950 29280 258028 29336
rect 257889 29278 258028 29280
rect 257889 29275 257955 29278
rect 258022 29276 258028 29278
rect 258092 29276 258098 29340
rect 262857 29338 262923 29341
rect 285622 29338 285628 29340
rect 262857 29336 285628 29338
rect 262857 29280 262862 29336
rect 262918 29280 285628 29336
rect 262857 29278 285628 29280
rect 262857 29275 262923 29278
rect 285622 29276 285628 29278
rect 285692 29276 285698 29340
rect 295241 29338 295307 29341
rect 296621 29338 296687 29341
rect 295241 29336 296687 29338
rect 295241 29280 295246 29336
rect 295302 29280 296626 29336
rect 296682 29280 296687 29336
rect 295241 29278 296687 29280
rect 295241 29275 295307 29278
rect 296621 29275 296687 29278
rect 317321 29338 317387 29341
rect 322197 29338 322263 29341
rect 327030 29338 327090 29550
rect 331857 29547 331923 29550
rect 396022 29548 396028 29612
rect 396092 29610 396098 29612
rect 396092 29550 405658 29610
rect 396092 29548 396098 29550
rect 405598 29476 405658 29550
rect 405590 29412 405596 29476
rect 405660 29412 405666 29476
rect 481582 29412 481588 29476
rect 481652 29474 481658 29476
rect 491201 29474 491267 29477
rect 481652 29472 491267 29474
rect 481652 29416 491206 29472
rect 491262 29416 491267 29472
rect 481652 29414 491267 29416
rect 481652 29412 481658 29414
rect 491201 29411 491267 29414
rect 317321 29336 317522 29338
rect 317321 29280 317326 29336
rect 317382 29280 317522 29336
rect 317321 29278 317522 29280
rect 317321 29275 317387 29278
rect 235758 29140 235764 29204
rect 235828 29202 235834 29204
rect 248413 29202 248479 29205
rect 235828 29200 248479 29202
rect 235828 29144 248418 29200
rect 248474 29144 248479 29200
rect 235828 29142 248479 29144
rect 235828 29140 235834 29142
rect 248413 29139 248479 29142
rect 296662 29140 296668 29204
rect 296732 29202 296738 29204
rect 306281 29202 306347 29205
rect 296732 29200 306347 29202
rect 296732 29144 306286 29200
rect 306342 29144 306347 29200
rect 296732 29142 306347 29144
rect 296732 29140 296738 29142
rect 306281 29139 306347 29142
rect 258022 29004 258028 29068
rect 258092 29066 258098 29068
rect 262857 29066 262923 29069
rect 258092 29064 262923 29066
rect 258092 29008 262862 29064
rect 262918 29008 262923 29064
rect 258092 29006 262923 29008
rect 317462 29066 317522 29278
rect 322197 29336 327090 29338
rect 322197 29280 322202 29336
rect 322258 29280 327090 29336
rect 322197 29278 327090 29280
rect 331857 29338 331923 29341
rect 376661 29338 376727 29341
rect 476021 29338 476087 29341
rect 331857 29336 340890 29338
rect 331857 29280 331862 29336
rect 331918 29280 340890 29336
rect 331857 29278 340890 29280
rect 322197 29275 322263 29278
rect 331857 29275 331923 29278
rect 322197 29066 322263 29069
rect 317462 29064 322263 29066
rect 317462 29008 322202 29064
rect 322258 29008 322263 29064
rect 317462 29006 322263 29008
rect 340830 29066 340890 29278
rect 376661 29336 379530 29338
rect 376661 29280 376666 29336
rect 376722 29280 379530 29336
rect 376661 29278 379530 29280
rect 376661 29275 376727 29278
rect 350582 29142 357450 29202
rect 350582 29066 350642 29142
rect 340830 29006 350642 29066
rect 357390 29100 357450 29142
rect 357390 29066 357634 29100
rect 367093 29066 367159 29069
rect 357390 29064 367159 29066
rect 357390 29040 367098 29064
rect 357574 29008 367098 29040
rect 367154 29008 367159 29064
rect 357574 29006 367159 29008
rect 258092 29004 258098 29006
rect 262857 29003 262923 29006
rect 322197 29003 322263 29006
rect 367093 29003 367159 29006
rect 377121 29066 377187 29069
rect 377305 29066 377371 29069
rect 377121 29064 377371 29066
rect 377121 29008 377126 29064
rect 377182 29008 377310 29064
rect 377366 29008 377371 29064
rect 377121 29006 377371 29008
rect 379470 29066 379530 29278
rect 466502 29336 476087 29338
rect 466502 29280 476026 29336
rect 476082 29280 476087 29336
rect 466502 29278 476087 29280
rect 396022 29202 396028 29204
rect 389222 29142 396028 29202
rect 389222 29066 389282 29142
rect 396022 29140 396028 29142
rect 396092 29140 396098 29204
rect 417877 29202 417943 29205
rect 408542 29200 417943 29202
rect 408542 29144 417882 29200
rect 417938 29144 417943 29200
rect 408542 29142 417943 29144
rect 379470 29006 389282 29066
rect 377121 29003 377187 29006
rect 377305 29003 377371 29006
rect 405590 29004 405596 29068
rect 405660 29066 405666 29068
rect 408542 29066 408602 29142
rect 417877 29139 417943 29142
rect 418797 29202 418863 29205
rect 437197 29202 437263 29205
rect 418797 29200 424978 29202
rect 418797 29144 418802 29200
rect 418858 29144 424978 29200
rect 418797 29142 424978 29144
rect 418797 29139 418863 29142
rect 405660 29006 408602 29066
rect 424918 29066 424978 29142
rect 427862 29200 437263 29202
rect 427862 29144 437202 29200
rect 437258 29144 437263 29200
rect 427862 29142 437263 29144
rect 427862 29066 427922 29142
rect 437197 29139 437263 29142
rect 437473 29202 437539 29205
rect 456517 29202 456583 29205
rect 437473 29200 444298 29202
rect 437473 29144 437478 29200
rect 437534 29144 444298 29200
rect 437473 29142 444298 29144
rect 437473 29139 437539 29142
rect 424918 29006 427922 29066
rect 444238 29066 444298 29142
rect 447182 29200 456583 29202
rect 447182 29144 456522 29200
rect 456578 29144 456583 29200
rect 447182 29142 456583 29144
rect 447182 29066 447242 29142
rect 456517 29139 456583 29142
rect 456977 29202 457043 29205
rect 456977 29200 463618 29202
rect 456977 29144 456982 29200
rect 457038 29144 463618 29200
rect 456977 29142 463618 29144
rect 456977 29139 457043 29142
rect 444238 29006 447242 29066
rect 463558 29066 463618 29142
rect 466502 29066 466562 29278
rect 476021 29275 476087 29278
rect 502241 29338 502307 29341
rect 583520 29338 584960 29428
rect 502241 29336 509250 29338
rect 502241 29280 502246 29336
rect 502302 29280 509250 29336
rect 502241 29278 509250 29280
rect 502241 29275 502307 29278
rect 476205 29202 476271 29205
rect 481582 29202 481588 29204
rect 476205 29200 481588 29202
rect 476205 29144 476210 29200
rect 476266 29144 481588 29200
rect 476205 29142 481588 29144
rect 476205 29139 476271 29142
rect 481582 29140 481588 29142
rect 481652 29140 481658 29204
rect 509190 29202 509250 29278
rect 518942 29278 528570 29338
rect 509190 29142 518818 29202
rect 463558 29006 466562 29066
rect 491201 29066 491267 29069
rect 492765 29066 492831 29069
rect 491201 29064 492831 29066
rect 491201 29008 491206 29064
rect 491262 29008 492770 29064
rect 492826 29008 492831 29064
rect 491201 29006 492831 29008
rect 518758 29066 518818 29142
rect 518942 29066 519002 29278
rect 528510 29202 528570 29278
rect 538262 29278 547890 29338
rect 528510 29142 538138 29202
rect 518758 29006 519002 29066
rect 538078 29066 538138 29142
rect 538262 29066 538322 29278
rect 547830 29202 547890 29278
rect 557582 29278 567210 29338
rect 547830 29142 557458 29202
rect 538078 29006 538322 29066
rect 557398 29066 557458 29142
rect 557582 29066 557642 29278
rect 567150 29202 567210 29278
rect 583342 29278 584960 29338
rect 583342 29202 583402 29278
rect 567150 29142 576778 29202
rect 557398 29006 557642 29066
rect 576718 29066 576778 29142
rect 576902 29142 583402 29202
rect 583520 29188 584960 29278
rect 576902 29066 576962 29142
rect 576718 29006 576962 29066
rect 405660 29004 405666 29006
rect 491201 29003 491267 29006
rect 492765 29003 492831 29006
rect 306281 28930 306347 28933
rect 307661 28930 307727 28933
rect 306281 28928 307727 28930
rect 306281 28872 306286 28928
rect 306342 28872 307666 28928
rect 307722 28872 307727 28928
rect 306281 28870 307727 28872
rect 306281 28867 306347 28870
rect 307661 28867 307727 28870
rect 315941 28930 316007 28933
rect 317321 28930 317387 28933
rect 315941 28928 317387 28930
rect 315941 28872 315946 28928
rect 316002 28872 317326 28928
rect 317382 28872 317387 28928
rect 315941 28870 317387 28872
rect 315941 28867 316007 28870
rect 317321 28867 317387 28870
rect 389449 22268 389515 22269
rect 389398 22266 389404 22268
rect 389358 22206 389404 22266
rect 389468 22264 389515 22268
rect 389510 22208 389515 22264
rect 389398 22204 389404 22206
rect 389468 22204 389515 22208
rect 389449 22203 389515 22204
rect 465574 21994 465580 21996
rect 614 21934 465580 21994
rect -960 21450 480 21540
rect 614 21450 674 21934
rect 465574 21932 465580 21934
rect 465644 21932 465650 21996
rect -960 21390 674 21450
rect -960 21300 480 21390
rect 251214 21388 251220 21452
rect 251284 21450 251290 21452
rect 251449 21450 251515 21453
rect 251284 21448 251515 21450
rect 251284 21392 251454 21448
rect 251510 21392 251515 21448
rect 251284 21390 251515 21392
rect 251284 21388 251290 21390
rect 251449 21387 251515 21390
rect 389357 18052 389423 18053
rect 389357 18050 389404 18052
rect 389312 18048 389404 18050
rect 389312 17992 389362 18048
rect 389312 17990 389404 17992
rect 389357 17988 389404 17990
rect 389468 17988 389474 18052
rect 389357 17987 389423 17988
rect 583520 17642 584960 17732
rect 583342 17582 584960 17642
rect 473302 17172 473308 17236
rect 473372 17234 473378 17236
rect 482921 17234 482987 17237
rect 473372 17232 482987 17234
rect 473372 17176 482926 17232
rect 482982 17176 482987 17232
rect 473372 17174 482987 17176
rect 473372 17172 473378 17174
rect 482921 17171 482987 17174
rect 405406 17098 405412 17100
rect 398606 17038 405412 17098
rect 338205 16962 338271 16965
rect 338205 16960 360210 16962
rect 338205 16904 338210 16960
rect 338266 16904 360210 16960
rect 338205 16902 360210 16904
rect 338205 16899 338271 16902
rect 231710 16764 231716 16828
rect 231780 16826 231786 16828
rect 241421 16826 241487 16829
rect 231780 16824 241487 16826
rect 231780 16768 241426 16824
rect 241482 16768 241487 16824
rect 231780 16766 241487 16768
rect 231780 16764 231786 16766
rect 241421 16763 241487 16766
rect 260966 16764 260972 16828
rect 261036 16826 261042 16828
rect 288341 16826 288407 16829
rect 298001 16826 298067 16829
rect 328269 16826 328335 16829
rect 261036 16766 273178 16826
rect 288260 16824 288450 16826
rect 288260 16768 288346 16824
rect 288402 16768 288450 16824
rect 288260 16766 288450 16768
rect 261036 16764 261042 16766
rect 241421 16690 241487 16693
rect 251081 16690 251147 16693
rect 241421 16688 251147 16690
rect 241421 16632 241426 16688
rect 241482 16632 251086 16688
rect 251142 16632 251147 16688
rect 241421 16630 251147 16632
rect 241421 16627 241487 16630
rect 251081 16627 251147 16630
rect 259361 16690 259427 16693
rect 260782 16690 260788 16692
rect 259361 16688 260788 16690
rect 259361 16632 259366 16688
rect 259422 16632 260788 16688
rect 259361 16630 260788 16632
rect 259361 16627 259427 16630
rect 260782 16628 260788 16630
rect 260852 16628 260858 16692
rect 273118 16588 273178 16766
rect 288341 16763 288450 16766
rect 298001 16824 298202 16826
rect 298001 16768 298006 16824
rect 298062 16768 298202 16824
rect 298001 16766 298202 16768
rect 298001 16763 298067 16766
rect 273302 16630 278882 16690
rect 273302 16588 273362 16630
rect 273118 16528 273362 16588
rect 278822 16554 278882 16630
rect 288390 16557 288450 16763
rect 288341 16554 288450 16557
rect 298001 16554 298067 16557
rect 278822 16552 298067 16554
rect 278822 16496 288346 16552
rect 288402 16496 298006 16552
rect 298062 16496 298067 16552
rect 278822 16494 298067 16496
rect 298142 16554 298202 16766
rect 327030 16824 328335 16826
rect 327030 16768 328274 16824
rect 328330 16768 328335 16824
rect 327030 16766 328335 16768
rect 360150 16826 360210 16902
rect 398606 16826 398666 17038
rect 405406 17036 405412 17038
rect 405476 17036 405482 17100
rect 487797 17098 487863 17101
rect 483062 17096 487863 17098
rect 483062 17040 487802 17096
rect 487858 17040 487863 17096
rect 483062 17038 487863 17040
rect 473302 16962 473308 16964
rect 466502 16902 473308 16962
rect 417877 16826 417943 16829
rect 360150 16766 369778 16826
rect 317321 16690 317387 16693
rect 322197 16690 322263 16693
rect 327030 16690 327090 16766
rect 328269 16763 328335 16766
rect 336733 16690 336799 16693
rect 317321 16688 317522 16690
rect 317321 16632 317326 16688
rect 317382 16632 317522 16688
rect 317321 16630 317522 16632
rect 317321 16627 317387 16630
rect 306414 16554 306420 16556
rect 298142 16494 306420 16554
rect 288341 16491 288407 16494
rect 298001 16491 298067 16494
rect 306414 16492 306420 16494
rect 306484 16492 306490 16556
rect 315941 16418 316007 16421
rect 317321 16418 317387 16421
rect 315941 16416 317387 16418
rect 315941 16360 315946 16416
rect 316002 16360 317326 16416
rect 317382 16360 317387 16416
rect 315941 16358 317387 16360
rect 317462 16418 317522 16630
rect 322197 16688 327090 16690
rect 322197 16632 322202 16688
rect 322258 16632 327090 16688
rect 322197 16630 327090 16632
rect 336598 16688 336799 16690
rect 336598 16632 336738 16688
rect 336794 16632 336799 16688
rect 336598 16630 336799 16632
rect 369718 16690 369778 16766
rect 389222 16766 398666 16826
rect 408542 16824 417943 16826
rect 408542 16768 417882 16824
rect 417938 16768 417943 16824
rect 408542 16766 417943 16768
rect 389222 16690 389282 16766
rect 369718 16630 389282 16690
rect 322197 16627 322263 16630
rect 328269 16554 328335 16557
rect 336598 16554 336658 16630
rect 336733 16627 336799 16630
rect 405590 16628 405596 16692
rect 405660 16690 405666 16692
rect 408542 16690 408602 16766
rect 417877 16763 417943 16766
rect 418153 16826 418219 16829
rect 437197 16826 437263 16829
rect 418153 16824 424978 16826
rect 418153 16768 418158 16824
rect 418214 16768 424978 16824
rect 418153 16766 424978 16768
rect 418153 16763 418219 16766
rect 405660 16630 408602 16690
rect 424918 16690 424978 16766
rect 427862 16824 437263 16826
rect 427862 16768 437202 16824
rect 437258 16768 437263 16824
rect 427862 16766 437263 16768
rect 427862 16690 427922 16766
rect 437197 16763 437263 16766
rect 437473 16826 437539 16829
rect 456517 16826 456583 16829
rect 437473 16824 444298 16826
rect 437473 16768 437478 16824
rect 437534 16768 444298 16824
rect 437473 16766 444298 16768
rect 437473 16763 437539 16766
rect 424918 16630 427922 16690
rect 444238 16690 444298 16766
rect 447182 16824 456583 16826
rect 447182 16768 456522 16824
rect 456578 16768 456583 16824
rect 447182 16766 456583 16768
rect 447182 16690 447242 16766
rect 456517 16763 456583 16766
rect 458817 16826 458883 16829
rect 458817 16824 463618 16826
rect 458817 16768 458822 16824
rect 458878 16768 463618 16824
rect 458817 16766 463618 16768
rect 458817 16763 458883 16766
rect 444238 16630 447242 16690
rect 463558 16690 463618 16766
rect 466502 16690 466562 16902
rect 473302 16900 473308 16902
rect 473372 16900 473378 16964
rect 482921 16826 482987 16829
rect 483062 16826 483122 17038
rect 487797 17035 487863 17038
rect 492622 16900 492628 16964
rect 492692 16962 492698 16964
rect 492692 16902 509250 16962
rect 492692 16900 492698 16902
rect 482921 16824 483122 16826
rect 482921 16768 482926 16824
rect 482982 16768 483122 16824
rect 482921 16766 483122 16768
rect 509190 16826 509250 16902
rect 518942 16902 528570 16962
rect 509190 16766 518818 16826
rect 482921 16763 482987 16766
rect 463558 16630 466562 16690
rect 487797 16690 487863 16693
rect 492622 16690 492628 16692
rect 487797 16688 492628 16690
rect 487797 16632 487802 16688
rect 487858 16632 492628 16688
rect 487797 16630 492628 16632
rect 405660 16628 405666 16630
rect 487797 16627 487863 16630
rect 492622 16628 492628 16630
rect 492692 16628 492698 16692
rect 518758 16690 518818 16766
rect 518942 16690 519002 16902
rect 528510 16826 528570 16902
rect 538262 16902 547890 16962
rect 528510 16766 538138 16826
rect 518758 16630 519002 16690
rect 538078 16690 538138 16766
rect 538262 16690 538322 16902
rect 547830 16826 547890 16902
rect 557582 16902 567210 16962
rect 547830 16766 557458 16826
rect 538078 16630 538322 16690
rect 557398 16690 557458 16766
rect 557582 16690 557642 16902
rect 567150 16826 567210 16902
rect 583342 16826 583402 17582
rect 583520 17492 584960 17582
rect 567150 16766 576778 16826
rect 557398 16630 557642 16690
rect 576718 16690 576778 16766
rect 576902 16766 583402 16826
rect 576902 16690 576962 16766
rect 576718 16630 576962 16690
rect 328269 16552 336658 16554
rect 328269 16496 328274 16552
rect 328330 16496 336658 16552
rect 328269 16494 336658 16496
rect 328269 16491 328335 16494
rect 322197 16418 322263 16421
rect 317462 16416 322263 16418
rect 317462 16360 322202 16416
rect 322258 16360 322263 16416
rect 317462 16358 322263 16360
rect 315941 16355 316007 16358
rect 317321 16355 317387 16358
rect 322197 16355 322263 16358
rect 306414 16084 306420 16148
rect 306484 16146 306490 16148
rect 315941 16146 316007 16149
rect 306484 16144 316007 16146
rect 306484 16088 315946 16144
rect 316002 16088 316007 16144
rect 306484 16086 316007 16088
rect 306484 16084 306490 16086
rect 315941 16083 316007 16086
rect 132585 8938 132651 8941
rect 284477 8938 284543 8941
rect 132585 8936 284543 8938
rect 132585 8880 132590 8936
rect 132646 8880 284482 8936
rect 284538 8880 284543 8936
rect 132585 8878 284543 8880
rect 132585 8875 132651 8878
rect 284477 8875 284543 8878
rect 251214 8332 251220 8396
rect 251284 8394 251290 8396
rect 251357 8394 251423 8397
rect 251284 8392 251423 8394
rect 251284 8336 251362 8392
rect 251418 8336 251423 8392
rect 251284 8334 251423 8336
rect 251284 8332 251290 8334
rect 251357 8331 251423 8334
rect 128997 7578 129063 7581
rect 283097 7578 283163 7581
rect 128997 7576 283163 7578
rect 128997 7520 129002 7576
rect 129058 7520 283102 7576
rect 283158 7520 283163 7576
rect 128997 7518 283163 7520
rect 128997 7515 129063 7518
rect 283097 7515 283163 7518
rect -960 7170 480 7260
rect 2773 7170 2839 7173
rect -960 7168 2839 7170
rect -960 7112 2778 7168
rect 2834 7112 2839 7168
rect -960 7110 2839 7112
rect -960 7020 480 7110
rect 2773 7107 2839 7110
rect 51625 6218 51691 6221
rect 249977 6218 250043 6221
rect 51625 6216 250043 6218
rect 51625 6160 51630 6216
rect 51686 6160 249982 6216
rect 250038 6160 250043 6216
rect 51625 6158 250043 6160
rect 51625 6155 51691 6158
rect 249977 6155 250043 6158
rect 583520 5796 584960 6036
rect 312077 4994 312143 4997
rect 315941 4994 316007 4997
rect 312077 4992 316007 4994
rect 312077 4936 312082 4992
rect 312138 4936 315946 4992
rect 316002 4936 316007 4992
rect 312077 4934 316007 4936
rect 312077 4931 312143 4934
rect 315941 4931 316007 4934
rect 208669 4858 208735 4861
rect 314653 4858 314719 4861
rect 208669 4856 314719 4858
rect 208669 4800 208674 4856
rect 208730 4800 314658 4856
rect 314714 4800 314719 4856
rect 208669 4798 314719 4800
rect 208669 4795 208735 4798
rect 314653 4795 314719 4798
rect 467741 4858 467807 4861
rect 576209 4858 576275 4861
rect 467741 4856 576275 4858
rect 467741 4800 467746 4856
rect 467802 4800 576214 4856
rect 576270 4800 576275 4856
rect 467741 4798 576275 4800
rect 467741 4795 467807 4798
rect 576209 4795 576275 4798
rect 354121 4042 354187 4045
rect 358169 4042 358235 4045
rect 354121 4040 358235 4042
rect 354121 3984 354126 4040
rect 354182 3984 358174 4040
rect 358230 3984 358235 4040
rect 354121 3982 358235 3984
rect 354121 3979 354187 3982
rect 358169 3979 358235 3982
rect 350625 3906 350691 3909
rect 354213 3906 354279 3909
rect 350625 3904 354279 3906
rect 350625 3848 350630 3904
rect 350686 3848 354218 3904
rect 354274 3848 354279 3904
rect 350625 3846 354279 3848
rect 350625 3843 350691 3846
rect 354213 3843 354279 3846
rect 6453 3362 6519 3365
rect 232037 3362 232103 3365
rect 6453 3360 232103 3362
rect 6453 3304 6458 3360
rect 6514 3304 232042 3360
rect 232098 3304 232103 3360
rect 6453 3302 232103 3304
rect 6453 3299 6519 3302
rect 232037 3299 232103 3302
rect 307385 3362 307451 3365
rect 356237 3362 356303 3365
rect 307385 3360 356303 3362
rect 307385 3304 307390 3360
rect 307446 3304 356242 3360
rect 356298 3304 356303 3360
rect 307385 3302 356303 3304
rect 307385 3299 307451 3302
rect 356237 3299 356303 3302
rect 468753 3362 468819 3365
rect 580993 3362 581059 3365
rect 468753 3360 581059 3362
rect 468753 3304 468758 3360
rect 468814 3304 580998 3360
rect 581054 3304 581059 3360
rect 468753 3302 581059 3304
rect 468753 3299 468819 3302
rect 580993 3299 581059 3302
rect 353661 3090 353727 3093
rect 356789 3090 356855 3093
rect 353661 3088 356855 3090
rect 353661 3032 353666 3088
rect 353722 3032 356794 3088
rect 356850 3032 356855 3088
rect 353661 3030 356855 3032
rect 353661 3027 353727 3030
rect 356789 3027 356855 3030
<< via3 >>
rect 467236 583068 467300 583132
rect 240916 582932 240980 582996
rect 240732 582796 240796 582860
rect 467052 582660 467116 582724
rect 231716 579260 231780 579324
rect 233004 579320 233068 579324
rect 233004 579264 233018 579320
rect 233018 579264 233068 579320
rect 233004 579260 233068 579264
rect 235764 579260 235828 579324
rect 237236 579320 237300 579324
rect 237236 579264 237250 579320
rect 237250 579264 237300 579320
rect 237236 579260 237300 579264
rect 239996 579260 240060 579324
rect 241284 579260 241348 579324
rect 243308 579320 243372 579324
rect 243308 579264 243322 579320
rect 243322 579264 243372 579320
rect 243308 579260 243372 579264
rect 249564 579320 249628 579324
rect 249564 579264 249578 579320
rect 249578 579264 249628 579320
rect 249564 579260 249628 579264
rect 465580 579260 465644 579324
rect 467236 486100 467300 486164
rect 242940 340580 243004 340644
rect 249564 340580 249628 340644
rect 240916 337996 240980 338060
rect 249564 336636 249628 336700
rect 249380 327116 249444 327180
rect 249380 321404 249444 321468
rect 249012 317460 249076 317524
rect 249012 309164 249076 309228
rect 249196 308892 249260 308956
rect 249196 302228 249260 302292
rect 249196 302092 249260 302156
rect 249196 298072 249260 298076
rect 249196 298016 249246 298072
rect 249246 298016 249260 298072
rect 249196 298012 249260 298016
rect 240732 295156 240796 295220
rect 249380 288492 249444 288556
rect 249380 288356 249444 288420
rect 249196 279032 249260 279036
rect 249196 278976 249246 279032
rect 249246 278976 249260 279032
rect 249196 278972 249260 278976
rect 249196 277340 249260 277404
rect 249380 267880 249444 267884
rect 249380 267824 249430 267880
rect 249430 267824 249444 267880
rect 249380 267820 249444 267824
rect 249380 263740 249444 263804
rect 249196 263468 249260 263532
rect 249380 241844 249444 241908
rect 249196 241708 249260 241772
rect 249196 241436 249260 241500
rect 366956 241496 367020 241500
rect 366956 241440 367006 241496
rect 367006 241440 367020 241496
rect 366956 241436 367020 241440
rect 249380 240892 249444 240956
rect 366956 231976 367020 231980
rect 366956 231920 367006 231976
rect 367006 231920 367020 231976
rect 366956 231916 367020 231920
rect 249380 224980 249444 225044
rect 249564 224708 249628 224772
rect 249196 217364 249260 217428
rect 249564 217364 249628 217428
rect 249196 212528 249260 212532
rect 249196 212472 249246 212528
rect 249246 212472 249260 212528
rect 249196 212468 249260 212472
rect 249564 205396 249628 205460
rect 249564 202872 249628 202876
rect 249564 202816 249614 202872
rect 249614 202816 249628 202872
rect 249564 202812 249628 202816
rect 272196 202872 272260 202876
rect 272196 202816 272210 202872
rect 272210 202816 272260 202872
rect 272196 202812 272260 202816
rect 249380 196556 249444 196620
rect 249380 191762 249444 191826
rect 272196 190496 272260 190500
rect 272196 190440 272246 190496
rect 272246 190440 272260 190496
rect 272196 190436 272260 190440
rect 249196 182200 249260 182204
rect 249196 182144 249246 182200
rect 249246 182144 249260 182200
rect 249196 182140 249260 182144
rect 249196 180644 249260 180708
rect 249748 173844 249812 173908
rect 366956 173904 367020 173908
rect 366956 173848 367006 173904
rect 367006 173848 367020 173904
rect 366956 173844 367020 173848
rect 249380 164188 249444 164252
rect 249748 164188 249812 164252
rect 366956 164248 367020 164252
rect 366956 164192 367006 164248
rect 367006 164192 367020 164248
rect 366956 164188 367020 164192
rect 324268 157660 324332 157724
rect 249380 157388 249444 157452
rect 324268 157388 324332 157452
rect 405412 157796 405476 157860
rect 405596 157388 405660 157452
rect 467052 123116 467116 123180
rect 389404 118764 389468 118828
rect 473308 111012 473372 111076
rect 243308 110740 243372 110804
rect 280108 110800 280172 110804
rect 280108 110744 280122 110800
rect 280122 110744 280172 110800
rect 280108 110740 280172 110744
rect 296668 110740 296732 110804
rect 280108 110528 280172 110532
rect 280108 110472 280122 110528
rect 280122 110472 280172 110528
rect 280108 110468 280172 110472
rect 296668 110468 296732 110532
rect 365668 110740 365732 110804
rect 357388 110604 357452 110668
rect 405412 110876 405476 110940
rect 405596 110468 405660 110532
rect 473308 110740 473372 110804
rect 492628 110740 492692 110804
rect 492628 110468 492692 110532
rect 357388 110332 357452 110396
rect 365668 110332 365732 110396
rect 389404 108896 389468 108900
rect 389404 108840 389454 108896
rect 389454 108840 389468 108896
rect 389404 108836 389468 108840
rect 265204 96384 265268 96388
rect 265204 96328 265218 96384
rect 265218 96328 265268 96384
rect 265204 96324 265268 96328
rect 265204 89040 265268 89044
rect 265204 88984 265254 89040
rect 265254 88984 265268 89040
rect 265204 88980 265268 88984
rect 396028 87484 396092 87548
rect 405596 87484 405660 87548
rect 299428 87348 299492 87412
rect 481588 87348 481652 87412
rect 251220 87212 251284 87276
rect 251220 87136 251284 87140
rect 251220 87080 251234 87136
rect 251234 87080 251284 87136
rect 251220 87076 251284 87080
rect 307708 87212 307772 87276
rect 299428 87076 299492 87140
rect 239996 86940 240060 87004
rect 307708 86940 307772 87004
rect 357388 87076 357452 87140
rect 357572 86940 357636 87004
rect 396028 87136 396092 87140
rect 396028 87080 396042 87136
rect 396042 87080 396092 87136
rect 396028 87076 396092 87080
rect 405596 86940 405660 87004
rect 481588 87076 481652 87140
rect 376708 76468 376772 76532
rect 395844 76468 395908 76532
rect 473308 76468 473372 76532
rect 241284 76060 241348 76124
rect 376708 76060 376772 76124
rect 395844 76060 395908 76124
rect 473308 76196 473372 76260
rect 492628 76196 492692 76260
rect 492628 75924 492692 75988
rect 287100 63956 287164 64020
rect 327028 63820 327092 63884
rect 287100 63684 287164 63748
rect 237236 63548 237300 63612
rect 327028 63548 327092 63612
rect 405412 63956 405476 64020
rect 405596 63548 405660 63612
rect 233004 40156 233068 40220
rect 327028 40292 327092 40356
rect 327028 40020 327092 40084
rect 405596 40292 405660 40356
rect 405596 40020 405660 40084
rect 285628 29548 285692 29612
rect 296668 29472 296732 29476
rect 296668 29416 296682 29472
rect 296682 29416 296732 29472
rect 296668 29412 296732 29416
rect 258028 29276 258092 29340
rect 285628 29276 285692 29340
rect 396028 29548 396092 29612
rect 405596 29412 405660 29476
rect 481588 29412 481652 29476
rect 235764 29140 235828 29204
rect 296668 29140 296732 29204
rect 258028 29004 258092 29068
rect 396028 29140 396092 29204
rect 405596 29004 405660 29068
rect 481588 29140 481652 29204
rect 389404 22264 389468 22268
rect 389404 22208 389454 22264
rect 389454 22208 389468 22264
rect 389404 22204 389468 22208
rect 465580 21932 465644 21996
rect 251220 21388 251284 21452
rect 389404 18048 389468 18052
rect 389404 17992 389418 18048
rect 389418 17992 389468 18048
rect 389404 17988 389468 17992
rect 473308 17172 473372 17236
rect 231716 16764 231780 16828
rect 260972 16764 261036 16828
rect 260788 16628 260852 16692
rect 405412 17036 405476 17100
rect 306420 16492 306484 16556
rect 405596 16628 405660 16692
rect 473308 16900 473372 16964
rect 492628 16900 492692 16964
rect 492628 16628 492692 16692
rect 306420 16084 306484 16148
rect 251220 8332 251284 8396
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 231715 579324 231781 579325
rect 231715 579260 231716 579324
rect 231780 579260 231781 579324
rect 231715 579259 231781 579260
rect 233003 579324 233069 579325
rect 233003 579260 233004 579324
rect 233068 579260 233069 579324
rect 233003 579259 233069 579260
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 231718 16829 231778 579259
rect 233006 40221 233066 579259
rect 234804 560454 235404 595898
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 235763 579324 235829 579325
rect 235763 579260 235764 579324
rect 235828 579260 235829 579324
rect 235763 579259 235829 579260
rect 237235 579324 237301 579325
rect 237235 579260 237236 579324
rect 237300 579260 237301 579324
rect 237235 579259 237301 579260
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 233003 40220 233069 40221
rect 233003 40156 233004 40220
rect 233068 40156 233069 40220
rect 233003 40155 233069 40156
rect 234804 20454 235404 55898
rect 235766 29205 235826 579259
rect 237238 63613 237298 579259
rect 238404 564054 239004 599498
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 240915 582996 240981 582997
rect 240915 582932 240916 582996
rect 240980 582932 240981 582996
rect 240915 582931 240981 582932
rect 240731 582860 240797 582861
rect 240731 582796 240732 582860
rect 240796 582796 240797 582860
rect 240731 582795 240797 582796
rect 239995 579324 240061 579325
rect 239995 579260 239996 579324
rect 240060 579260 240061 579324
rect 239995 579259 240061 579260
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 237235 63612 237301 63613
rect 237235 63548 237236 63612
rect 237300 63548 237301 63612
rect 237235 63547 237301 63548
rect 238404 60054 239004 95498
rect 239998 87005 240058 579259
rect 240734 295221 240794 582795
rect 240918 338061 240978 582931
rect 241283 579324 241349 579325
rect 241283 579260 241284 579324
rect 241348 579260 241349 579324
rect 241283 579259 241349 579260
rect 240915 338060 240981 338061
rect 240915 337996 240916 338060
rect 240980 337996 240981 338060
rect 240915 337995 240981 337996
rect 240731 295220 240797 295221
rect 240731 295156 240732 295220
rect 240796 295156 240797 295220
rect 240731 295155 240797 295156
rect 239995 87004 240061 87005
rect 239995 86940 239996 87004
rect 240060 86940 240061 87004
rect 239995 86939 240061 86940
rect 241286 76125 241346 579259
rect 242004 567654 242604 603098
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 243307 579324 243373 579325
rect 243307 579260 243308 579324
rect 243372 579260 243373 579324
rect 243307 579259 243373 579260
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 243310 437610 243370 579259
rect 243126 437550 243370 437610
rect 245604 571254 246204 606698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 249563 579324 249629 579325
rect 249563 579260 249564 579324
rect 249628 579260 249629 579324
rect 249563 579259 249629 579260
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 243126 436930 243186 437550
rect 243126 436870 243370 436930
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 241654 396218 241714 404142
rect 242004 387654 242604 423098
rect 242942 413898 243002 432022
rect 242942 404378 243002 412302
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242942 350658 243002 395982
rect 242942 340645 243002 346342
rect 242939 340644 243005 340645
rect 242939 340580 242940 340644
rect 243004 340580 243005 340644
rect 242939 340579 243005 340580
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 243310 110805 243370 436870
rect 245604 427254 246204 462698
rect 249566 432170 249626 579259
rect 249382 432110 249626 432170
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 249382 431578 249442 432110
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 249566 346578 249626 349062
rect 249563 340644 249629 340645
rect 249563 340580 249564 340644
rect 249628 340580 249629 340644
rect 249563 340579 249629 340580
rect 249566 336701 249626 340579
rect 249563 336700 249629 336701
rect 249563 336636 249564 336700
rect 249628 336636 249629 336700
rect 249563 336635 249629 336636
rect 249379 327180 249445 327181
rect 249379 327116 249380 327180
rect 249444 327116 249445 327180
rect 249379 327115 249445 327116
rect 249382 321469 249442 327115
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 249379 321468 249445 321469
rect 249379 321404 249380 321468
rect 249444 321404 249445 321468
rect 249379 321403 249445 321404
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 249011 317524 249077 317525
rect 249011 317460 249012 317524
rect 249076 317460 249077 317524
rect 249011 317459 249077 317460
rect 249014 309229 249074 317459
rect 249011 309228 249077 309229
rect 249011 309164 249012 309228
rect 249076 309164 249077 309228
rect 249011 309163 249077 309164
rect 249195 308956 249261 308957
rect 249195 308892 249196 308956
rect 249260 308892 249261 308956
rect 249195 308891 249261 308892
rect 249198 302293 249258 308891
rect 249195 302292 249261 302293
rect 249195 302228 249196 302292
rect 249260 302228 249261 302292
rect 249195 302227 249261 302228
rect 249195 302156 249261 302157
rect 249195 302092 249196 302156
rect 249260 302092 249261 302156
rect 249195 302091 249261 302092
rect 249198 298077 249258 302091
rect 249195 298076 249261 298077
rect 249195 298012 249196 298076
rect 249260 298012 249261 298076
rect 249195 298011 249261 298012
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 249379 288556 249445 288557
rect 249379 288492 249380 288556
rect 249444 288492 249445 288556
rect 249379 288491 249445 288492
rect 249382 288421 249442 288491
rect 249379 288420 249445 288421
rect 249379 288356 249380 288420
rect 249444 288356 249445 288420
rect 249379 288355 249445 288356
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 249195 279036 249261 279037
rect 249195 278972 249196 279036
rect 249260 278972 249261 279036
rect 249195 278971 249261 278972
rect 249198 277405 249258 278971
rect 249195 277404 249261 277405
rect 249195 277340 249196 277404
rect 249260 277340 249261 277404
rect 249195 277339 249261 277340
rect 249379 267884 249445 267885
rect 249379 267820 249380 267884
rect 249444 267820 249445 267884
rect 249379 267819 249445 267820
rect 249382 263805 249442 267819
rect 249379 263804 249445 263805
rect 249379 263740 249380 263804
rect 249444 263740 249445 263804
rect 249379 263739 249445 263740
rect 249195 263532 249261 263533
rect 249195 263468 249196 263532
rect 249260 263468 249261 263532
rect 249195 263467 249261 263468
rect 249198 259538 249258 263467
rect 249566 253330 249626 259302
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 249382 253270 249626 253330
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 249382 241909 249442 253270
rect 249379 241908 249445 241909
rect 249379 241844 249380 241908
rect 249444 241844 249445 241908
rect 249379 241843 249445 241844
rect 249195 241772 249261 241773
rect 249195 241708 249196 241772
rect 249260 241708 249261 241772
rect 249195 241707 249261 241708
rect 249198 241501 249258 241707
rect 249195 241500 249261 241501
rect 249195 241436 249196 241500
rect 249260 241436 249261 241500
rect 249195 241435 249261 241436
rect 249379 240956 249445 240957
rect 249379 240892 249380 240956
rect 249444 240892 249445 240956
rect 249379 240891 249445 240892
rect 249382 225045 249442 240891
rect 249379 225044 249445 225045
rect 249379 224980 249380 225044
rect 249444 224980 249445 225044
rect 249379 224979 249445 224980
rect 249563 224772 249629 224773
rect 249563 224708 249564 224772
rect 249628 224708 249629 224772
rect 249563 224707 249629 224708
rect 249566 217429 249626 224707
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 249195 217428 249261 217429
rect 249195 217364 249196 217428
rect 249260 217364 249261 217428
rect 249195 217363 249261 217364
rect 249563 217428 249629 217429
rect 249563 217364 249564 217428
rect 249628 217364 249629 217428
rect 249563 217363 249629 217364
rect 249198 212533 249258 217363
rect 249195 212532 249261 212533
rect 249195 212468 249196 212532
rect 249260 212468 249261 212532
rect 249195 212467 249261 212468
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 249563 205460 249629 205461
rect 249563 205396 249564 205460
rect 249628 205396 249629 205460
rect 249563 205395 249629 205396
rect 249566 202877 249626 205395
rect 249563 202876 249629 202877
rect 249563 202812 249564 202876
rect 249628 202812 249629 202876
rect 249563 202811 249629 202812
rect 249379 196620 249445 196621
rect 249379 196556 249380 196620
rect 249444 196556 249445 196620
rect 249379 196555 249445 196556
rect 249382 191827 249442 196555
rect 249379 191826 249445 191827
rect 249379 191762 249380 191826
rect 249444 191762 249445 191826
rect 249379 191761 249445 191762
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 249195 182204 249261 182205
rect 249195 182140 249196 182204
rect 249260 182140 249261 182204
rect 249195 182139 249261 182140
rect 249198 180709 249258 182139
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 249195 180708 249261 180709
rect 249195 180644 249196 180708
rect 249260 180644 249261 180708
rect 249195 180643 249261 180644
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 249747 173908 249813 173909
rect 249747 173844 249748 173908
rect 249812 173844 249813 173908
rect 249747 173843 249813 173844
rect 249750 164253 249810 173843
rect 249379 164252 249445 164253
rect 249379 164188 249380 164252
rect 249444 164188 249445 164252
rect 249379 164187 249445 164188
rect 249747 164252 249813 164253
rect 249747 164188 249748 164252
rect 249812 164188 249813 164252
rect 249747 164187 249813 164188
rect 249382 157453 249442 164187
rect 249379 157452 249445 157453
rect 249379 157388 249380 157452
rect 249444 157388 249445 157452
rect 249379 157387 249445 157388
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 243307 110804 243373 110805
rect 243307 110740 243308 110804
rect 243372 110740 243373 110804
rect 243307 110739 243373 110740
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 241283 76124 241349 76125
rect 241283 76060 241284 76124
rect 241348 76060 241349 76124
rect 241283 76059 241349 76060
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 235763 29204 235829 29205
rect 235763 29140 235764 29204
rect 235828 29140 235829 29204
rect 235763 29139 235829 29140
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 231715 16828 231781 16829
rect 231715 16764 231716 16828
rect 231780 16764 231781 16828
rect 231715 16763 231781 16764
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 251219 87276 251285 87277
rect 251219 87212 251220 87276
rect 251284 87212 251285 87276
rect 251219 87211 251285 87212
rect 251222 87141 251282 87211
rect 251219 87140 251285 87141
rect 251219 87076 251220 87140
rect 251284 87076 251285 87140
rect 251219 87075 251285 87076
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 251219 21452 251285 21453
rect 251219 21388 251220 21452
rect 251284 21388 251285 21452
rect 251219 21387 251285 21388
rect 251222 8397 251282 21387
rect 251219 8396 251285 8397
rect 251219 8332 251220 8396
rect 251284 8332 251285 8396
rect 251219 8331 251285 8332
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 258027 29340 258093 29341
rect 258027 29276 258028 29340
rect 258092 29276 258093 29340
rect 258027 29275 258093 29276
rect 258030 29069 258090 29275
rect 258027 29068 258093 29069
rect 258027 29004 258028 29068
rect 258092 29004 258093 29068
rect 258027 29003 258093 29004
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 9654 260604 45098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 272195 202876 272261 202877
rect 272195 202812 272196 202876
rect 272260 202812 272261 202876
rect 272195 202811 272261 202812
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 272198 190501 272258 202811
rect 272195 190500 272261 190501
rect 272195 190436 272196 190500
rect 272260 190436 272261 190500
rect 272195 190435 272261 190436
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 265203 96388 265269 96389
rect 265203 96324 265204 96388
rect 265268 96324 265269 96388
rect 265203 96323 265269 96324
rect 265206 89045 265266 96323
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 265203 89044 265269 89045
rect 265203 88980 265204 89044
rect 265268 88980 265269 89044
rect 265203 88979 265269 88980
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 260971 16828 261037 16829
rect 260971 16764 260972 16828
rect 261036 16764 261037 16828
rect 260971 16763 261037 16764
rect 260787 16692 260853 16693
rect 260787 16628 260788 16692
rect 260852 16690 260853 16692
rect 260974 16690 261034 16763
rect 260852 16630 261034 16690
rect 260852 16628 260853 16630
rect 260787 16627 260853 16628
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 280107 110804 280173 110805
rect 280107 110740 280108 110804
rect 280172 110740 280173 110804
rect 280107 110739 280173 110740
rect 280110 110533 280170 110739
rect 280107 110532 280173 110533
rect 280107 110468 280108 110532
rect 280172 110468 280173 110532
rect 280107 110467 280173 110468
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 287099 64020 287165 64021
rect 287099 63956 287100 64020
rect 287164 63956 287165 64020
rect 287099 63955 287165 63956
rect 287102 63749 287162 63955
rect 287099 63748 287165 63749
rect 287099 63684 287100 63748
rect 287164 63684 287165 63748
rect 287099 63683 287165 63684
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 285627 29612 285693 29613
rect 285627 29548 285628 29612
rect 285692 29548 285693 29612
rect 285627 29547 285693 29548
rect 285630 29341 285690 29547
rect 285627 29340 285693 29341
rect 285627 29276 285628 29340
rect 285692 29276 285693 29340
rect 285627 29275 285693 29276
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 296667 110804 296733 110805
rect 296667 110740 296668 110804
rect 296732 110740 296733 110804
rect 296667 110739 296733 110740
rect 296670 110533 296730 110739
rect 296667 110532 296733 110533
rect 296667 110468 296668 110532
rect 296732 110468 296733 110532
rect 296667 110467 296733 110468
rect 299427 87412 299493 87413
rect 299427 87348 299428 87412
rect 299492 87348 299493 87412
rect 299427 87347 299493 87348
rect 299430 87141 299490 87347
rect 299427 87140 299493 87141
rect 299427 87076 299428 87140
rect 299492 87076 299493 87140
rect 299427 87075 299493 87076
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 296667 29476 296733 29477
rect 296667 29412 296668 29476
rect 296732 29412 296733 29476
rect 296667 29411 296733 29412
rect 296670 29205 296730 29411
rect 296667 29204 296733 29205
rect 296667 29140 296668 29204
rect 296732 29140 296733 29204
rect 296667 29139 296733 29140
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 13254 300204 48698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 307707 87276 307773 87277
rect 307707 87212 307708 87276
rect 307772 87212 307773 87276
rect 307707 87211 307773 87212
rect 307710 87005 307770 87211
rect 307707 87004 307773 87005
rect 307707 86940 307708 87004
rect 307772 86940 307773 87004
rect 307707 86939 307773 86940
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306419 16556 306485 16557
rect 306419 16492 306420 16556
rect 306484 16492 306485 16556
rect 306419 16491 306485 16492
rect 306422 16149 306482 16491
rect 306419 16148 306485 16149
rect 306419 16084 306420 16148
rect 306484 16084 306485 16148
rect 306419 16083 306485 16084
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324267 157724 324333 157725
rect 324267 157660 324268 157724
rect 324332 157660 324333 157724
rect 324267 157659 324333 157660
rect 324270 157453 324330 157659
rect 324267 157452 324333 157453
rect 324267 157388 324268 157452
rect 324332 157388 324333 157452
rect 324267 157387 324333 157388
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 327027 63884 327093 63885
rect 327027 63820 327028 63884
rect 327092 63820 327093 63884
rect 327027 63819 327093 63820
rect 327030 63613 327090 63819
rect 327027 63612 327093 63613
rect 327027 63548 327028 63612
rect 327092 63548 327093 63612
rect 327027 63547 327093 63548
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 327027 40356 327093 40357
rect 327027 40292 327028 40356
rect 327092 40292 327093 40356
rect 327027 40291 327093 40292
rect 327030 40085 327090 40291
rect 327027 40084 327093 40085
rect 327027 40020 327028 40084
rect 327092 40020 327093 40084
rect 327027 40019 327093 40020
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 357387 110668 357453 110669
rect 357387 110604 357388 110668
rect 357452 110604 357453 110668
rect 357387 110603 357453 110604
rect 357390 110397 357450 110603
rect 360804 110454 361404 145898
rect 357387 110396 357453 110397
rect 357387 110332 357388 110396
rect 357452 110332 357453 110396
rect 357387 110331 357453 110332
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 357390 87350 357634 87410
rect 357390 87141 357450 87350
rect 357387 87140 357453 87141
rect 357387 87076 357388 87140
rect 357452 87076 357453 87140
rect 357387 87075 357453 87076
rect 357574 87005 357634 87350
rect 357571 87004 357637 87005
rect 357571 86940 357572 87004
rect 357636 86940 357637 87004
rect 357571 86939 357637 86940
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 366955 241500 367021 241501
rect 366955 241436 366956 241500
rect 367020 241436 367021 241500
rect 366955 241435 367021 241436
rect 366958 231981 367018 241435
rect 366955 231980 367021 231981
rect 366955 231916 366956 231980
rect 367020 231916 367021 231980
rect 366955 231915 367021 231916
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 366955 173908 367021 173909
rect 366955 173844 366956 173908
rect 367020 173844 367021 173908
rect 366955 173843 367021 173844
rect 366958 164253 367018 173843
rect 366955 164252 367021 164253
rect 366955 164188 366956 164252
rect 367020 164188 367021 164252
rect 366955 164187 367021 164188
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 365667 110804 365733 110805
rect 365667 110740 365668 110804
rect 365732 110740 365733 110804
rect 365667 110739 365733 110740
rect 365670 110397 365730 110739
rect 365667 110396 365733 110397
rect 365667 110332 365668 110396
rect 365732 110332 365733 110396
rect 365667 110331 365733 110332
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 376707 76532 376773 76533
rect 376707 76468 376708 76532
rect 376772 76468 376773 76532
rect 376707 76467 376773 76468
rect 376710 76125 376770 76467
rect 376707 76124 376773 76125
rect 376707 76060 376708 76124
rect 376772 76060 376773 76124
rect 376707 76059 376773 76060
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389403 118828 389469 118829
rect 389403 118764 389404 118828
rect 389468 118764 389469 118828
rect 389403 118763 389469 118764
rect 389406 108901 389466 118763
rect 389403 108900 389469 108901
rect 389403 108836 389404 108900
rect 389468 108836 389469 108900
rect 389403 108835 389469 108836
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396027 87548 396093 87549
rect 396027 87484 396028 87548
rect 396092 87484 396093 87548
rect 396027 87483 396093 87484
rect 396030 87141 396090 87483
rect 396027 87140 396093 87141
rect 396027 87076 396028 87140
rect 396092 87076 396093 87140
rect 396027 87075 396093 87076
rect 395843 76532 395909 76533
rect 395843 76468 395844 76532
rect 395908 76468 395909 76532
rect 395843 76467 395909 76468
rect 395846 76125 395906 76467
rect 395843 76124 395909 76125
rect 395843 76060 395844 76124
rect 395908 76060 395909 76124
rect 395843 76059 395909 76060
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 389403 22268 389469 22269
rect 389403 22204 389404 22268
rect 389468 22204 389469 22268
rect 389403 22203 389469 22204
rect 389406 18053 389466 22203
rect 389403 18052 389469 18053
rect 389403 17988 389404 18052
rect 389468 17988 389469 18052
rect 389403 17987 389469 17988
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396027 29612 396093 29613
rect 396027 29548 396028 29612
rect 396092 29548 396093 29612
rect 396027 29547 396093 29548
rect 396030 29205 396090 29547
rect 396027 29204 396093 29205
rect 396027 29140 396028 29204
rect 396092 29140 396093 29204
rect 396027 29139 396093 29140
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 405411 157860 405477 157861
rect 405411 157796 405412 157860
rect 405476 157796 405477 157860
rect 405411 157795 405477 157796
rect 405414 157450 405474 157795
rect 405595 157452 405661 157453
rect 405595 157450 405596 157452
rect 405414 157390 405596 157450
rect 405595 157388 405596 157390
rect 405660 157388 405661 157452
rect 405595 157387 405661 157388
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 405411 110940 405477 110941
rect 405411 110876 405412 110940
rect 405476 110876 405477 110940
rect 405411 110875 405477 110876
rect 405414 110530 405474 110875
rect 405595 110532 405661 110533
rect 405595 110530 405596 110532
rect 405414 110470 405596 110530
rect 405595 110468 405596 110470
rect 405660 110468 405661 110532
rect 405595 110467 405661 110468
rect 405595 87548 405661 87549
rect 405595 87484 405596 87548
rect 405660 87484 405661 87548
rect 405595 87483 405661 87484
rect 405598 87005 405658 87483
rect 405595 87004 405661 87005
rect 405595 86940 405596 87004
rect 405660 86940 405661 87004
rect 405595 86939 405661 86940
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 405411 64020 405477 64021
rect 405411 63956 405412 64020
rect 405476 63956 405477 64020
rect 405411 63955 405477 63956
rect 405414 63610 405474 63955
rect 405595 63612 405661 63613
rect 405595 63610 405596 63612
rect 405414 63550 405596 63610
rect 405595 63548 405596 63550
rect 405660 63548 405661 63612
rect 405595 63547 405661 63548
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 405595 40356 405661 40357
rect 405595 40292 405596 40356
rect 405660 40292 405661 40356
rect 405595 40291 405661 40292
rect 405598 40085 405658 40291
rect 405595 40084 405661 40085
rect 405595 40020 405596 40084
rect 405660 40020 405661 40084
rect 405595 40019 405661 40020
rect 405595 29476 405661 29477
rect 405595 29412 405596 29476
rect 405660 29412 405661 29476
rect 405595 29411 405661 29412
rect 405598 29069 405658 29411
rect 405595 29068 405661 29069
rect 405595 29004 405596 29068
rect 405660 29004 405661 29068
rect 405595 29003 405661 29004
rect 405411 17100 405477 17101
rect 405411 17036 405412 17100
rect 405476 17036 405477 17100
rect 405411 17035 405477 17036
rect 405414 16690 405474 17035
rect 405595 16692 405661 16693
rect 405595 16690 405596 16692
rect 405414 16630 405596 16690
rect 405595 16628 405596 16630
rect 405660 16628 405661 16692
rect 405595 16627 405661 16628
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 467235 583132 467301 583133
rect 467235 583068 467236 583132
rect 467300 583068 467301 583132
rect 467235 583067 467301 583068
rect 467051 582724 467117 582725
rect 467051 582660 467052 582724
rect 467116 582660 467117 582724
rect 467051 582659 467117 582660
rect 465579 579324 465645 579325
rect 465579 579260 465580 579324
rect 465644 579260 465645 579324
rect 465579 579259 465645 579260
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 465582 21997 465642 579259
rect 467054 123181 467114 582659
rect 467238 486165 467298 583067
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 467235 486164 467301 486165
rect 467235 486100 467236 486164
rect 467300 486100 467301 486164
rect 467235 486099 467301 486100
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 467051 123180 467117 123181
rect 467051 123116 467052 123180
rect 467116 123116 467117 123180
rect 467051 123115 467117 123116
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 465579 21996 465645 21997
rect 465579 21932 465580 21996
rect 465644 21932 465645 21996
rect 465579 21931 465645 21932
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 473307 111076 473373 111077
rect 473307 111012 473308 111076
rect 473372 111012 473373 111076
rect 473307 111011 473373 111012
rect 473310 110805 473370 111011
rect 473307 110804 473373 110805
rect 473307 110740 473308 110804
rect 473372 110740 473373 110804
rect 473307 110739 473373 110740
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 473307 76532 473373 76533
rect 473307 76468 473308 76532
rect 473372 76468 473373 76532
rect 473307 76467 473373 76468
rect 473310 76261 473370 76467
rect 473307 76260 473373 76261
rect 473307 76196 473308 76260
rect 473372 76196 473373 76260
rect 473307 76195 473373 76196
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 473307 17236 473373 17237
rect 473307 17172 473308 17236
rect 473372 17172 473373 17236
rect 473307 17171 473373 17172
rect 473310 16965 473370 17171
rect 473307 16964 473373 16965
rect 473307 16900 473308 16964
rect 473372 16900 473373 16964
rect 473307 16899 473373 16900
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 481587 87412 481653 87413
rect 481587 87348 481588 87412
rect 481652 87348 481653 87412
rect 481587 87347 481653 87348
rect 481590 87141 481650 87347
rect 481587 87140 481653 87141
rect 481587 87076 481588 87140
rect 481652 87076 481653 87140
rect 481587 87075 481653 87076
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 481587 29476 481653 29477
rect 481587 29412 481588 29476
rect 481652 29412 481653 29476
rect 481587 29411 481653 29412
rect 481590 29205 481650 29411
rect 481587 29204 481653 29205
rect 481587 29140 481588 29204
rect 481652 29140 481653 29204
rect 481587 29139 481653 29140
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 492627 110804 492693 110805
rect 492627 110740 492628 110804
rect 492692 110740 492693 110804
rect 492627 110739 492693 110740
rect 492630 110533 492690 110739
rect 492627 110532 492693 110533
rect 492627 110468 492628 110532
rect 492692 110468 492693 110532
rect 492627 110467 492693 110468
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 492627 76260 492693 76261
rect 492627 76196 492628 76260
rect 492692 76196 492693 76260
rect 492627 76195 492693 76196
rect 492630 75989 492690 76195
rect 492627 75988 492693 75989
rect 492627 75924 492628 75988
rect 492692 75924 492693 75988
rect 492627 75923 492693 75924
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 492627 16964 492693 16965
rect 492627 16900 492628 16964
rect 492692 16900 492693 16964
rect 492627 16899 492693 16900
rect 492630 16693 492690 16899
rect 492627 16692 492693 16693
rect 492627 16628 492628 16692
rect 492692 16628 492693 16692
rect 492627 16627 492693 16628
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 242854 432022 243090 432258
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 241566 404142 241802 404378
rect 241566 395982 241802 396218
rect 242854 413662 243090 413898
rect 242854 412302 243090 412538
rect 242854 404142 243090 404378
rect 242854 395982 243090 396218
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242854 350422 243090 350658
rect 242854 346342 243090 346578
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 249294 431342 249530 431578
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 249478 349062 249714 349298
rect 249478 346342 249714 346578
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 249110 259302 249346 259538
rect 249478 259302 249714 259538
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect 242812 432258 248284 432300
rect 242812 432022 242854 432258
rect 243090 432022 248284 432258
rect 242812 431980 248284 432022
rect 247964 431620 248284 431980
rect 247964 431578 249572 431620
rect 247964 431342 249294 431578
rect 249530 431342 249572 431578
rect 247964 431300 249572 431342
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect 242812 413898 243316 413940
rect 242812 413662 242854 413898
rect 243090 413662 243316 413898
rect 242812 413620 243316 413662
rect 242996 412580 243316 413620
rect 242812 412538 243316 412580
rect 242812 412302 242854 412538
rect 243090 412302 243316 412538
rect 242812 412260 243316 412302
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect 241524 404378 243132 404420
rect 241524 404142 241566 404378
rect 241802 404142 242854 404378
rect 243090 404142 243132 404378
rect 241524 404100 243132 404142
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect 241524 396218 243132 396260
rect 241524 395982 241566 396218
rect 241802 395982 242854 396218
rect 243090 395982 243132 396218
rect 241524 395940 243132 395982
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect 242812 350658 249756 350700
rect 242812 350422 242854 350658
rect 243090 350422 249756 350658
rect 242812 350380 249756 350422
rect 249436 349298 249756 350380
rect 249436 349062 249478 349298
rect 249714 349062 249756 349298
rect 249436 349020 249756 349062
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect 242812 346578 249756 346620
rect 242812 346342 242854 346578
rect 243090 346342 249478 346578
rect 249714 346342 249756 346578
rect 242812 346300 249756 346342
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect 249068 259538 249756 259580
rect 249068 259302 249110 259538
rect 249346 259302 249478 259538
rect 249714 259302 249756 259538
rect 249068 259260 249756 259302
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use user_proj_example  mprj
timestamp 1608158347
transform 1 0 230000 0 1 340000
box 0 0 239540 240000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
